----------------------------------------------------------------
-- Copyright 2020 University of Alberta

-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at

--     http://www.apache.org/licenses/LICENSE-2.0

-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
----------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.vnir;

package img_buffer_pkg is
    --Generating 10 buffers for each, allowing for storage of up to 10 rows
    constant NUM_SWIR_ROW_FIFO : integer := 10;
    constant NUM_VNIR_ROW_FIFO : integer := 10;

    --Number of bits in swir and vnir fifo
    constant SWIR_FIFO_WORD_LENGTH : integer := 64;
    constant VNIR_FIFO_WORD_LENGTH : integer := 160;

    --vnir & swir row fragments are split into their respective FIFO word lengths
    subtype vnir_fragment_t is std_logic_vector (VNIR_FIFO_WORD_LENGTH-1 downto 0);
    subtype swir_fragment_t is std_logic_vector (SWIR_FIFO_WORD_LENGTH-1 downto 0);

    --The links between the vnir and swir fifos
    type vnir_link_a is array of (0 to NUM_VNIR_ROW_FIFO-1) of vnir_fragement_t;
    type swir_link_a is array of (0 to NUM_SWIR_ROW_FIFO-1) of swir_fragment_t;

    type row_type_buffer_a is array of (0 to NUM_VNIR_ROW_FIFO-1) of vnir.row_type_t;

    
end package img_buffer_pkg;
