----------------------------------------------------------------
-- Copyright 2020 University of Alberta

-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at

--     http://www.apache.org/licenses/LICENSE-2.0

-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
----------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.spi_types.all;
use work.vnir_types.all;

entity collate_rows_tb is
end entity;

architecture tests of collate_rows_tb is

	constant clock_period	: time := 20 ns;

	signal clock            : std_logic := '0';
	signal reset_n          : std_logic := '1';
	signal pixels           : vnir_pixel_vector_t(0 to 4-1);
	signal pixels_available	: std_logic := '0';
	signal row_red          : vnir_row_t;
	signal row_blue         : vnir_row_t;
	signal row_nir          : vnir_row_t;
	signal rows_available   : std_logic := '0';

    component collate_rows is
    port (
        clock            : in std_logic;
        reset_n          : in std_logic;
        pixels_in        : in vnir_pixel_vector_t(0 to 4-1);
        pixels_available : in std_logic;
        red              : out vnir_row_t;
        blue             : out vnir_row_t;
        nir              : out vnir_row_t;
        rows_available   : out std_logic
    );
    end component collate_rows;

    type vnir_row_window_t is array(0 to 9) of vnir_row_t;
    type data_t is array(0 to 2) of vnir_row_window_t;
    constant data : data_t := (
        0 => (
            0 => (0 => to_unsigned(2732, 12), 1 => to_unsigned(2607, 12), 2 => to_unsigned(1653, 12), 3 => to_unsigned(3264, 12), 4 => to_unsigned(835, 12), 5 => to_unsigned(763, 12), 6 => to_unsigned(1731, 12), 7 => to_unsigned(3431, 12), 8 => to_unsigned(1033, 12), 9 => to_unsigned(3795, 12), 10 => to_unsigned(277, 12), 11 => to_unsigned(1778, 12), 12 => to_unsigned(1828, 12), 13 => to_unsigned(2647, 12), 14 => to_unsigned(3142, 12), 15 => to_unsigned(3544, 12), 16 => to_unsigned(2648, 12), 17 => to_unsigned(3468, 12), 18 => to_unsigned(2362, 12), 19 => to_unsigned(705, 12), 20 => to_unsigned(3558, 12), 21 => to_unsigned(2599, 12), 22 => to_unsigned(2135, 12), 23 => to_unsigned(2222, 12), 24 => to_unsigned(3672, 12), 25 => to_unsigned(2897, 12), 26 => to_unsigned(1701, 12), 27 => to_unsigned(537, 12), 28 => to_unsigned(2893, 12), 29 => to_unsigned(2120, 12), 30 => to_unsigned(2825, 12), 31 => to_unsigned(1940, 12), 32 => to_unsigned(2163, 12), 33 => to_unsigned(976, 12), 34 => to_unsigned(755, 12), 35 => to_unsigned(3781, 12), 36 => to_unsigned(2046, 12), 37 => to_unsigned(1871, 12), 38 => to_unsigned(3503, 12), 39 => to_unsigned(2496, 12), 40 => to_unsigned(2898, 12), 41 => to_unsigned(99, 12), 42 => to_unsigned(2008, 12), 43 => to_unsigned(3249, 12), 44 => to_unsigned(755, 12), 45 => to_unsigned(797, 12), 46 => to_unsigned(659, 12), 47 => to_unsigned(3219, 12), 48 => to_unsigned(2958, 12), 49 => to_unsigned(423, 12), 50 => to_unsigned(3360, 12), 51 => to_unsigned(4033, 12), 52 => to_unsigned(3337, 12), 53 => to_unsigned(2745, 12), 54 => to_unsigned(639, 12), 55 => to_unsigned(544, 12), 56 => to_unsigned(2591, 12), 57 => to_unsigned(714, 12), 58 => to_unsigned(2292, 12), 59 => to_unsigned(151, 12), 60 => to_unsigned(2723, 12), 61 => to_unsigned(2558, 12), 62 => to_unsigned(3531, 12), 63 => to_unsigned(2930, 12), 64 => to_unsigned(1207, 12), 65 => to_unsigned(2076, 12), 66 => to_unsigned(802, 12), 67 => to_unsigned(2176, 12), 68 => to_unsigned(2176, 12), 69 => to_unsigned(1956, 12), 70 => to_unsigned(3125, 12), 71 => to_unsigned(1925, 12), 72 => to_unsigned(3622, 12), 73 => to_unsigned(3560, 12), 74 => to_unsigned(756, 12), 75 => to_unsigned(273, 12), 76 => to_unsigned(2383, 12), 77 => to_unsigned(388, 12), 78 => to_unsigned(1641, 12), 79 => to_unsigned(3114, 12), 80 => to_unsigned(1466, 12), 81 => to_unsigned(2591, 12), 82 => to_unsigned(888, 12), 83 => to_unsigned(257, 12), 84 => to_unsigned(1345, 12), 85 => to_unsigned(4071, 12), 86 => to_unsigned(4009, 12), 87 => to_unsigned(2105, 12), 88 => to_unsigned(2339, 12), 89 => to_unsigned(3942, 12), 90 => to_unsigned(3191, 12), 91 => to_unsigned(2827, 12), 92 => to_unsigned(430, 12), 93 => to_unsigned(3154, 12), 94 => to_unsigned(91, 12), 95 => to_unsigned(1920, 12), 96 => to_unsigned(2446, 12), 97 => to_unsigned(2659, 12), 98 => to_unsigned(1589, 12), 99 => to_unsigned(2956, 12), 100 => to_unsigned(2681, 12), 101 => to_unsigned(4010, 12), 102 => to_unsigned(84, 12), 103 => to_unsigned(2251, 12), 104 => to_unsigned(324, 12), 105 => to_unsigned(774, 12), 106 => to_unsigned(3012, 12), 107 => to_unsigned(1071, 12), 108 => to_unsigned(639, 12), 109 => to_unsigned(2036, 12), 110 => to_unsigned(1155, 12), 111 => to_unsigned(972, 12), 112 => to_unsigned(2916, 12), 113 => to_unsigned(1204, 12), 114 => to_unsigned(2024, 12), 115 => to_unsigned(3918, 12), 116 => to_unsigned(1167, 12), 117 => to_unsigned(1684, 12), 118 => to_unsigned(3299, 12), 119 => to_unsigned(3002, 12), 120 => to_unsigned(2839, 12), 121 => to_unsigned(2767, 12), 122 => to_unsigned(2957, 12), 123 => to_unsigned(373, 12), 124 => to_unsigned(1877, 12), 125 => to_unsigned(560, 12), 126 => to_unsigned(1329, 12), 127 => to_unsigned(1605, 12), 128 => to_unsigned(2217, 12), 129 => to_unsigned(1699, 12), 130 => to_unsigned(1472, 12), 131 => to_unsigned(3167, 12), 132 => to_unsigned(3269, 12), 133 => to_unsigned(3678, 12), 134 => to_unsigned(256, 12), 135 => to_unsigned(1905, 12), 136 => to_unsigned(3762, 12), 137 => to_unsigned(1316, 12), 138 => to_unsigned(1954, 12), 139 => to_unsigned(816, 12), 140 => to_unsigned(3933, 12), 141 => to_unsigned(2435, 12), 142 => to_unsigned(1634, 12), 143 => to_unsigned(3626, 12), 144 => to_unsigned(973, 12), 145 => to_unsigned(368, 12), 146 => to_unsigned(2023, 12), 147 => to_unsigned(2965, 12), 148 => to_unsigned(201, 12), 149 => to_unsigned(2431, 12), 150 => to_unsigned(1536, 12), 151 => to_unsigned(1930, 12), 152 => to_unsigned(2418, 12), 153 => to_unsigned(555, 12), 154 => to_unsigned(954, 12), 155 => to_unsigned(3455, 12), 156 => to_unsigned(2071, 12), 157 => to_unsigned(1723, 12), 158 => to_unsigned(130, 12), 159 => to_unsigned(2425, 12), 160 => to_unsigned(2146, 12), 161 => to_unsigned(3646, 12), 162 => to_unsigned(931, 12), 163 => to_unsigned(2782, 12), 164 => to_unsigned(2171, 12), 165 => to_unsigned(1987, 12), 166 => to_unsigned(2642, 12), 167 => to_unsigned(1966, 12), 168 => to_unsigned(2787, 12), 169 => to_unsigned(3220, 12), 170 => to_unsigned(209, 12), 171 => to_unsigned(2610, 12), 172 => to_unsigned(1435, 12), 173 => to_unsigned(2830, 12), 174 => to_unsigned(3113, 12), 175 => to_unsigned(3130, 12), 176 => to_unsigned(2753, 12), 177 => to_unsigned(3108, 12), 178 => to_unsigned(2826, 12), 179 => to_unsigned(86, 12), 180 => to_unsigned(3115, 12), 181 => to_unsigned(872, 12), 182 => to_unsigned(2059, 12), 183 => to_unsigned(2818, 12), 184 => to_unsigned(307, 12), 185 => to_unsigned(1104, 12), 186 => to_unsigned(2080, 12), 187 => to_unsigned(1206, 12), 188 => to_unsigned(1152, 12), 189 => to_unsigned(2854, 12), 190 => to_unsigned(275, 12), 191 => to_unsigned(1198, 12), 192 => to_unsigned(1578, 12), 193 => to_unsigned(1395, 12), 194 => to_unsigned(1208, 12), 195 => to_unsigned(2492, 12), 196 => to_unsigned(2536, 12), 197 => to_unsigned(3661, 12), 198 => to_unsigned(2334, 12), 199 => to_unsigned(1304, 12), 200 => to_unsigned(637, 12), 201 => to_unsigned(770, 12), 202 => to_unsigned(3587, 12), 203 => to_unsigned(94, 12), 204 => to_unsigned(3298, 12), 205 => to_unsigned(1899, 12), 206 => to_unsigned(3341, 12), 207 => to_unsigned(1904, 12), 208 => to_unsigned(2344, 12), 209 => to_unsigned(1352, 12), 210 => to_unsigned(3091, 12), 211 => to_unsigned(607, 12), 212 => to_unsigned(3912, 12), 213 => to_unsigned(1434, 12), 214 => to_unsigned(2498, 12), 215 => to_unsigned(1272, 12), 216 => to_unsigned(180, 12), 217 => to_unsigned(2371, 12), 218 => to_unsigned(3052, 12), 219 => to_unsigned(3901, 12), 220 => to_unsigned(3854, 12), 221 => to_unsigned(3936, 12), 222 => to_unsigned(3332, 12), 223 => to_unsigned(4035, 12), 224 => to_unsigned(749, 12), 225 => to_unsigned(2187, 12), 226 => to_unsigned(1020, 12), 227 => to_unsigned(2646, 12), 228 => to_unsigned(3533, 12), 229 => to_unsigned(2937, 12), 230 => to_unsigned(1645, 12), 231 => to_unsigned(843, 12), 232 => to_unsigned(2744, 12), 233 => to_unsigned(1552, 12), 234 => to_unsigned(3224, 12), 235 => to_unsigned(925, 12), 236 => to_unsigned(2197, 12), 237 => to_unsigned(1134, 12), 238 => to_unsigned(25, 12), 239 => to_unsigned(1488, 12), 240 => to_unsigned(956, 12), 241 => to_unsigned(1913, 12), 242 => to_unsigned(2934, 12), 243 => to_unsigned(1141, 12), 244 => to_unsigned(1469, 12), 245 => to_unsigned(1619, 12), 246 => to_unsigned(2721, 12), 247 => to_unsigned(1896, 12), 248 => to_unsigned(928, 12), 249 => to_unsigned(3300, 12), 250 => to_unsigned(1531, 12), 251 => to_unsigned(2811, 12), 252 => to_unsigned(2169, 12), 253 => to_unsigned(1350, 12), 254 => to_unsigned(469, 12), 255 => to_unsigned(2335, 12), 256 => to_unsigned(525, 12), 257 => to_unsigned(1863, 12), 258 => to_unsigned(1720, 12), 259 => to_unsigned(1176, 12), 260 => to_unsigned(591, 12), 261 => to_unsigned(2089, 12), 262 => to_unsigned(2322, 12), 263 => to_unsigned(3624, 12), 264 => to_unsigned(3510, 12), 265 => to_unsigned(207, 12), 266 => to_unsigned(2827, 12), 267 => to_unsigned(166, 12), 268 => to_unsigned(2159, 12), 269 => to_unsigned(3421, 12), 270 => to_unsigned(4089, 12), 271 => to_unsigned(1153, 12), 272 => to_unsigned(2783, 12), 273 => to_unsigned(1910, 12), 274 => to_unsigned(2860, 12), 275 => to_unsigned(216, 12), 276 => to_unsigned(3453, 12), 277 => to_unsigned(24, 12), 278 => to_unsigned(67, 12), 279 => to_unsigned(3026, 12), 280 => to_unsigned(1007, 12), 281 => to_unsigned(3843, 12), 282 => to_unsigned(2282, 12), 283 => to_unsigned(1740, 12), 284 => to_unsigned(2022, 12), 285 => to_unsigned(291, 12), 286 => to_unsigned(1750, 12), 287 => to_unsigned(1022, 12), 288 => to_unsigned(2749, 12), 289 => to_unsigned(3781, 12), 290 => to_unsigned(2775, 12), 291 => to_unsigned(2603, 12), 292 => to_unsigned(2080, 12), 293 => to_unsigned(3083, 12), 294 => to_unsigned(1640, 12), 295 => to_unsigned(2260, 12), 296 => to_unsigned(1162, 12), 297 => to_unsigned(1718, 12), 298 => to_unsigned(4075, 12), 299 => to_unsigned(1445, 12), 300 => to_unsigned(3709, 12), 301 => to_unsigned(3740, 12), 302 => to_unsigned(623, 12), 303 => to_unsigned(3560, 12), 304 => to_unsigned(770, 12), 305 => to_unsigned(1563, 12), 306 => to_unsigned(4051, 12), 307 => to_unsigned(1241, 12), 308 => to_unsigned(2711, 12), 309 => to_unsigned(821, 12), 310 => to_unsigned(307, 12), 311 => to_unsigned(1198, 12), 312 => to_unsigned(1172, 12), 313 => to_unsigned(2997, 12), 314 => to_unsigned(1565, 12), 315 => to_unsigned(3651, 12), 316 => to_unsigned(2595, 12), 317 => to_unsigned(807, 12), 318 => to_unsigned(3465, 12), 319 => to_unsigned(2121, 12), 320 => to_unsigned(297, 12), 321 => to_unsigned(2967, 12), 322 => to_unsigned(3971, 12), 323 => to_unsigned(3886, 12), 324 => to_unsigned(730, 12), 325 => to_unsigned(1970, 12), 326 => to_unsigned(2924, 12), 327 => to_unsigned(1795, 12), 328 => to_unsigned(1823, 12), 329 => to_unsigned(2825, 12), 330 => to_unsigned(3466, 12), 331 => to_unsigned(3611, 12), 332 => to_unsigned(429, 12), 333 => to_unsigned(199, 12), 334 => to_unsigned(1447, 12), 335 => to_unsigned(1085, 12), 336 => to_unsigned(2389, 12), 337 => to_unsigned(865, 12), 338 => to_unsigned(3116, 12), 339 => to_unsigned(2850, 12), 340 => to_unsigned(1954, 12), 341 => to_unsigned(1112, 12), 342 => to_unsigned(2081, 12), 343 => to_unsigned(2693, 12), 344 => to_unsigned(2280, 12), 345 => to_unsigned(767, 12), 346 => to_unsigned(2084, 12), 347 => to_unsigned(1792, 12), 348 => to_unsigned(1483, 12), 349 => to_unsigned(2338, 12), 350 => to_unsigned(197, 12), 351 => to_unsigned(894, 12), 352 => to_unsigned(1973, 12), 353 => to_unsigned(1278, 12), 354 => to_unsigned(3152, 12), 355 => to_unsigned(1470, 12), 356 => to_unsigned(136, 12), 357 => to_unsigned(2237, 12), 358 => to_unsigned(2177, 12), 359 => to_unsigned(2257, 12), 360 => to_unsigned(1392, 12), 361 => to_unsigned(2339, 12), 362 => to_unsigned(1400, 12), 363 => to_unsigned(3419, 12), 364 => to_unsigned(168, 12), 365 => to_unsigned(1908, 12), 366 => to_unsigned(2852, 12), 367 => to_unsigned(176, 12), 368 => to_unsigned(1561, 12), 369 => to_unsigned(323, 12), 370 => to_unsigned(3943, 12), 371 => to_unsigned(508, 12), 372 => to_unsigned(2851, 12), 373 => to_unsigned(3186, 12), 374 => to_unsigned(1822, 12), 375 => to_unsigned(1053, 12), 376 => to_unsigned(1777, 12), 377 => to_unsigned(3361, 12), 378 => to_unsigned(146, 12), 379 => to_unsigned(1297, 12), 380 => to_unsigned(221, 12), 381 => to_unsigned(2388, 12), 382 => to_unsigned(509, 12), 383 => to_unsigned(2562, 12), 384 => to_unsigned(2117, 12), 385 => to_unsigned(1381, 12), 386 => to_unsigned(908, 12), 387 => to_unsigned(556, 12), 388 => to_unsigned(885, 12), 389 => to_unsigned(2813, 12), 390 => to_unsigned(1346, 12), 391 => to_unsigned(3695, 12), 392 => to_unsigned(2139, 12), 393 => to_unsigned(3413, 12), 394 => to_unsigned(423, 12), 395 => to_unsigned(3623, 12), 396 => to_unsigned(4043, 12), 397 => to_unsigned(3734, 12), 398 => to_unsigned(3486, 12), 399 => to_unsigned(3729, 12), 400 => to_unsigned(2758, 12), 401 => to_unsigned(967, 12), 402 => to_unsigned(274, 12), 403 => to_unsigned(860, 12), 404 => to_unsigned(2091, 12), 405 => to_unsigned(1107, 12), 406 => to_unsigned(433, 12), 407 => to_unsigned(809, 12), 408 => to_unsigned(2141, 12), 409 => to_unsigned(1198, 12), 410 => to_unsigned(1429, 12), 411 => to_unsigned(201, 12), 412 => to_unsigned(3929, 12), 413 => to_unsigned(2546, 12), 414 => to_unsigned(2528, 12), 415 => to_unsigned(2011, 12), 416 => to_unsigned(329, 12), 417 => to_unsigned(3612, 12), 418 => to_unsigned(4075, 12), 419 => to_unsigned(209, 12), 420 => to_unsigned(2665, 12), 421 => to_unsigned(1978, 12), 422 => to_unsigned(3968, 12), 423 => to_unsigned(4054, 12), 424 => to_unsigned(3647, 12), 425 => to_unsigned(1040, 12), 426 => to_unsigned(2154, 12), 427 => to_unsigned(164, 12), 428 => to_unsigned(606, 12), 429 => to_unsigned(3608, 12), 430 => to_unsigned(2676, 12), 431 => to_unsigned(1215, 12), 432 => to_unsigned(1219, 12), 433 => to_unsigned(1331, 12), 434 => to_unsigned(136, 12), 435 => to_unsigned(952, 12), 436 => to_unsigned(859, 12), 437 => to_unsigned(3165, 12), 438 => to_unsigned(1915, 12), 439 => to_unsigned(2798, 12), 440 => to_unsigned(1111, 12), 441 => to_unsigned(160, 12), 442 => to_unsigned(2195, 12), 443 => to_unsigned(584, 12), 444 => to_unsigned(2503, 12), 445 => to_unsigned(1111, 12), 446 => to_unsigned(3085, 12), 447 => to_unsigned(3386, 12), 448 => to_unsigned(1617, 12), 449 => to_unsigned(1144, 12), 450 => to_unsigned(1908, 12), 451 => to_unsigned(2999, 12), 452 => to_unsigned(2880, 12), 453 => to_unsigned(2763, 12), 454 => to_unsigned(732, 12), 455 => to_unsigned(932, 12), 456 => to_unsigned(281, 12), 457 => to_unsigned(800, 12), 458 => to_unsigned(3498, 12), 459 => to_unsigned(3854, 12), 460 => to_unsigned(470, 12), 461 => to_unsigned(1308, 12), 462 => to_unsigned(3348, 12), 463 => to_unsigned(4050, 12), 464 => to_unsigned(3396, 12), 465 => to_unsigned(1558, 12), 466 => to_unsigned(1251, 12), 467 => to_unsigned(2938, 12), 468 => to_unsigned(595, 12), 469 => to_unsigned(647, 12), 470 => to_unsigned(4040, 12), 471 => to_unsigned(573, 12), 472 => to_unsigned(2701, 12), 473 => to_unsigned(1541, 12), 474 => to_unsigned(256, 12), 475 => to_unsigned(3208, 12), 476 => to_unsigned(3279, 12), 477 => to_unsigned(2511, 12), 478 => to_unsigned(4021, 12), 479 => to_unsigned(1163, 12), 480 => to_unsigned(1028, 12), 481 => to_unsigned(2471, 12), 482 => to_unsigned(348, 12), 483 => to_unsigned(2989, 12), 484 => to_unsigned(1306, 12), 485 => to_unsigned(586, 12), 486 => to_unsigned(1844, 12), 487 => to_unsigned(1006, 12), 488 => to_unsigned(3505, 12), 489 => to_unsigned(3291, 12), 490 => to_unsigned(2867, 12), 491 => to_unsigned(739, 12), 492 => to_unsigned(873, 12), 493 => to_unsigned(786, 12), 494 => to_unsigned(3445, 12), 495 => to_unsigned(1314, 12), 496 => to_unsigned(3635, 12), 497 => to_unsigned(3742, 12), 498 => to_unsigned(437, 12), 499 => to_unsigned(3898, 12), 500 => to_unsigned(4011, 12), 501 => to_unsigned(1847, 12), 502 => to_unsigned(1532, 12), 503 => to_unsigned(1020, 12), 504 => to_unsigned(2834, 12), 505 => to_unsigned(941, 12), 506 => to_unsigned(2903, 12), 507 => to_unsigned(449, 12), 508 => to_unsigned(3398, 12), 509 => to_unsigned(1514, 12), 510 => to_unsigned(3125, 12), 511 => to_unsigned(816, 12), 512 => to_unsigned(3166, 12), 513 => to_unsigned(2107, 12), 514 => to_unsigned(2384, 12), 515 => to_unsigned(1690, 12), 516 => to_unsigned(1660, 12), 517 => to_unsigned(163, 12), 518 => to_unsigned(3642, 12), 519 => to_unsigned(945, 12), 520 => to_unsigned(1130, 12), 521 => to_unsigned(201, 12), 522 => to_unsigned(3372, 12), 523 => to_unsigned(1805, 12), 524 => to_unsigned(2937, 12), 525 => to_unsigned(1862, 12), 526 => to_unsigned(550, 12), 527 => to_unsigned(3751, 12), 528 => to_unsigned(1672, 12), 529 => to_unsigned(3085, 12), 530 => to_unsigned(2040, 12), 531 => to_unsigned(903, 12), 532 => to_unsigned(1744, 12), 533 => to_unsigned(3064, 12), 534 => to_unsigned(2582, 12), 535 => to_unsigned(504, 12), 536 => to_unsigned(3919, 12), 537 => to_unsigned(2009, 12), 538 => to_unsigned(1800, 12), 539 => to_unsigned(3811, 12), 540 => to_unsigned(3846, 12), 541 => to_unsigned(3281, 12), 542 => to_unsigned(1479, 12), 543 => to_unsigned(2516, 12), 544 => to_unsigned(1497, 12), 545 => to_unsigned(4034, 12), 546 => to_unsigned(1596, 12), 547 => to_unsigned(400, 12), 548 => to_unsigned(3128, 12), 549 => to_unsigned(2930, 12), 550 => to_unsigned(3821, 12), 551 => to_unsigned(2711, 12), 552 => to_unsigned(280, 12), 553 => to_unsigned(1028, 12), 554 => to_unsigned(2660, 12), 555 => to_unsigned(1004, 12), 556 => to_unsigned(2353, 12), 557 => to_unsigned(2391, 12), 558 => to_unsigned(1566, 12), 559 => to_unsigned(3638, 12), 560 => to_unsigned(153, 12), 561 => to_unsigned(3860, 12), 562 => to_unsigned(3425, 12), 563 => to_unsigned(2405, 12), 564 => to_unsigned(2745, 12), 565 => to_unsigned(407, 12), 566 => to_unsigned(3483, 12), 567 => to_unsigned(1053, 12), 568 => to_unsigned(2977, 12), 569 => to_unsigned(1395, 12), 570 => to_unsigned(3893, 12), 571 => to_unsigned(2679, 12), 572 => to_unsigned(2995, 12), 573 => to_unsigned(854, 12), 574 => to_unsigned(2550, 12), 575 => to_unsigned(7, 12), 576 => to_unsigned(2665, 12), 577 => to_unsigned(3057, 12), 578 => to_unsigned(2185, 12), 579 => to_unsigned(2742, 12), 580 => to_unsigned(3968, 12), 581 => to_unsigned(851, 12), 582 => to_unsigned(1400, 12), 583 => to_unsigned(932, 12), 584 => to_unsigned(3793, 12), 585 => to_unsigned(3220, 12), 586 => to_unsigned(3957, 12), 587 => to_unsigned(3056, 12), 588 => to_unsigned(3331, 12), 589 => to_unsigned(126, 12), 590 => to_unsigned(1834, 12), 591 => to_unsigned(577, 12), 592 => to_unsigned(1556, 12), 593 => to_unsigned(804, 12), 594 => to_unsigned(1348, 12), 595 => to_unsigned(3024, 12), 596 => to_unsigned(112, 12), 597 => to_unsigned(1967, 12), 598 => to_unsigned(650, 12), 599 => to_unsigned(237, 12), 600 => to_unsigned(1384, 12), 601 => to_unsigned(990, 12), 602 => to_unsigned(1883, 12), 603 => to_unsigned(1579, 12), 604 => to_unsigned(63, 12), 605 => to_unsigned(3999, 12), 606 => to_unsigned(3988, 12), 607 => to_unsigned(2502, 12), 608 => to_unsigned(1289, 12), 609 => to_unsigned(3516, 12), 610 => to_unsigned(603, 12), 611 => to_unsigned(2671, 12), 612 => to_unsigned(1443, 12), 613 => to_unsigned(2387, 12), 614 => to_unsigned(1868, 12), 615 => to_unsigned(1298, 12), 616 => to_unsigned(3441, 12), 617 => to_unsigned(3914, 12), 618 => to_unsigned(2274, 12), 619 => to_unsigned(1249, 12), 620 => to_unsigned(1963, 12), 621 => to_unsigned(1667, 12), 622 => to_unsigned(2956, 12), 623 => to_unsigned(3300, 12), 624 => to_unsigned(3898, 12), 625 => to_unsigned(3969, 12), 626 => to_unsigned(2417, 12), 627 => to_unsigned(3200, 12), 628 => to_unsigned(807, 12), 629 => to_unsigned(1048, 12), 630 => to_unsigned(698, 12), 631 => to_unsigned(292, 12), 632 => to_unsigned(2403, 12), 633 => to_unsigned(837, 12), 634 => to_unsigned(2182, 12), 635 => to_unsigned(3, 12), 636 => to_unsigned(1250, 12), 637 => to_unsigned(2937, 12), 638 => to_unsigned(680, 12), 639 => to_unsigned(2492, 12), 640 => to_unsigned(1441, 12), 641 => to_unsigned(3356, 12), 642 => to_unsigned(2884, 12), 643 => to_unsigned(26, 12), 644 => to_unsigned(736, 12), 645 => to_unsigned(2296, 12), 646 => to_unsigned(365, 12), 647 => to_unsigned(1971, 12), 648 => to_unsigned(3273, 12), 649 => to_unsigned(1461, 12), 650 => to_unsigned(197, 12), 651 => to_unsigned(929, 12), 652 => to_unsigned(1671, 12), 653 => to_unsigned(2685, 12), 654 => to_unsigned(606, 12), 655 => to_unsigned(2120, 12), 656 => to_unsigned(246, 12), 657 => to_unsigned(2900, 12), 658 => to_unsigned(1159, 12), 659 => to_unsigned(1731, 12), 660 => to_unsigned(2261, 12), 661 => to_unsigned(3547, 12), 662 => to_unsigned(3692, 12), 663 => to_unsigned(3395, 12), 664 => to_unsigned(2150, 12), 665 => to_unsigned(3924, 12), 666 => to_unsigned(2375, 12), 667 => to_unsigned(595, 12), 668 => to_unsigned(1247, 12), 669 => to_unsigned(2304, 12), 670 => to_unsigned(3717, 12), 671 => to_unsigned(3419, 12), 672 => to_unsigned(1131, 12), 673 => to_unsigned(2974, 12), 674 => to_unsigned(1993, 12), 675 => to_unsigned(2003, 12), 676 => to_unsigned(3591, 12), 677 => to_unsigned(3221, 12), 678 => to_unsigned(2021, 12), 679 => to_unsigned(3548, 12), 680 => to_unsigned(1416, 12), 681 => to_unsigned(1707, 12), 682 => to_unsigned(1582, 12), 683 => to_unsigned(0, 12), 684 => to_unsigned(3432, 12), 685 => to_unsigned(691, 12), 686 => to_unsigned(1574, 12), 687 => to_unsigned(1113, 12), 688 => to_unsigned(3146, 12), 689 => to_unsigned(2547, 12), 690 => to_unsigned(2786, 12), 691 => to_unsigned(2683, 12), 692 => to_unsigned(343, 12), 693 => to_unsigned(3168, 12), 694 => to_unsigned(2899, 12), 695 => to_unsigned(282, 12), 696 => to_unsigned(2766, 12), 697 => to_unsigned(2080, 12), 698 => to_unsigned(3187, 12), 699 => to_unsigned(2502, 12), 700 => to_unsigned(1889, 12), 701 => to_unsigned(428, 12), 702 => to_unsigned(827, 12), 703 => to_unsigned(1849, 12), 704 => to_unsigned(2738, 12), 705 => to_unsigned(2221, 12), 706 => to_unsigned(1769, 12), 707 => to_unsigned(3204, 12), 708 => to_unsigned(3513, 12), 709 => to_unsigned(93, 12), 710 => to_unsigned(3419, 12), 711 => to_unsigned(1425, 12), 712 => to_unsigned(2467, 12), 713 => to_unsigned(3778, 12), 714 => to_unsigned(404, 12), 715 => to_unsigned(941, 12), 716 => to_unsigned(1209, 12), 717 => to_unsigned(975, 12), 718 => to_unsigned(375, 12), 719 => to_unsigned(3748, 12), 720 => to_unsigned(3945, 12), 721 => to_unsigned(2750, 12), 722 => to_unsigned(3588, 12), 723 => to_unsigned(497, 12), 724 => to_unsigned(3570, 12), 725 => to_unsigned(3277, 12), 726 => to_unsigned(1438, 12), 727 => to_unsigned(1389, 12), 728 => to_unsigned(1879, 12), 729 => to_unsigned(738, 12), 730 => to_unsigned(419, 12), 731 => to_unsigned(2633, 12), 732 => to_unsigned(3290, 12), 733 => to_unsigned(1975, 12), 734 => to_unsigned(1562, 12), 735 => to_unsigned(1398, 12), 736 => to_unsigned(1046, 12), 737 => to_unsigned(460, 12), 738 => to_unsigned(2767, 12), 739 => to_unsigned(3426, 12), 740 => to_unsigned(3674, 12), 741 => to_unsigned(3123, 12), 742 => to_unsigned(3046, 12), 743 => to_unsigned(1838, 12), 744 => to_unsigned(3792, 12), 745 => to_unsigned(3645, 12), 746 => to_unsigned(1468, 12), 747 => to_unsigned(2863, 12), 748 => to_unsigned(2042, 12), 749 => to_unsigned(2152, 12), 750 => to_unsigned(640, 12), 751 => to_unsigned(3466, 12), 752 => to_unsigned(4043, 12), 753 => to_unsigned(1933, 12), 754 => to_unsigned(327, 12), 755 => to_unsigned(606, 12), 756 => to_unsigned(1542, 12), 757 => to_unsigned(3757, 12), 758 => to_unsigned(3317, 12), 759 => to_unsigned(1438, 12), 760 => to_unsigned(1551, 12), 761 => to_unsigned(2217, 12), 762 => to_unsigned(2214, 12), 763 => to_unsigned(1333, 12), 764 => to_unsigned(2987, 12), 765 => to_unsigned(594, 12), 766 => to_unsigned(3463, 12), 767 => to_unsigned(3292, 12), 768 => to_unsigned(2881, 12), 769 => to_unsigned(1705, 12), 770 => to_unsigned(2882, 12), 771 => to_unsigned(3186, 12), 772 => to_unsigned(2908, 12), 773 => to_unsigned(334, 12), 774 => to_unsigned(741, 12), 775 => to_unsigned(1243, 12), 776 => to_unsigned(3318, 12), 777 => to_unsigned(100, 12), 778 => to_unsigned(2463, 12), 779 => to_unsigned(2269, 12), 780 => to_unsigned(1202, 12), 781 => to_unsigned(3580, 12), 782 => to_unsigned(174, 12), 783 => to_unsigned(605, 12), 784 => to_unsigned(3698, 12), 785 => to_unsigned(3745, 12), 786 => to_unsigned(780, 12), 787 => to_unsigned(3808, 12), 788 => to_unsigned(1769, 12), 789 => to_unsigned(848, 12), 790 => to_unsigned(1090, 12), 791 => to_unsigned(1480, 12), 792 => to_unsigned(1011, 12), 793 => to_unsigned(2173, 12), 794 => to_unsigned(1162, 12), 795 => to_unsigned(624, 12), 796 => to_unsigned(2778, 12), 797 => to_unsigned(1179, 12), 798 => to_unsigned(696, 12), 799 => to_unsigned(3192, 12), 800 => to_unsigned(321, 12), 801 => to_unsigned(2496, 12), 802 => to_unsigned(2757, 12), 803 => to_unsigned(3928, 12), 804 => to_unsigned(3362, 12), 805 => to_unsigned(4047, 12), 806 => to_unsigned(2051, 12), 807 => to_unsigned(2748, 12), 808 => to_unsigned(3310, 12), 809 => to_unsigned(3749, 12), 810 => to_unsigned(3243, 12), 811 => to_unsigned(1747, 12), 812 => to_unsigned(2904, 12), 813 => to_unsigned(3654, 12), 814 => to_unsigned(3732, 12), 815 => to_unsigned(902, 12), 816 => to_unsigned(3868, 12), 817 => to_unsigned(627, 12), 818 => to_unsigned(902, 12), 819 => to_unsigned(834, 12), 820 => to_unsigned(604, 12), 821 => to_unsigned(4060, 12), 822 => to_unsigned(3686, 12), 823 => to_unsigned(869, 12), 824 => to_unsigned(3451, 12), 825 => to_unsigned(3781, 12), 826 => to_unsigned(1133, 12), 827 => to_unsigned(1353, 12), 828 => to_unsigned(100, 12), 829 => to_unsigned(694, 12), 830 => to_unsigned(845, 12), 831 => to_unsigned(1941, 12), 832 => to_unsigned(1531, 12), 833 => to_unsigned(671, 12), 834 => to_unsigned(3665, 12), 835 => to_unsigned(3107, 12), 836 => to_unsigned(237, 12), 837 => to_unsigned(3315, 12), 838 => to_unsigned(2298, 12), 839 => to_unsigned(2440, 12), 840 => to_unsigned(2814, 12), 841 => to_unsigned(1305, 12), 842 => to_unsigned(21, 12), 843 => to_unsigned(2477, 12), 844 => to_unsigned(1253, 12), 845 => to_unsigned(2006, 12), 846 => to_unsigned(400, 12), 847 => to_unsigned(1177, 12), 848 => to_unsigned(1006, 12), 849 => to_unsigned(3191, 12), 850 => to_unsigned(1701, 12), 851 => to_unsigned(3967, 12), 852 => to_unsigned(1409, 12), 853 => to_unsigned(1413, 12), 854 => to_unsigned(1734, 12), 855 => to_unsigned(2444, 12), 856 => to_unsigned(3418, 12), 857 => to_unsigned(586, 12), 858 => to_unsigned(3067, 12), 859 => to_unsigned(950, 12), 860 => to_unsigned(3150, 12), 861 => to_unsigned(830, 12), 862 => to_unsigned(1608, 12), 863 => to_unsigned(2247, 12), 864 => to_unsigned(3885, 12), 865 => to_unsigned(3205, 12), 866 => to_unsigned(3631, 12), 867 => to_unsigned(699, 12), 868 => to_unsigned(1194, 12), 869 => to_unsigned(451, 12), 870 => to_unsigned(2186, 12), 871 => to_unsigned(754, 12), 872 => to_unsigned(1337, 12), 873 => to_unsigned(3547, 12), 874 => to_unsigned(1369, 12), 875 => to_unsigned(387, 12), 876 => to_unsigned(1149, 12), 877 => to_unsigned(2766, 12), 878 => to_unsigned(3922, 12), 879 => to_unsigned(1221, 12), 880 => to_unsigned(1722, 12), 881 => to_unsigned(1924, 12), 882 => to_unsigned(3089, 12), 883 => to_unsigned(709, 12), 884 => to_unsigned(447, 12), 885 => to_unsigned(350, 12), 886 => to_unsigned(664, 12), 887 => to_unsigned(3715, 12), 888 => to_unsigned(325, 12), 889 => to_unsigned(424, 12), 890 => to_unsigned(164, 12), 891 => to_unsigned(3642, 12), 892 => to_unsigned(1201, 12), 893 => to_unsigned(3511, 12), 894 => to_unsigned(2712, 12), 895 => to_unsigned(673, 12), 896 => to_unsigned(1938, 12), 897 => to_unsigned(3937, 12), 898 => to_unsigned(462, 12), 899 => to_unsigned(753, 12), 900 => to_unsigned(3207, 12), 901 => to_unsigned(1973, 12), 902 => to_unsigned(747, 12), 903 => to_unsigned(46, 12), 904 => to_unsigned(3568, 12), 905 => to_unsigned(3060, 12), 906 => to_unsigned(2687, 12), 907 => to_unsigned(2977, 12), 908 => to_unsigned(337, 12), 909 => to_unsigned(1181, 12), 910 => to_unsigned(3596, 12), 911 => to_unsigned(3702, 12), 912 => to_unsigned(1838, 12), 913 => to_unsigned(2934, 12), 914 => to_unsigned(288, 12), 915 => to_unsigned(3874, 12), 916 => to_unsigned(115, 12), 917 => to_unsigned(1623, 12), 918 => to_unsigned(2684, 12), 919 => to_unsigned(409, 12), 920 => to_unsigned(3246, 12), 921 => to_unsigned(2546, 12), 922 => to_unsigned(3947, 12), 923 => to_unsigned(3636, 12), 924 => to_unsigned(4073, 12), 925 => to_unsigned(622, 12), 926 => to_unsigned(1600, 12), 927 => to_unsigned(3404, 12), 928 => to_unsigned(3958, 12), 929 => to_unsigned(2633, 12), 930 => to_unsigned(146, 12), 931 => to_unsigned(2820, 12), 932 => to_unsigned(1799, 12), 933 => to_unsigned(2691, 12), 934 => to_unsigned(1072, 12), 935 => to_unsigned(3148, 12), 936 => to_unsigned(2341, 12), 937 => to_unsigned(116, 12), 938 => to_unsigned(1517, 12), 939 => to_unsigned(1584, 12), 940 => to_unsigned(2157, 12), 941 => to_unsigned(2002, 12), 942 => to_unsigned(2227, 12), 943 => to_unsigned(2609, 12), 944 => to_unsigned(3143, 12), 945 => to_unsigned(3930, 12), 946 => to_unsigned(3505, 12), 947 => to_unsigned(4078, 12), 948 => to_unsigned(1309, 12), 949 => to_unsigned(515, 12), 950 => to_unsigned(74, 12), 951 => to_unsigned(3668, 12), 952 => to_unsigned(2538, 12), 953 => to_unsigned(3393, 12), 954 => to_unsigned(1911, 12), 955 => to_unsigned(3604, 12), 956 => to_unsigned(3280, 12), 957 => to_unsigned(1066, 12), 958 => to_unsigned(1522, 12), 959 => to_unsigned(28, 12), 960 => to_unsigned(1434, 12), 961 => to_unsigned(2903, 12), 962 => to_unsigned(3252, 12), 963 => to_unsigned(2352, 12), 964 => to_unsigned(1986, 12), 965 => to_unsigned(1638, 12), 966 => to_unsigned(777, 12), 967 => to_unsigned(3330, 12), 968 => to_unsigned(3444, 12), 969 => to_unsigned(2924, 12), 970 => to_unsigned(1769, 12), 971 => to_unsigned(857, 12), 972 => to_unsigned(1404, 12), 973 => to_unsigned(885, 12), 974 => to_unsigned(612, 12), 975 => to_unsigned(90, 12), 976 => to_unsigned(1092, 12), 977 => to_unsigned(617, 12), 978 => to_unsigned(1546, 12), 979 => to_unsigned(12, 12), 980 => to_unsigned(1640, 12), 981 => to_unsigned(2273, 12), 982 => to_unsigned(2469, 12), 983 => to_unsigned(167, 12), 984 => to_unsigned(928, 12), 985 => to_unsigned(1402, 12), 986 => to_unsigned(3361, 12), 987 => to_unsigned(922, 12), 988 => to_unsigned(99, 12), 989 => to_unsigned(3289, 12), 990 => to_unsigned(2354, 12), 991 => to_unsigned(2392, 12), 992 => to_unsigned(3282, 12), 993 => to_unsigned(1812, 12), 994 => to_unsigned(734, 12), 995 => to_unsigned(3740, 12), 996 => to_unsigned(1608, 12), 997 => to_unsigned(1298, 12), 998 => to_unsigned(1433, 12), 999 => to_unsigned(920, 12), 1000 => to_unsigned(3623, 12), 1001 => to_unsigned(3306, 12), 1002 => to_unsigned(1659, 12), 1003 => to_unsigned(284, 12), 1004 => to_unsigned(1688, 12), 1005 => to_unsigned(3730, 12), 1006 => to_unsigned(3779, 12), 1007 => to_unsigned(2220, 12), 1008 => to_unsigned(3795, 12), 1009 => to_unsigned(2349, 12), 1010 => to_unsigned(2870, 12), 1011 => to_unsigned(0, 12), 1012 => to_unsigned(2186, 12), 1013 => to_unsigned(707, 12), 1014 => to_unsigned(1926, 12), 1015 => to_unsigned(1755, 12), 1016 => to_unsigned(1891, 12), 1017 => to_unsigned(2489, 12), 1018 => to_unsigned(4038, 12), 1019 => to_unsigned(2963, 12), 1020 => to_unsigned(1186, 12), 1021 => to_unsigned(2098, 12), 1022 => to_unsigned(2290, 12), 1023 => to_unsigned(870, 12), 1024 => to_unsigned(2068, 12), 1025 => to_unsigned(2731, 12), 1026 => to_unsigned(630, 12), 1027 => to_unsigned(2176, 12), 1028 => to_unsigned(1508, 12), 1029 => to_unsigned(2413, 12), 1030 => to_unsigned(105, 12), 1031 => to_unsigned(3778, 12), 1032 => to_unsigned(225, 12), 1033 => to_unsigned(3724, 12), 1034 => to_unsigned(1807, 12), 1035 => to_unsigned(3190, 12), 1036 => to_unsigned(2593, 12), 1037 => to_unsigned(2199, 12), 1038 => to_unsigned(1932, 12), 1039 => to_unsigned(3973, 12), 1040 => to_unsigned(3110, 12), 1041 => to_unsigned(3841, 12), 1042 => to_unsigned(266, 12), 1043 => to_unsigned(3078, 12), 1044 => to_unsigned(3965, 12), 1045 => to_unsigned(1286, 12), 1046 => to_unsigned(614, 12), 1047 => to_unsigned(4006, 12), 1048 => to_unsigned(331, 12), 1049 => to_unsigned(1394, 12), 1050 => to_unsigned(1365, 12), 1051 => to_unsigned(3454, 12), 1052 => to_unsigned(2418, 12), 1053 => to_unsigned(2738, 12), 1054 => to_unsigned(3891, 12), 1055 => to_unsigned(3330, 12), 1056 => to_unsigned(3404, 12), 1057 => to_unsigned(669, 12), 1058 => to_unsigned(1545, 12), 1059 => to_unsigned(627, 12), 1060 => to_unsigned(968, 12), 1061 => to_unsigned(389, 12), 1062 => to_unsigned(2676, 12), 1063 => to_unsigned(181, 12), 1064 => to_unsigned(2283, 12), 1065 => to_unsigned(193, 12), 1066 => to_unsigned(3883, 12), 1067 => to_unsigned(2639, 12), 1068 => to_unsigned(3134, 12), 1069 => to_unsigned(2380, 12), 1070 => to_unsigned(2607, 12), 1071 => to_unsigned(2636, 12), 1072 => to_unsigned(1685, 12), 1073 => to_unsigned(120, 12), 1074 => to_unsigned(1810, 12), 1075 => to_unsigned(2393, 12), 1076 => to_unsigned(525, 12), 1077 => to_unsigned(222, 12), 1078 => to_unsigned(3676, 12), 1079 => to_unsigned(236, 12), 1080 => to_unsigned(2153, 12), 1081 => to_unsigned(3285, 12), 1082 => to_unsigned(3590, 12), 1083 => to_unsigned(612, 12), 1084 => to_unsigned(3632, 12), 1085 => to_unsigned(1576, 12), 1086 => to_unsigned(922, 12), 1087 => to_unsigned(3230, 12), 1088 => to_unsigned(3461, 12), 1089 => to_unsigned(2191, 12), 1090 => to_unsigned(959, 12), 1091 => to_unsigned(3557, 12), 1092 => to_unsigned(3109, 12), 1093 => to_unsigned(3643, 12), 1094 => to_unsigned(3697, 12), 1095 => to_unsigned(95, 12), 1096 => to_unsigned(2400, 12), 1097 => to_unsigned(2544, 12), 1098 => to_unsigned(2256, 12), 1099 => to_unsigned(2336, 12), 1100 => to_unsigned(62, 12), 1101 => to_unsigned(2442, 12), 1102 => to_unsigned(2444, 12), 1103 => to_unsigned(1629, 12), 1104 => to_unsigned(3904, 12), 1105 => to_unsigned(1437, 12), 1106 => to_unsigned(2394, 12), 1107 => to_unsigned(2023, 12), 1108 => to_unsigned(150, 12), 1109 => to_unsigned(403, 12), 1110 => to_unsigned(2437, 12), 1111 => to_unsigned(2852, 12), 1112 => to_unsigned(595, 12), 1113 => to_unsigned(127, 12), 1114 => to_unsigned(1508, 12), 1115 => to_unsigned(1797, 12), 1116 => to_unsigned(3420, 12), 1117 => to_unsigned(2508, 12), 1118 => to_unsigned(3226, 12), 1119 => to_unsigned(3825, 12), 1120 => to_unsigned(1107, 12), 1121 => to_unsigned(3980, 12), 1122 => to_unsigned(2022, 12), 1123 => to_unsigned(1159, 12), 1124 => to_unsigned(3252, 12), 1125 => to_unsigned(592, 12), 1126 => to_unsigned(2461, 12), 1127 => to_unsigned(1024, 12), 1128 => to_unsigned(3799, 12), 1129 => to_unsigned(2767, 12), 1130 => to_unsigned(3914, 12), 1131 => to_unsigned(3836, 12), 1132 => to_unsigned(3715, 12), 1133 => to_unsigned(573, 12), 1134 => to_unsigned(2371, 12), 1135 => to_unsigned(3216, 12), 1136 => to_unsigned(1904, 12), 1137 => to_unsigned(1481, 12), 1138 => to_unsigned(3668, 12), 1139 => to_unsigned(116, 12), 1140 => to_unsigned(741, 12), 1141 => to_unsigned(3839, 12), 1142 => to_unsigned(824, 12), 1143 => to_unsigned(1342, 12), 1144 => to_unsigned(3000, 12), 1145 => to_unsigned(2608, 12), 1146 => to_unsigned(1169, 12), 1147 => to_unsigned(1909, 12), 1148 => to_unsigned(4025, 12), 1149 => to_unsigned(3593, 12), 1150 => to_unsigned(492, 12), 1151 => to_unsigned(1214, 12), 1152 => to_unsigned(2127, 12), 1153 => to_unsigned(742, 12), 1154 => to_unsigned(3278, 12), 1155 => to_unsigned(417, 12), 1156 => to_unsigned(1924, 12), 1157 => to_unsigned(2960, 12), 1158 => to_unsigned(2276, 12), 1159 => to_unsigned(1863, 12), 1160 => to_unsigned(3390, 12), 1161 => to_unsigned(3863, 12), 1162 => to_unsigned(3931, 12), 1163 => to_unsigned(2414, 12), 1164 => to_unsigned(7, 12), 1165 => to_unsigned(2557, 12), 1166 => to_unsigned(790, 12), 1167 => to_unsigned(1890, 12), 1168 => to_unsigned(2206, 12), 1169 => to_unsigned(1782, 12), 1170 => to_unsigned(1616, 12), 1171 => to_unsigned(1179, 12), 1172 => to_unsigned(3631, 12), 1173 => to_unsigned(495, 12), 1174 => to_unsigned(626, 12), 1175 => to_unsigned(2571, 12), 1176 => to_unsigned(2007, 12), 1177 => to_unsigned(1870, 12), 1178 => to_unsigned(4071, 12), 1179 => to_unsigned(798, 12), 1180 => to_unsigned(2138, 12), 1181 => to_unsigned(2338, 12), 1182 => to_unsigned(2614, 12), 1183 => to_unsigned(1873, 12), 1184 => to_unsigned(2723, 12), 1185 => to_unsigned(3143, 12), 1186 => to_unsigned(2925, 12), 1187 => to_unsigned(3899, 12), 1188 => to_unsigned(624, 12), 1189 => to_unsigned(421, 12), 1190 => to_unsigned(1092, 12), 1191 => to_unsigned(437, 12), 1192 => to_unsigned(3085, 12), 1193 => to_unsigned(2149, 12), 1194 => to_unsigned(787, 12), 1195 => to_unsigned(3947, 12), 1196 => to_unsigned(3336, 12), 1197 => to_unsigned(2912, 12), 1198 => to_unsigned(1745, 12), 1199 => to_unsigned(1221, 12), 1200 => to_unsigned(2428, 12), 1201 => to_unsigned(100, 12), 1202 => to_unsigned(1409, 12), 1203 => to_unsigned(765, 12), 1204 => to_unsigned(1181, 12), 1205 => to_unsigned(901, 12), 1206 => to_unsigned(4048, 12), 1207 => to_unsigned(230, 12), 1208 => to_unsigned(504, 12), 1209 => to_unsigned(1960, 12), 1210 => to_unsigned(2710, 12), 1211 => to_unsigned(3102, 12), 1212 => to_unsigned(2303, 12), 1213 => to_unsigned(2579, 12), 1214 => to_unsigned(1796, 12), 1215 => to_unsigned(660, 12), 1216 => to_unsigned(2922, 12), 1217 => to_unsigned(2634, 12), 1218 => to_unsigned(123, 12), 1219 => to_unsigned(3523, 12), 1220 => to_unsigned(3286, 12), 1221 => to_unsigned(2364, 12), 1222 => to_unsigned(2789, 12), 1223 => to_unsigned(1274, 12), 1224 => to_unsigned(1629, 12), 1225 => to_unsigned(681, 12), 1226 => to_unsigned(1576, 12), 1227 => to_unsigned(2236, 12), 1228 => to_unsigned(1233, 12), 1229 => to_unsigned(691, 12), 1230 => to_unsigned(1320, 12), 1231 => to_unsigned(2107, 12), 1232 => to_unsigned(2538, 12), 1233 => to_unsigned(1502, 12), 1234 => to_unsigned(2589, 12), 1235 => to_unsigned(2273, 12), 1236 => to_unsigned(3678, 12), 1237 => to_unsigned(3310, 12), 1238 => to_unsigned(3749, 12), 1239 => to_unsigned(382, 12), 1240 => to_unsigned(2264, 12), 1241 => to_unsigned(3344, 12), 1242 => to_unsigned(2915, 12), 1243 => to_unsigned(3239, 12), 1244 => to_unsigned(3741, 12), 1245 => to_unsigned(508, 12), 1246 => to_unsigned(3137, 12), 1247 => to_unsigned(3863, 12), 1248 => to_unsigned(3272, 12), 1249 => to_unsigned(1408, 12), 1250 => to_unsigned(1111, 12), 1251 => to_unsigned(3877, 12), 1252 => to_unsigned(1391, 12), 1253 => to_unsigned(2495, 12), 1254 => to_unsigned(2458, 12), 1255 => to_unsigned(729, 12), 1256 => to_unsigned(1369, 12), 1257 => to_unsigned(3206, 12), 1258 => to_unsigned(2264, 12), 1259 => to_unsigned(1527, 12), 1260 => to_unsigned(2511, 12), 1261 => to_unsigned(1125, 12), 1262 => to_unsigned(1321, 12), 1263 => to_unsigned(1937, 12), 1264 => to_unsigned(4048, 12), 1265 => to_unsigned(3952, 12), 1266 => to_unsigned(3115, 12), 1267 => to_unsigned(1134, 12), 1268 => to_unsigned(3525, 12), 1269 => to_unsigned(374, 12), 1270 => to_unsigned(2963, 12), 1271 => to_unsigned(2799, 12), 1272 => to_unsigned(1814, 12), 1273 => to_unsigned(3437, 12), 1274 => to_unsigned(3979, 12), 1275 => to_unsigned(2571, 12), 1276 => to_unsigned(2977, 12), 1277 => to_unsigned(3975, 12), 1278 => to_unsigned(2167, 12), 1279 => to_unsigned(282, 12), 1280 => to_unsigned(560, 12), 1281 => to_unsigned(3271, 12), 1282 => to_unsigned(239, 12), 1283 => to_unsigned(2742, 12), 1284 => to_unsigned(608, 12), 1285 => to_unsigned(356, 12), 1286 => to_unsigned(1874, 12), 1287 => to_unsigned(2647, 12), 1288 => to_unsigned(1429, 12), 1289 => to_unsigned(1534, 12), 1290 => to_unsigned(2562, 12), 1291 => to_unsigned(3336, 12), 1292 => to_unsigned(3338, 12), 1293 => to_unsigned(2309, 12), 1294 => to_unsigned(3366, 12), 1295 => to_unsigned(2982, 12), 1296 => to_unsigned(612, 12), 1297 => to_unsigned(449, 12), 1298 => to_unsigned(1653, 12), 1299 => to_unsigned(571, 12), 1300 => to_unsigned(3748, 12), 1301 => to_unsigned(901, 12), 1302 => to_unsigned(2309, 12), 1303 => to_unsigned(2086, 12), 1304 => to_unsigned(3747, 12), 1305 => to_unsigned(2136, 12), 1306 => to_unsigned(4017, 12), 1307 => to_unsigned(1743, 12), 1308 => to_unsigned(3412, 12), 1309 => to_unsigned(2418, 12), 1310 => to_unsigned(1289, 12), 1311 => to_unsigned(4087, 12), 1312 => to_unsigned(3204, 12), 1313 => to_unsigned(2993, 12), 1314 => to_unsigned(3096, 12), 1315 => to_unsigned(1630, 12), 1316 => to_unsigned(3458, 12), 1317 => to_unsigned(3923, 12), 1318 => to_unsigned(3971, 12), 1319 => to_unsigned(3661, 12), 1320 => to_unsigned(1291, 12), 1321 => to_unsigned(397, 12), 1322 => to_unsigned(2532, 12), 1323 => to_unsigned(2129, 12), 1324 => to_unsigned(1178, 12), 1325 => to_unsigned(4038, 12), 1326 => to_unsigned(1711, 12), 1327 => to_unsigned(1634, 12), 1328 => to_unsigned(1557, 12), 1329 => to_unsigned(3988, 12), 1330 => to_unsigned(1706, 12), 1331 => to_unsigned(3962, 12), 1332 => to_unsigned(2489, 12), 1333 => to_unsigned(1169, 12), 1334 => to_unsigned(613, 12), 1335 => to_unsigned(4057, 12), 1336 => to_unsigned(3316, 12), 1337 => to_unsigned(2517, 12), 1338 => to_unsigned(183, 12), 1339 => to_unsigned(3684, 12), 1340 => to_unsigned(3268, 12), 1341 => to_unsigned(111, 12), 1342 => to_unsigned(1250, 12), 1343 => to_unsigned(2827, 12), 1344 => to_unsigned(4066, 12), 1345 => to_unsigned(2145, 12), 1346 => to_unsigned(2286, 12), 1347 => to_unsigned(2451, 12), 1348 => to_unsigned(3952, 12), 1349 => to_unsigned(1035, 12), 1350 => to_unsigned(3041, 12), 1351 => to_unsigned(1561, 12), 1352 => to_unsigned(1121, 12), 1353 => to_unsigned(1375, 12), 1354 => to_unsigned(2349, 12), 1355 => to_unsigned(2822, 12), 1356 => to_unsigned(2649, 12), 1357 => to_unsigned(3928, 12), 1358 => to_unsigned(2541, 12), 1359 => to_unsigned(2598, 12), 1360 => to_unsigned(51, 12), 1361 => to_unsigned(1040, 12), 1362 => to_unsigned(3991, 12), 1363 => to_unsigned(3802, 12), 1364 => to_unsigned(771, 12), 1365 => to_unsigned(1882, 12), 1366 => to_unsigned(430, 12), 1367 => to_unsigned(3706, 12), 1368 => to_unsigned(1437, 12), 1369 => to_unsigned(770, 12), 1370 => to_unsigned(645, 12), 1371 => to_unsigned(1401, 12), 1372 => to_unsigned(4039, 12), 1373 => to_unsigned(2831, 12), 1374 => to_unsigned(2894, 12), 1375 => to_unsigned(1443, 12), 1376 => to_unsigned(2228, 12), 1377 => to_unsigned(1383, 12), 1378 => to_unsigned(3958, 12), 1379 => to_unsigned(2311, 12), 1380 => to_unsigned(2739, 12), 1381 => to_unsigned(3430, 12), 1382 => to_unsigned(761, 12), 1383 => to_unsigned(947, 12), 1384 => to_unsigned(3997, 12), 1385 => to_unsigned(695, 12), 1386 => to_unsigned(625, 12), 1387 => to_unsigned(395, 12), 1388 => to_unsigned(2499, 12), 1389 => to_unsigned(1741, 12), 1390 => to_unsigned(3962, 12), 1391 => to_unsigned(3383, 12), 1392 => to_unsigned(3672, 12), 1393 => to_unsigned(2555, 12), 1394 => to_unsigned(3324, 12), 1395 => to_unsigned(504, 12), 1396 => to_unsigned(1860, 12), 1397 => to_unsigned(3189, 12), 1398 => to_unsigned(2419, 12), 1399 => to_unsigned(3542, 12), 1400 => to_unsigned(1209, 12), 1401 => to_unsigned(2397, 12), 1402 => to_unsigned(2662, 12), 1403 => to_unsigned(907, 12), 1404 => to_unsigned(3790, 12), 1405 => to_unsigned(3666, 12), 1406 => to_unsigned(4057, 12), 1407 => to_unsigned(3308, 12), 1408 => to_unsigned(3, 12), 1409 => to_unsigned(165, 12), 1410 => to_unsigned(1415, 12), 1411 => to_unsigned(1821, 12), 1412 => to_unsigned(1102, 12), 1413 => to_unsigned(3851, 12), 1414 => to_unsigned(3017, 12), 1415 => to_unsigned(523, 12), 1416 => to_unsigned(2832, 12), 1417 => to_unsigned(3132, 12), 1418 => to_unsigned(2683, 12), 1419 => to_unsigned(103, 12), 1420 => to_unsigned(1727, 12), 1421 => to_unsigned(699, 12), 1422 => to_unsigned(2177, 12), 1423 => to_unsigned(1938, 12), 1424 => to_unsigned(3765, 12), 1425 => to_unsigned(1308, 12), 1426 => to_unsigned(448, 12), 1427 => to_unsigned(853, 12), 1428 => to_unsigned(3800, 12), 1429 => to_unsigned(1609, 12), 1430 => to_unsigned(2952, 12), 1431 => to_unsigned(4050, 12), 1432 => to_unsigned(3467, 12), 1433 => to_unsigned(2524, 12), 1434 => to_unsigned(2421, 12), 1435 => to_unsigned(1971, 12), 1436 => to_unsigned(2897, 12), 1437 => to_unsigned(439, 12), 1438 => to_unsigned(3087, 12), 1439 => to_unsigned(131, 12), 1440 => to_unsigned(1130, 12), 1441 => to_unsigned(2520, 12), 1442 => to_unsigned(213, 12), 1443 => to_unsigned(3356, 12), 1444 => to_unsigned(3898, 12), 1445 => to_unsigned(3797, 12), 1446 => to_unsigned(1614, 12), 1447 => to_unsigned(2927, 12), 1448 => to_unsigned(833, 12), 1449 => to_unsigned(844, 12), 1450 => to_unsigned(1291, 12), 1451 => to_unsigned(1305, 12), 1452 => to_unsigned(1383, 12), 1453 => to_unsigned(1803, 12), 1454 => to_unsigned(858, 12), 1455 => to_unsigned(749, 12), 1456 => to_unsigned(1442, 12), 1457 => to_unsigned(1921, 12), 1458 => to_unsigned(3070, 12), 1459 => to_unsigned(656, 12), 1460 => to_unsigned(3329, 12), 1461 => to_unsigned(2576, 12), 1462 => to_unsigned(2593, 12), 1463 => to_unsigned(3105, 12), 1464 => to_unsigned(3244, 12), 1465 => to_unsigned(1510, 12), 1466 => to_unsigned(808, 12), 1467 => to_unsigned(2376, 12), 1468 => to_unsigned(2253, 12), 1469 => to_unsigned(1130, 12), 1470 => to_unsigned(595, 12), 1471 => to_unsigned(754, 12), 1472 => to_unsigned(1440, 12), 1473 => to_unsigned(919, 12), 1474 => to_unsigned(324, 12), 1475 => to_unsigned(1439, 12), 1476 => to_unsigned(662, 12), 1477 => to_unsigned(3136, 12), 1478 => to_unsigned(3813, 12), 1479 => to_unsigned(3359, 12), 1480 => to_unsigned(79, 12), 1481 => to_unsigned(83, 12), 1482 => to_unsigned(2831, 12), 1483 => to_unsigned(2867, 12), 1484 => to_unsigned(3577, 12), 1485 => to_unsigned(3468, 12), 1486 => to_unsigned(2733, 12), 1487 => to_unsigned(1034, 12), 1488 => to_unsigned(1524, 12), 1489 => to_unsigned(1641, 12), 1490 => to_unsigned(848, 12), 1491 => to_unsigned(3142, 12), 1492 => to_unsigned(2069, 12), 1493 => to_unsigned(3806, 12), 1494 => to_unsigned(1731, 12), 1495 => to_unsigned(1360, 12), 1496 => to_unsigned(1344, 12), 1497 => to_unsigned(1153, 12), 1498 => to_unsigned(1842, 12), 1499 => to_unsigned(2912, 12), 1500 => to_unsigned(363, 12), 1501 => to_unsigned(1019, 12), 1502 => to_unsigned(466, 12), 1503 => to_unsigned(2386, 12), 1504 => to_unsigned(697, 12), 1505 => to_unsigned(3478, 12), 1506 => to_unsigned(3855, 12), 1507 => to_unsigned(911, 12), 1508 => to_unsigned(3612, 12), 1509 => to_unsigned(3399, 12), 1510 => to_unsigned(1307, 12), 1511 => to_unsigned(2264, 12), 1512 => to_unsigned(313, 12), 1513 => to_unsigned(2874, 12), 1514 => to_unsigned(2264, 12), 1515 => to_unsigned(1996, 12), 1516 => to_unsigned(2317, 12), 1517 => to_unsigned(1938, 12), 1518 => to_unsigned(78, 12), 1519 => to_unsigned(4046, 12), 1520 => to_unsigned(1812, 12), 1521 => to_unsigned(1607, 12), 1522 => to_unsigned(1719, 12), 1523 => to_unsigned(3372, 12), 1524 => to_unsigned(2283, 12), 1525 => to_unsigned(3317, 12), 1526 => to_unsigned(3163, 12), 1527 => to_unsigned(2092, 12), 1528 => to_unsigned(3855, 12), 1529 => to_unsigned(2045, 12), 1530 => to_unsigned(1623, 12), 1531 => to_unsigned(1995, 12), 1532 => to_unsigned(1613, 12), 1533 => to_unsigned(510, 12), 1534 => to_unsigned(3485, 12), 1535 => to_unsigned(1631, 12), 1536 => to_unsigned(110, 12), 1537 => to_unsigned(3794, 12), 1538 => to_unsigned(3716, 12), 1539 => to_unsigned(540, 12), 1540 => to_unsigned(1729, 12), 1541 => to_unsigned(2097, 12), 1542 => to_unsigned(945, 12), 1543 => to_unsigned(2391, 12), 1544 => to_unsigned(3641, 12), 1545 => to_unsigned(3792, 12), 1546 => to_unsigned(3113, 12), 1547 => to_unsigned(1498, 12), 1548 => to_unsigned(1776, 12), 1549 => to_unsigned(1218, 12), 1550 => to_unsigned(2991, 12), 1551 => to_unsigned(2321, 12), 1552 => to_unsigned(3092, 12), 1553 => to_unsigned(2726, 12), 1554 => to_unsigned(1344, 12), 1555 => to_unsigned(3718, 12), 1556 => to_unsigned(236, 12), 1557 => to_unsigned(662, 12), 1558 => to_unsigned(2127, 12), 1559 => to_unsigned(2122, 12), 1560 => to_unsigned(1186, 12), 1561 => to_unsigned(3752, 12), 1562 => to_unsigned(2726, 12), 1563 => to_unsigned(3062, 12), 1564 => to_unsigned(1685, 12), 1565 => to_unsigned(3874, 12), 1566 => to_unsigned(373, 12), 1567 => to_unsigned(3232, 12), 1568 => to_unsigned(2474, 12), 1569 => to_unsigned(1407, 12), 1570 => to_unsigned(3372, 12), 1571 => to_unsigned(611, 12), 1572 => to_unsigned(1833, 12), 1573 => to_unsigned(2809, 12), 1574 => to_unsigned(2919, 12), 1575 => to_unsigned(3995, 12), 1576 => to_unsigned(1787, 12), 1577 => to_unsigned(2352, 12), 1578 => to_unsigned(1407, 12), 1579 => to_unsigned(1674, 12), 1580 => to_unsigned(1348, 12), 1581 => to_unsigned(1297, 12), 1582 => to_unsigned(2819, 12), 1583 => to_unsigned(3685, 12), 1584 => to_unsigned(1630, 12), 1585 => to_unsigned(471, 12), 1586 => to_unsigned(2333, 12), 1587 => to_unsigned(614, 12), 1588 => to_unsigned(1659, 12), 1589 => to_unsigned(3230, 12), 1590 => to_unsigned(1227, 12), 1591 => to_unsigned(450, 12), 1592 => to_unsigned(3549, 12), 1593 => to_unsigned(3388, 12), 1594 => to_unsigned(2695, 12), 1595 => to_unsigned(2739, 12), 1596 => to_unsigned(2292, 12), 1597 => to_unsigned(2633, 12), 1598 => to_unsigned(3543, 12), 1599 => to_unsigned(1984, 12), 1600 => to_unsigned(2032, 12), 1601 => to_unsigned(401, 12), 1602 => to_unsigned(1704, 12), 1603 => to_unsigned(243, 12), 1604 => to_unsigned(2581, 12), 1605 => to_unsigned(1630, 12), 1606 => to_unsigned(1946, 12), 1607 => to_unsigned(3215, 12), 1608 => to_unsigned(2800, 12), 1609 => to_unsigned(1809, 12), 1610 => to_unsigned(2314, 12), 1611 => to_unsigned(1681, 12), 1612 => to_unsigned(2179, 12), 1613 => to_unsigned(3047, 12), 1614 => to_unsigned(3657, 12), 1615 => to_unsigned(797, 12), 1616 => to_unsigned(3267, 12), 1617 => to_unsigned(2503, 12), 1618 => to_unsigned(464, 12), 1619 => to_unsigned(2274, 12), 1620 => to_unsigned(3716, 12), 1621 => to_unsigned(445, 12), 1622 => to_unsigned(1882, 12), 1623 => to_unsigned(1124, 12), 1624 => to_unsigned(2182, 12), 1625 => to_unsigned(32, 12), 1626 => to_unsigned(3153, 12), 1627 => to_unsigned(1655, 12), 1628 => to_unsigned(2422, 12), 1629 => to_unsigned(1781, 12), 1630 => to_unsigned(2341, 12), 1631 => to_unsigned(2679, 12), 1632 => to_unsigned(1307, 12), 1633 => to_unsigned(1075, 12), 1634 => to_unsigned(1614, 12), 1635 => to_unsigned(4027, 12), 1636 => to_unsigned(1622, 12), 1637 => to_unsigned(1631, 12), 1638 => to_unsigned(2056, 12), 1639 => to_unsigned(3384, 12), 1640 => to_unsigned(2845, 12), 1641 => to_unsigned(2716, 12), 1642 => to_unsigned(2015, 12), 1643 => to_unsigned(1442, 12), 1644 => to_unsigned(186, 12), 1645 => to_unsigned(1919, 12), 1646 => to_unsigned(3966, 12), 1647 => to_unsigned(4049, 12), 1648 => to_unsigned(1500, 12), 1649 => to_unsigned(2159, 12), 1650 => to_unsigned(3728, 12), 1651 => to_unsigned(4040, 12), 1652 => to_unsigned(1595, 12), 1653 => to_unsigned(247, 12), 1654 => to_unsigned(1004, 12), 1655 => to_unsigned(1031, 12), 1656 => to_unsigned(2956, 12), 1657 => to_unsigned(1312, 12), 1658 => to_unsigned(3796, 12), 1659 => to_unsigned(747, 12), 1660 => to_unsigned(75, 12), 1661 => to_unsigned(3293, 12), 1662 => to_unsigned(1064, 12), 1663 => to_unsigned(1024, 12), 1664 => to_unsigned(212, 12), 1665 => to_unsigned(1133, 12), 1666 => to_unsigned(2652, 12), 1667 => to_unsigned(3277, 12), 1668 => to_unsigned(1189, 12), 1669 => to_unsigned(2479, 12), 1670 => to_unsigned(573, 12), 1671 => to_unsigned(103, 12), 1672 => to_unsigned(1970, 12), 1673 => to_unsigned(580, 12), 1674 => to_unsigned(494, 12), 1675 => to_unsigned(3020, 12), 1676 => to_unsigned(3769, 12), 1677 => to_unsigned(887, 12), 1678 => to_unsigned(4069, 12), 1679 => to_unsigned(4080, 12), 1680 => to_unsigned(1156, 12), 1681 => to_unsigned(2665, 12), 1682 => to_unsigned(2596, 12), 1683 => to_unsigned(336, 12), 1684 => to_unsigned(2514, 12), 1685 => to_unsigned(165, 12), 1686 => to_unsigned(734, 12), 1687 => to_unsigned(373, 12), 1688 => to_unsigned(1518, 12), 1689 => to_unsigned(3363, 12), 1690 => to_unsigned(1968, 12), 1691 => to_unsigned(1664, 12), 1692 => to_unsigned(1585, 12), 1693 => to_unsigned(3257, 12), 1694 => to_unsigned(265, 12), 1695 => to_unsigned(2098, 12), 1696 => to_unsigned(2785, 12), 1697 => to_unsigned(1200, 12), 1698 => to_unsigned(4081, 12), 1699 => to_unsigned(524, 12), 1700 => to_unsigned(3782, 12), 1701 => to_unsigned(3708, 12), 1702 => to_unsigned(2547, 12), 1703 => to_unsigned(1956, 12), 1704 => to_unsigned(1123, 12), 1705 => to_unsigned(358, 12), 1706 => to_unsigned(1060, 12), 1707 => to_unsigned(3358, 12), 1708 => to_unsigned(1650, 12), 1709 => to_unsigned(3219, 12), 1710 => to_unsigned(3494, 12), 1711 => to_unsigned(428, 12), 1712 => to_unsigned(35, 12), 1713 => to_unsigned(782, 12), 1714 => to_unsigned(2077, 12), 1715 => to_unsigned(4019, 12), 1716 => to_unsigned(60, 12), 1717 => to_unsigned(1016, 12), 1718 => to_unsigned(3409, 12), 1719 => to_unsigned(2883, 12), 1720 => to_unsigned(1821, 12), 1721 => to_unsigned(155, 12), 1722 => to_unsigned(3203, 12), 1723 => to_unsigned(1057, 12), 1724 => to_unsigned(3829, 12), 1725 => to_unsigned(435, 12), 1726 => to_unsigned(3958, 12), 1727 => to_unsigned(1435, 12), 1728 => to_unsigned(3300, 12), 1729 => to_unsigned(56, 12), 1730 => to_unsigned(2325, 12), 1731 => to_unsigned(679, 12), 1732 => to_unsigned(3818, 12), 1733 => to_unsigned(3402, 12), 1734 => to_unsigned(2589, 12), 1735 => to_unsigned(2289, 12), 1736 => to_unsigned(2973, 12), 1737 => to_unsigned(957, 12), 1738 => to_unsigned(1594, 12), 1739 => to_unsigned(1816, 12), 1740 => to_unsigned(114, 12), 1741 => to_unsigned(3344, 12), 1742 => to_unsigned(2496, 12), 1743 => to_unsigned(3940, 12), 1744 => to_unsigned(2018, 12), 1745 => to_unsigned(2683, 12), 1746 => to_unsigned(2061, 12), 1747 => to_unsigned(769, 12), 1748 => to_unsigned(3835, 12), 1749 => to_unsigned(258, 12), 1750 => to_unsigned(1858, 12), 1751 => to_unsigned(2195, 12), 1752 => to_unsigned(2548, 12), 1753 => to_unsigned(3834, 12), 1754 => to_unsigned(1484, 12), 1755 => to_unsigned(3742, 12), 1756 => to_unsigned(1575, 12), 1757 => to_unsigned(3541, 12), 1758 => to_unsigned(1613, 12), 1759 => to_unsigned(2993, 12), 1760 => to_unsigned(1306, 12), 1761 => to_unsigned(371, 12), 1762 => to_unsigned(1164, 12), 1763 => to_unsigned(3313, 12), 1764 => to_unsigned(960, 12), 1765 => to_unsigned(2305, 12), 1766 => to_unsigned(3492, 12), 1767 => to_unsigned(3850, 12), 1768 => to_unsigned(3946, 12), 1769 => to_unsigned(2336, 12), 1770 => to_unsigned(1534, 12), 1771 => to_unsigned(3356, 12), 1772 => to_unsigned(2746, 12), 1773 => to_unsigned(2754, 12), 1774 => to_unsigned(2780, 12), 1775 => to_unsigned(1089, 12), 1776 => to_unsigned(1229, 12), 1777 => to_unsigned(2387, 12), 1778 => to_unsigned(2607, 12), 1779 => to_unsigned(2641, 12), 1780 => to_unsigned(420, 12), 1781 => to_unsigned(3271, 12), 1782 => to_unsigned(1333, 12), 1783 => to_unsigned(1734, 12), 1784 => to_unsigned(649, 12), 1785 => to_unsigned(3599, 12), 1786 => to_unsigned(2834, 12), 1787 => to_unsigned(1181, 12), 1788 => to_unsigned(693, 12), 1789 => to_unsigned(3004, 12), 1790 => to_unsigned(554, 12), 1791 => to_unsigned(2514, 12), 1792 => to_unsigned(2690, 12), 1793 => to_unsigned(2845, 12), 1794 => to_unsigned(2449, 12), 1795 => to_unsigned(2083, 12), 1796 => to_unsigned(2936, 12), 1797 => to_unsigned(3347, 12), 1798 => to_unsigned(3984, 12), 1799 => to_unsigned(3607, 12), 1800 => to_unsigned(3724, 12), 1801 => to_unsigned(355, 12), 1802 => to_unsigned(2925, 12), 1803 => to_unsigned(1720, 12), 1804 => to_unsigned(1730, 12), 1805 => to_unsigned(2836, 12), 1806 => to_unsigned(3203, 12), 1807 => to_unsigned(81, 12), 1808 => to_unsigned(2988, 12), 1809 => to_unsigned(2086, 12), 1810 => to_unsigned(3114, 12), 1811 => to_unsigned(3018, 12), 1812 => to_unsigned(549, 12), 1813 => to_unsigned(362, 12), 1814 => to_unsigned(552, 12), 1815 => to_unsigned(1903, 12), 1816 => to_unsigned(3867, 12), 1817 => to_unsigned(1668, 12), 1818 => to_unsigned(1459, 12), 1819 => to_unsigned(2454, 12), 1820 => to_unsigned(2725, 12), 1821 => to_unsigned(2851, 12), 1822 => to_unsigned(542, 12), 1823 => to_unsigned(1799, 12), 1824 => to_unsigned(3032, 12), 1825 => to_unsigned(1624, 12), 1826 => to_unsigned(239, 12), 1827 => to_unsigned(1935, 12), 1828 => to_unsigned(2442, 12), 1829 => to_unsigned(3219, 12), 1830 => to_unsigned(2893, 12), 1831 => to_unsigned(2023, 12), 1832 => to_unsigned(1848, 12), 1833 => to_unsigned(2021, 12), 1834 => to_unsigned(4071, 12), 1835 => to_unsigned(1938, 12), 1836 => to_unsigned(3527, 12), 1837 => to_unsigned(60, 12), 1838 => to_unsigned(24, 12), 1839 => to_unsigned(160, 12), 1840 => to_unsigned(3436, 12), 1841 => to_unsigned(3367, 12), 1842 => to_unsigned(2932, 12), 1843 => to_unsigned(3176, 12), 1844 => to_unsigned(1406, 12), 1845 => to_unsigned(367, 12), 1846 => to_unsigned(116, 12), 1847 => to_unsigned(2020, 12), 1848 => to_unsigned(2026, 12), 1849 => to_unsigned(16, 12), 1850 => to_unsigned(948, 12), 1851 => to_unsigned(2266, 12), 1852 => to_unsigned(4072, 12), 1853 => to_unsigned(2256, 12), 1854 => to_unsigned(814, 12), 1855 => to_unsigned(3296, 12), 1856 => to_unsigned(2654, 12), 1857 => to_unsigned(1876, 12), 1858 => to_unsigned(3863, 12), 1859 => to_unsigned(3727, 12), 1860 => to_unsigned(172, 12), 1861 => to_unsigned(2643, 12), 1862 => to_unsigned(1143, 12), 1863 => to_unsigned(1591, 12), 1864 => to_unsigned(1378, 12), 1865 => to_unsigned(3483, 12), 1866 => to_unsigned(2349, 12), 1867 => to_unsigned(3042, 12), 1868 => to_unsigned(1361, 12), 1869 => to_unsigned(3799, 12), 1870 => to_unsigned(3483, 12), 1871 => to_unsigned(3661, 12), 1872 => to_unsigned(432, 12), 1873 => to_unsigned(2007, 12), 1874 => to_unsigned(2910, 12), 1875 => to_unsigned(1413, 12), 1876 => to_unsigned(377, 12), 1877 => to_unsigned(231, 12), 1878 => to_unsigned(737, 12), 1879 => to_unsigned(881, 12), 1880 => to_unsigned(994, 12), 1881 => to_unsigned(1820, 12), 1882 => to_unsigned(3316, 12), 1883 => to_unsigned(3137, 12), 1884 => to_unsigned(2116, 12), 1885 => to_unsigned(2773, 12), 1886 => to_unsigned(2504, 12), 1887 => to_unsigned(1788, 12), 1888 => to_unsigned(370, 12), 1889 => to_unsigned(2977, 12), 1890 => to_unsigned(1398, 12), 1891 => to_unsigned(3555, 12), 1892 => to_unsigned(1584, 12), 1893 => to_unsigned(1123, 12), 1894 => to_unsigned(4057, 12), 1895 => to_unsigned(1605, 12), 1896 => to_unsigned(1985, 12), 1897 => to_unsigned(1635, 12), 1898 => to_unsigned(2119, 12), 1899 => to_unsigned(2561, 12), 1900 => to_unsigned(129, 12), 1901 => to_unsigned(199, 12), 1902 => to_unsigned(3737, 12), 1903 => to_unsigned(1124, 12), 1904 => to_unsigned(2637, 12), 1905 => to_unsigned(3692, 12), 1906 => to_unsigned(3250, 12), 1907 => to_unsigned(1435, 12), 1908 => to_unsigned(96, 12), 1909 => to_unsigned(1579, 12), 1910 => to_unsigned(3859, 12), 1911 => to_unsigned(2402, 12), 1912 => to_unsigned(1325, 12), 1913 => to_unsigned(100, 12), 1914 => to_unsigned(336, 12), 1915 => to_unsigned(112, 12), 1916 => to_unsigned(3306, 12), 1917 => to_unsigned(889, 12), 1918 => to_unsigned(2987, 12), 1919 => to_unsigned(3523, 12), 1920 => to_unsigned(2568, 12), 1921 => to_unsigned(2259, 12), 1922 => to_unsigned(2990, 12), 1923 => to_unsigned(2624, 12), 1924 => to_unsigned(372, 12), 1925 => to_unsigned(3988, 12), 1926 => to_unsigned(3168, 12), 1927 => to_unsigned(1506, 12), 1928 => to_unsigned(875, 12), 1929 => to_unsigned(2437, 12), 1930 => to_unsigned(341, 12), 1931 => to_unsigned(2328, 12), 1932 => to_unsigned(1026, 12), 1933 => to_unsigned(2557, 12), 1934 => to_unsigned(3069, 12), 1935 => to_unsigned(3527, 12), 1936 => to_unsigned(1132, 12), 1937 => to_unsigned(2251, 12), 1938 => to_unsigned(243, 12), 1939 => to_unsigned(3868, 12), 1940 => to_unsigned(374, 12), 1941 => to_unsigned(863, 12), 1942 => to_unsigned(65, 12), 1943 => to_unsigned(2512, 12), 1944 => to_unsigned(2418, 12), 1945 => to_unsigned(210, 12), 1946 => to_unsigned(3470, 12), 1947 => to_unsigned(3605, 12), 1948 => to_unsigned(1135, 12), 1949 => to_unsigned(1903, 12), 1950 => to_unsigned(2245, 12), 1951 => to_unsigned(801, 12), 1952 => to_unsigned(3690, 12), 1953 => to_unsigned(1154, 12), 1954 => to_unsigned(539, 12), 1955 => to_unsigned(2792, 12), 1956 => to_unsigned(375, 12), 1957 => to_unsigned(3219, 12), 1958 => to_unsigned(3983, 12), 1959 => to_unsigned(839, 12), 1960 => to_unsigned(2028, 12), 1961 => to_unsigned(2845, 12), 1962 => to_unsigned(1443, 12), 1963 => to_unsigned(2785, 12), 1964 => to_unsigned(2352, 12), 1965 => to_unsigned(945, 12), 1966 => to_unsigned(848, 12), 1967 => to_unsigned(184, 12), 1968 => to_unsigned(319, 12), 1969 => to_unsigned(3544, 12), 1970 => to_unsigned(1466, 12), 1971 => to_unsigned(901, 12), 1972 => to_unsigned(1843, 12), 1973 => to_unsigned(1274, 12), 1974 => to_unsigned(573, 12), 1975 => to_unsigned(3178, 12), 1976 => to_unsigned(2515, 12), 1977 => to_unsigned(3345, 12), 1978 => to_unsigned(2093, 12), 1979 => to_unsigned(992, 12), 1980 => to_unsigned(1598, 12), 1981 => to_unsigned(3094, 12), 1982 => to_unsigned(1249, 12), 1983 => to_unsigned(3686, 12), 1984 => to_unsigned(3721, 12), 1985 => to_unsigned(2821, 12), 1986 => to_unsigned(1356, 12), 1987 => to_unsigned(1597, 12), 1988 => to_unsigned(2218, 12), 1989 => to_unsigned(759, 12), 1990 => to_unsigned(400, 12), 1991 => to_unsigned(3387, 12), 1992 => to_unsigned(273, 12), 1993 => to_unsigned(3268, 12), 1994 => to_unsigned(1340, 12), 1995 => to_unsigned(1689, 12), 1996 => to_unsigned(1166, 12), 1997 => to_unsigned(877, 12), 1998 => to_unsigned(3901, 12), 1999 => to_unsigned(181, 12), 2000 => to_unsigned(81, 12), 2001 => to_unsigned(3613, 12), 2002 => to_unsigned(2246, 12), 2003 => to_unsigned(28, 12), 2004 => to_unsigned(3786, 12), 2005 => to_unsigned(3717, 12), 2006 => to_unsigned(2532, 12), 2007 => to_unsigned(484, 12), 2008 => to_unsigned(2388, 12), 2009 => to_unsigned(4023, 12), 2010 => to_unsigned(498, 12), 2011 => to_unsigned(178, 12), 2012 => to_unsigned(3670, 12), 2013 => to_unsigned(2229, 12), 2014 => to_unsigned(1802, 12), 2015 => to_unsigned(3627, 12), 2016 => to_unsigned(3003, 12), 2017 => to_unsigned(1438, 12), 2018 => to_unsigned(1851, 12), 2019 => to_unsigned(1166, 12), 2020 => to_unsigned(2035, 12), 2021 => to_unsigned(1456, 12), 2022 => to_unsigned(632, 12), 2023 => to_unsigned(1405, 12), 2024 => to_unsigned(1080, 12), 2025 => to_unsigned(449, 12), 2026 => to_unsigned(1896, 12), 2027 => to_unsigned(3975, 12), 2028 => to_unsigned(3013, 12), 2029 => to_unsigned(2191, 12), 2030 => to_unsigned(631, 12), 2031 => to_unsigned(3049, 12), 2032 => to_unsigned(2356, 12), 2033 => to_unsigned(2336, 12), 2034 => to_unsigned(3159, 12), 2035 => to_unsigned(1998, 12), 2036 => to_unsigned(2978, 12), 2037 => to_unsigned(1565, 12), 2038 => to_unsigned(2099, 12), 2039 => to_unsigned(3545, 12), 2040 => to_unsigned(437, 12), 2041 => to_unsigned(2820, 12), 2042 => to_unsigned(1216, 12), 2043 => to_unsigned(3963, 12), 2044 => to_unsigned(2202, 12), 2045 => to_unsigned(1492, 12), 2046 => to_unsigned(2437, 12), 2047 => to_unsigned(2426, 12)),
            1 => (0 => to_unsigned(2904, 12), 1 => to_unsigned(2321, 12), 2 => to_unsigned(1988, 12), 3 => to_unsigned(2360, 12), 4 => to_unsigned(2208, 12), 5 => to_unsigned(1265, 12), 6 => to_unsigned(337, 12), 7 => to_unsigned(1608, 12), 8 => to_unsigned(73, 12), 9 => to_unsigned(740, 12), 10 => to_unsigned(1439, 12), 11 => to_unsigned(2398, 12), 12 => to_unsigned(3401, 12), 13 => to_unsigned(364, 12), 14 => to_unsigned(3248, 12), 15 => to_unsigned(739, 12), 16 => to_unsigned(1440, 12), 17 => to_unsigned(1294, 12), 18 => to_unsigned(573, 12), 19 => to_unsigned(3415, 12), 20 => to_unsigned(416, 12), 21 => to_unsigned(2360, 12), 22 => to_unsigned(412, 12), 23 => to_unsigned(171, 12), 24 => to_unsigned(1121, 12), 25 => to_unsigned(178, 12), 26 => to_unsigned(2862, 12), 27 => to_unsigned(2156, 12), 28 => to_unsigned(1864, 12), 29 => to_unsigned(2469, 12), 30 => to_unsigned(2680, 12), 31 => to_unsigned(2050, 12), 32 => to_unsigned(785, 12), 33 => to_unsigned(143, 12), 34 => to_unsigned(707, 12), 35 => to_unsigned(1365, 12), 36 => to_unsigned(1520, 12), 37 => to_unsigned(754, 12), 38 => to_unsigned(3165, 12), 39 => to_unsigned(1893, 12), 40 => to_unsigned(3192, 12), 41 => to_unsigned(2710, 12), 42 => to_unsigned(1234, 12), 43 => to_unsigned(3591, 12), 44 => to_unsigned(823, 12), 45 => to_unsigned(2225, 12), 46 => to_unsigned(1050, 12), 47 => to_unsigned(760, 12), 48 => to_unsigned(644, 12), 49 => to_unsigned(3181, 12), 50 => to_unsigned(89, 12), 51 => to_unsigned(1050, 12), 52 => to_unsigned(3772, 12), 53 => to_unsigned(2291, 12), 54 => to_unsigned(3695, 12), 55 => to_unsigned(1619, 12), 56 => to_unsigned(2638, 12), 57 => to_unsigned(658, 12), 58 => to_unsigned(3193, 12), 59 => to_unsigned(2656, 12), 60 => to_unsigned(2395, 12), 61 => to_unsigned(2852, 12), 62 => to_unsigned(3430, 12), 63 => to_unsigned(3476, 12), 64 => to_unsigned(1407, 12), 65 => to_unsigned(1516, 12), 66 => to_unsigned(387, 12), 67 => to_unsigned(1682, 12), 68 => to_unsigned(205, 12), 69 => to_unsigned(2099, 12), 70 => to_unsigned(561, 12), 71 => to_unsigned(3615, 12), 72 => to_unsigned(2529, 12), 73 => to_unsigned(1682, 12), 74 => to_unsigned(2316, 12), 75 => to_unsigned(2671, 12), 76 => to_unsigned(4059, 12), 77 => to_unsigned(2279, 12), 78 => to_unsigned(2914, 12), 79 => to_unsigned(3911, 12), 80 => to_unsigned(3678, 12), 81 => to_unsigned(2861, 12), 82 => to_unsigned(3792, 12), 83 => to_unsigned(2113, 12), 84 => to_unsigned(2136, 12), 85 => to_unsigned(2320, 12), 86 => to_unsigned(2349, 12), 87 => to_unsigned(2431, 12), 88 => to_unsigned(2267, 12), 89 => to_unsigned(165, 12), 90 => to_unsigned(434, 12), 91 => to_unsigned(2456, 12), 92 => to_unsigned(1968, 12), 93 => to_unsigned(1228, 12), 94 => to_unsigned(1028, 12), 95 => to_unsigned(1008, 12), 96 => to_unsigned(947, 12), 97 => to_unsigned(1198, 12), 98 => to_unsigned(3112, 12), 99 => to_unsigned(3982, 12), 100 => to_unsigned(3313, 12), 101 => to_unsigned(2442, 12), 102 => to_unsigned(3483, 12), 103 => to_unsigned(3406, 12), 104 => to_unsigned(870, 12), 105 => to_unsigned(1421, 12), 106 => to_unsigned(3588, 12), 107 => to_unsigned(726, 12), 108 => to_unsigned(1295, 12), 109 => to_unsigned(3101, 12), 110 => to_unsigned(974, 12), 111 => to_unsigned(3242, 12), 112 => to_unsigned(3737, 12), 113 => to_unsigned(1227, 12), 114 => to_unsigned(479, 12), 115 => to_unsigned(3291, 12), 116 => to_unsigned(2582, 12), 117 => to_unsigned(3182, 12), 118 => to_unsigned(811, 12), 119 => to_unsigned(1492, 12), 120 => to_unsigned(3767, 12), 121 => to_unsigned(2813, 12), 122 => to_unsigned(1154, 12), 123 => to_unsigned(3737, 12), 124 => to_unsigned(1661, 12), 125 => to_unsigned(2168, 12), 126 => to_unsigned(1664, 12), 127 => to_unsigned(3423, 12), 128 => to_unsigned(184, 12), 129 => to_unsigned(3182, 12), 130 => to_unsigned(3782, 12), 131 => to_unsigned(978, 12), 132 => to_unsigned(2646, 12), 133 => to_unsigned(2238, 12), 134 => to_unsigned(3839, 12), 135 => to_unsigned(3630, 12), 136 => to_unsigned(763, 12), 137 => to_unsigned(1113, 12), 138 => to_unsigned(2765, 12), 139 => to_unsigned(1676, 12), 140 => to_unsigned(2366, 12), 141 => to_unsigned(293, 12), 142 => to_unsigned(4051, 12), 143 => to_unsigned(2207, 12), 144 => to_unsigned(887, 12), 145 => to_unsigned(3996, 12), 146 => to_unsigned(2363, 12), 147 => to_unsigned(1528, 12), 148 => to_unsigned(339, 12), 149 => to_unsigned(3880, 12), 150 => to_unsigned(1384, 12), 151 => to_unsigned(1401, 12), 152 => to_unsigned(3673, 12), 153 => to_unsigned(4079, 12), 154 => to_unsigned(3869, 12), 155 => to_unsigned(2844, 12), 156 => to_unsigned(1076, 12), 157 => to_unsigned(3370, 12), 158 => to_unsigned(2698, 12), 159 => to_unsigned(3796, 12), 160 => to_unsigned(1297, 12), 161 => to_unsigned(640, 12), 162 => to_unsigned(3751, 12), 163 => to_unsigned(38, 12), 164 => to_unsigned(1506, 12), 165 => to_unsigned(193, 12), 166 => to_unsigned(3632, 12), 167 => to_unsigned(2262, 12), 168 => to_unsigned(3117, 12), 169 => to_unsigned(1146, 12), 170 => to_unsigned(2737, 12), 171 => to_unsigned(1558, 12), 172 => to_unsigned(231, 12), 173 => to_unsigned(1534, 12), 174 => to_unsigned(3420, 12), 175 => to_unsigned(1345, 12), 176 => to_unsigned(1365, 12), 177 => to_unsigned(1858, 12), 178 => to_unsigned(1568, 12), 179 => to_unsigned(2482, 12), 180 => to_unsigned(1350, 12), 181 => to_unsigned(2662, 12), 182 => to_unsigned(2979, 12), 183 => to_unsigned(2037, 12), 184 => to_unsigned(484, 12), 185 => to_unsigned(2199, 12), 186 => to_unsigned(4083, 12), 187 => to_unsigned(2170, 12), 188 => to_unsigned(2130, 12), 189 => to_unsigned(1126, 12), 190 => to_unsigned(89, 12), 191 => to_unsigned(750, 12), 192 => to_unsigned(2127, 12), 193 => to_unsigned(3185, 12), 194 => to_unsigned(155, 12), 195 => to_unsigned(3925, 12), 196 => to_unsigned(1537, 12), 197 => to_unsigned(2313, 12), 198 => to_unsigned(115, 12), 199 => to_unsigned(1873, 12), 200 => to_unsigned(395, 12), 201 => to_unsigned(1088, 12), 202 => to_unsigned(2295, 12), 203 => to_unsigned(1859, 12), 204 => to_unsigned(3577, 12), 205 => to_unsigned(3261, 12), 206 => to_unsigned(54, 12), 207 => to_unsigned(1316, 12), 208 => to_unsigned(2516, 12), 209 => to_unsigned(3198, 12), 210 => to_unsigned(19, 12), 211 => to_unsigned(1007, 12), 212 => to_unsigned(3781, 12), 213 => to_unsigned(724, 12), 214 => to_unsigned(2685, 12), 215 => to_unsigned(3774, 12), 216 => to_unsigned(3268, 12), 217 => to_unsigned(1193, 12), 218 => to_unsigned(208, 12), 219 => to_unsigned(2704, 12), 220 => to_unsigned(2233, 12), 221 => to_unsigned(3717, 12), 222 => to_unsigned(2144, 12), 223 => to_unsigned(2326, 12), 224 => to_unsigned(1155, 12), 225 => to_unsigned(1416, 12), 226 => to_unsigned(830, 12), 227 => to_unsigned(1884, 12), 228 => to_unsigned(1193, 12), 229 => to_unsigned(1866, 12), 230 => to_unsigned(102, 12), 231 => to_unsigned(1628, 12), 232 => to_unsigned(3167, 12), 233 => to_unsigned(2156, 12), 234 => to_unsigned(907, 12), 235 => to_unsigned(930, 12), 236 => to_unsigned(91, 12), 237 => to_unsigned(1841, 12), 238 => to_unsigned(583, 12), 239 => to_unsigned(1447, 12), 240 => to_unsigned(2918, 12), 241 => to_unsigned(2935, 12), 242 => to_unsigned(3130, 12), 243 => to_unsigned(1029, 12), 244 => to_unsigned(1097, 12), 245 => to_unsigned(1880, 12), 246 => to_unsigned(140, 12), 247 => to_unsigned(2792, 12), 248 => to_unsigned(1249, 12), 249 => to_unsigned(3899, 12), 250 => to_unsigned(718, 12), 251 => to_unsigned(2029, 12), 252 => to_unsigned(3599, 12), 253 => to_unsigned(1028, 12), 254 => to_unsigned(1942, 12), 255 => to_unsigned(1716, 12), 256 => to_unsigned(2114, 12), 257 => to_unsigned(3911, 12), 258 => to_unsigned(3437, 12), 259 => to_unsigned(2376, 12), 260 => to_unsigned(3333, 12), 261 => to_unsigned(551, 12), 262 => to_unsigned(335, 12), 263 => to_unsigned(3919, 12), 264 => to_unsigned(3881, 12), 265 => to_unsigned(3033, 12), 266 => to_unsigned(662, 12), 267 => to_unsigned(2521, 12), 268 => to_unsigned(1241, 12), 269 => to_unsigned(915, 12), 270 => to_unsigned(3902, 12), 271 => to_unsigned(797, 12), 272 => to_unsigned(1801, 12), 273 => to_unsigned(3467, 12), 274 => to_unsigned(2941, 12), 275 => to_unsigned(2147, 12), 276 => to_unsigned(3610, 12), 277 => to_unsigned(2919, 12), 278 => to_unsigned(1279, 12), 279 => to_unsigned(3794, 12), 280 => to_unsigned(3656, 12), 281 => to_unsigned(255, 12), 282 => to_unsigned(1665, 12), 283 => to_unsigned(3939, 12), 284 => to_unsigned(2674, 12), 285 => to_unsigned(2289, 12), 286 => to_unsigned(3758, 12), 287 => to_unsigned(1335, 12), 288 => to_unsigned(1546, 12), 289 => to_unsigned(3786, 12), 290 => to_unsigned(1304, 12), 291 => to_unsigned(2559, 12), 292 => to_unsigned(1375, 12), 293 => to_unsigned(1067, 12), 294 => to_unsigned(987, 12), 295 => to_unsigned(1677, 12), 296 => to_unsigned(974, 12), 297 => to_unsigned(55, 12), 298 => to_unsigned(2053, 12), 299 => to_unsigned(407, 12), 300 => to_unsigned(2090, 12), 301 => to_unsigned(1639, 12), 302 => to_unsigned(3121, 12), 303 => to_unsigned(1381, 12), 304 => to_unsigned(870, 12), 305 => to_unsigned(1611, 12), 306 => to_unsigned(1909, 12), 307 => to_unsigned(3000, 12), 308 => to_unsigned(3499, 12), 309 => to_unsigned(152, 12), 310 => to_unsigned(3409, 12), 311 => to_unsigned(1557, 12), 312 => to_unsigned(2014, 12), 313 => to_unsigned(3218, 12), 314 => to_unsigned(63, 12), 315 => to_unsigned(1369, 12), 316 => to_unsigned(1565, 12), 317 => to_unsigned(3365, 12), 318 => to_unsigned(2993, 12), 319 => to_unsigned(1192, 12), 320 => to_unsigned(497, 12), 321 => to_unsigned(2410, 12), 322 => to_unsigned(3295, 12), 323 => to_unsigned(103, 12), 324 => to_unsigned(3339, 12), 325 => to_unsigned(312, 12), 326 => to_unsigned(4085, 12), 327 => to_unsigned(3519, 12), 328 => to_unsigned(2190, 12), 329 => to_unsigned(1312, 12), 330 => to_unsigned(2241, 12), 331 => to_unsigned(1145, 12), 332 => to_unsigned(373, 12), 333 => to_unsigned(833, 12), 334 => to_unsigned(2084, 12), 335 => to_unsigned(1786, 12), 336 => to_unsigned(2073, 12), 337 => to_unsigned(4044, 12), 338 => to_unsigned(2120, 12), 339 => to_unsigned(2098, 12), 340 => to_unsigned(2572, 12), 341 => to_unsigned(2968, 12), 342 => to_unsigned(147, 12), 343 => to_unsigned(1731, 12), 344 => to_unsigned(2442, 12), 345 => to_unsigned(2567, 12), 346 => to_unsigned(948, 12), 347 => to_unsigned(3164, 12), 348 => to_unsigned(3598, 12), 349 => to_unsigned(2504, 12), 350 => to_unsigned(46, 12), 351 => to_unsigned(1251, 12), 352 => to_unsigned(35, 12), 353 => to_unsigned(2257, 12), 354 => to_unsigned(1175, 12), 355 => to_unsigned(2109, 12), 356 => to_unsigned(1653, 12), 357 => to_unsigned(1205, 12), 358 => to_unsigned(524, 12), 359 => to_unsigned(1453, 12), 360 => to_unsigned(3591, 12), 361 => to_unsigned(506, 12), 362 => to_unsigned(1455, 12), 363 => to_unsigned(2158, 12), 364 => to_unsigned(679, 12), 365 => to_unsigned(3934, 12), 366 => to_unsigned(1683, 12), 367 => to_unsigned(1258, 12), 368 => to_unsigned(1901, 12), 369 => to_unsigned(946, 12), 370 => to_unsigned(3649, 12), 371 => to_unsigned(2987, 12), 372 => to_unsigned(594, 12), 373 => to_unsigned(1486, 12), 374 => to_unsigned(2043, 12), 375 => to_unsigned(1113, 12), 376 => to_unsigned(101, 12), 377 => to_unsigned(2424, 12), 378 => to_unsigned(184, 12), 379 => to_unsigned(2632, 12), 380 => to_unsigned(2738, 12), 381 => to_unsigned(2082, 12), 382 => to_unsigned(986, 12), 383 => to_unsigned(523, 12), 384 => to_unsigned(2668, 12), 385 => to_unsigned(3211, 12), 386 => to_unsigned(2408, 12), 387 => to_unsigned(2468, 12), 388 => to_unsigned(3966, 12), 389 => to_unsigned(3249, 12), 390 => to_unsigned(4044, 12), 391 => to_unsigned(2001, 12), 392 => to_unsigned(1247, 12), 393 => to_unsigned(4042, 12), 394 => to_unsigned(1840, 12), 395 => to_unsigned(586, 12), 396 => to_unsigned(3211, 12), 397 => to_unsigned(2653, 12), 398 => to_unsigned(1570, 12), 399 => to_unsigned(714, 12), 400 => to_unsigned(3532, 12), 401 => to_unsigned(2801, 12), 402 => to_unsigned(3367, 12), 403 => to_unsigned(2416, 12), 404 => to_unsigned(1546, 12), 405 => to_unsigned(770, 12), 406 => to_unsigned(1401, 12), 407 => to_unsigned(1007, 12), 408 => to_unsigned(75, 12), 409 => to_unsigned(1966, 12), 410 => to_unsigned(3123, 12), 411 => to_unsigned(2548, 12), 412 => to_unsigned(4009, 12), 413 => to_unsigned(4090, 12), 414 => to_unsigned(3163, 12), 415 => to_unsigned(3715, 12), 416 => to_unsigned(2320, 12), 417 => to_unsigned(3391, 12), 418 => to_unsigned(2880, 12), 419 => to_unsigned(3853, 12), 420 => to_unsigned(3878, 12), 421 => to_unsigned(260, 12), 422 => to_unsigned(2563, 12), 423 => to_unsigned(915, 12), 424 => to_unsigned(593, 12), 425 => to_unsigned(3216, 12), 426 => to_unsigned(2430, 12), 427 => to_unsigned(2887, 12), 428 => to_unsigned(664, 12), 429 => to_unsigned(1291, 12), 430 => to_unsigned(150, 12), 431 => to_unsigned(3644, 12), 432 => to_unsigned(1243, 12), 433 => to_unsigned(642, 12), 434 => to_unsigned(904, 12), 435 => to_unsigned(1096, 12), 436 => to_unsigned(1753, 12), 437 => to_unsigned(2342, 12), 438 => to_unsigned(1588, 12), 439 => to_unsigned(3809, 12), 440 => to_unsigned(2392, 12), 441 => to_unsigned(3391, 12), 442 => to_unsigned(2965, 12), 443 => to_unsigned(2564, 12), 444 => to_unsigned(2463, 12), 445 => to_unsigned(755, 12), 446 => to_unsigned(2251, 12), 447 => to_unsigned(2725, 12), 448 => to_unsigned(1799, 12), 449 => to_unsigned(3734, 12), 450 => to_unsigned(3708, 12), 451 => to_unsigned(1322, 12), 452 => to_unsigned(2235, 12), 453 => to_unsigned(2783, 12), 454 => to_unsigned(310, 12), 455 => to_unsigned(1993, 12), 456 => to_unsigned(3955, 12), 457 => to_unsigned(1459, 12), 458 => to_unsigned(2642, 12), 459 => to_unsigned(3863, 12), 460 => to_unsigned(3155, 12), 461 => to_unsigned(1817, 12), 462 => to_unsigned(1849, 12), 463 => to_unsigned(3269, 12), 464 => to_unsigned(2393, 12), 465 => to_unsigned(301, 12), 466 => to_unsigned(3439, 12), 467 => to_unsigned(1624, 12), 468 => to_unsigned(1971, 12), 469 => to_unsigned(1339, 12), 470 => to_unsigned(1964, 12), 471 => to_unsigned(1178, 12), 472 => to_unsigned(3704, 12), 473 => to_unsigned(2677, 12), 474 => to_unsigned(2987, 12), 475 => to_unsigned(633, 12), 476 => to_unsigned(416, 12), 477 => to_unsigned(1822, 12), 478 => to_unsigned(1678, 12), 479 => to_unsigned(3399, 12), 480 => to_unsigned(96, 12), 481 => to_unsigned(1725, 12), 482 => to_unsigned(513, 12), 483 => to_unsigned(3574, 12), 484 => to_unsigned(2479, 12), 485 => to_unsigned(3452, 12), 486 => to_unsigned(2413, 12), 487 => to_unsigned(3190, 12), 488 => to_unsigned(3243, 12), 489 => to_unsigned(2522, 12), 490 => to_unsigned(1039, 12), 491 => to_unsigned(3908, 12), 492 => to_unsigned(1226, 12), 493 => to_unsigned(2133, 12), 494 => to_unsigned(3751, 12), 495 => to_unsigned(106, 12), 496 => to_unsigned(3563, 12), 497 => to_unsigned(1630, 12), 498 => to_unsigned(3542, 12), 499 => to_unsigned(256, 12), 500 => to_unsigned(1617, 12), 501 => to_unsigned(3258, 12), 502 => to_unsigned(3084, 12), 503 => to_unsigned(1243, 12), 504 => to_unsigned(2859, 12), 505 => to_unsigned(950, 12), 506 => to_unsigned(2429, 12), 507 => to_unsigned(431, 12), 508 => to_unsigned(790, 12), 509 => to_unsigned(2847, 12), 510 => to_unsigned(372, 12), 511 => to_unsigned(3106, 12), 512 => to_unsigned(2018, 12), 513 => to_unsigned(3882, 12), 514 => to_unsigned(3396, 12), 515 => to_unsigned(3962, 12), 516 => to_unsigned(830, 12), 517 => to_unsigned(3876, 12), 518 => to_unsigned(3923, 12), 519 => to_unsigned(2220, 12), 520 => to_unsigned(721, 12), 521 => to_unsigned(2288, 12), 522 => to_unsigned(3439, 12), 523 => to_unsigned(198, 12), 524 => to_unsigned(262, 12), 525 => to_unsigned(3504, 12), 526 => to_unsigned(1417, 12), 527 => to_unsigned(3612, 12), 528 => to_unsigned(77, 12), 529 => to_unsigned(1720, 12), 530 => to_unsigned(2441, 12), 531 => to_unsigned(469, 12), 532 => to_unsigned(1858, 12), 533 => to_unsigned(2569, 12), 534 => to_unsigned(1134, 12), 535 => to_unsigned(3064, 12), 536 => to_unsigned(1188, 12), 537 => to_unsigned(284, 12), 538 => to_unsigned(1524, 12), 539 => to_unsigned(3136, 12), 540 => to_unsigned(970, 12), 541 => to_unsigned(892, 12), 542 => to_unsigned(1165, 12), 543 => to_unsigned(3307, 12), 544 => to_unsigned(1538, 12), 545 => to_unsigned(2469, 12), 546 => to_unsigned(3015, 12), 547 => to_unsigned(3159, 12), 548 => to_unsigned(1758, 12), 549 => to_unsigned(4049, 12), 550 => to_unsigned(1539, 12), 551 => to_unsigned(111, 12), 552 => to_unsigned(2018, 12), 553 => to_unsigned(2896, 12), 554 => to_unsigned(1779, 12), 555 => to_unsigned(594, 12), 556 => to_unsigned(818, 12), 557 => to_unsigned(1981, 12), 558 => to_unsigned(2538, 12), 559 => to_unsigned(978, 12), 560 => to_unsigned(28, 12), 561 => to_unsigned(1827, 12), 562 => to_unsigned(309, 12), 563 => to_unsigned(3866, 12), 564 => to_unsigned(3441, 12), 565 => to_unsigned(1383, 12), 566 => to_unsigned(1578, 12), 567 => to_unsigned(3886, 12), 568 => to_unsigned(197, 12), 569 => to_unsigned(2588, 12), 570 => to_unsigned(127, 12), 571 => to_unsigned(171, 12), 572 => to_unsigned(1107, 12), 573 => to_unsigned(62, 12), 574 => to_unsigned(2890, 12), 575 => to_unsigned(3274, 12), 576 => to_unsigned(2697, 12), 577 => to_unsigned(1243, 12), 578 => to_unsigned(739, 12), 579 => to_unsigned(2891, 12), 580 => to_unsigned(2912, 12), 581 => to_unsigned(166, 12), 582 => to_unsigned(2079, 12), 583 => to_unsigned(3827, 12), 584 => to_unsigned(3990, 12), 585 => to_unsigned(3454, 12), 586 => to_unsigned(1883, 12), 587 => to_unsigned(1849, 12), 588 => to_unsigned(3093, 12), 589 => to_unsigned(3809, 12), 590 => to_unsigned(3901, 12), 591 => to_unsigned(3564, 12), 592 => to_unsigned(3881, 12), 593 => to_unsigned(2419, 12), 594 => to_unsigned(875, 12), 595 => to_unsigned(2403, 12), 596 => to_unsigned(3241, 12), 597 => to_unsigned(2298, 12), 598 => to_unsigned(3735, 12), 599 => to_unsigned(3325, 12), 600 => to_unsigned(2792, 12), 601 => to_unsigned(1844, 12), 602 => to_unsigned(279, 12), 603 => to_unsigned(1146, 12), 604 => to_unsigned(3912, 12), 605 => to_unsigned(3625, 12), 606 => to_unsigned(3309, 12), 607 => to_unsigned(828, 12), 608 => to_unsigned(815, 12), 609 => to_unsigned(1679, 12), 610 => to_unsigned(1060, 12), 611 => to_unsigned(1985, 12), 612 => to_unsigned(2654, 12), 613 => to_unsigned(2021, 12), 614 => to_unsigned(810, 12), 615 => to_unsigned(3838, 12), 616 => to_unsigned(512, 12), 617 => to_unsigned(4051, 12), 618 => to_unsigned(2950, 12), 619 => to_unsigned(733, 12), 620 => to_unsigned(3139, 12), 621 => to_unsigned(287, 12), 622 => to_unsigned(2845, 12), 623 => to_unsigned(2064, 12), 624 => to_unsigned(1987, 12), 625 => to_unsigned(2330, 12), 626 => to_unsigned(4093, 12), 627 => to_unsigned(1286, 12), 628 => to_unsigned(233, 12), 629 => to_unsigned(3557, 12), 630 => to_unsigned(267, 12), 631 => to_unsigned(3409, 12), 632 => to_unsigned(2871, 12), 633 => to_unsigned(893, 12), 634 => to_unsigned(1323, 12), 635 => to_unsigned(2371, 12), 636 => to_unsigned(532, 12), 637 => to_unsigned(475, 12), 638 => to_unsigned(511, 12), 639 => to_unsigned(2679, 12), 640 => to_unsigned(1500, 12), 641 => to_unsigned(270, 12), 642 => to_unsigned(270, 12), 643 => to_unsigned(2128, 12), 644 => to_unsigned(3555, 12), 645 => to_unsigned(447, 12), 646 => to_unsigned(373, 12), 647 => to_unsigned(3814, 12), 648 => to_unsigned(43, 12), 649 => to_unsigned(3227, 12), 650 => to_unsigned(3430, 12), 651 => to_unsigned(3799, 12), 652 => to_unsigned(916, 12), 653 => to_unsigned(1019, 12), 654 => to_unsigned(2583, 12), 655 => to_unsigned(1314, 12), 656 => to_unsigned(3360, 12), 657 => to_unsigned(2881, 12), 658 => to_unsigned(1302, 12), 659 => to_unsigned(2837, 12), 660 => to_unsigned(441, 12), 661 => to_unsigned(2628, 12), 662 => to_unsigned(3885, 12), 663 => to_unsigned(1000, 12), 664 => to_unsigned(4007, 12), 665 => to_unsigned(792, 12), 666 => to_unsigned(2390, 12), 667 => to_unsigned(2321, 12), 668 => to_unsigned(4020, 12), 669 => to_unsigned(3546, 12), 670 => to_unsigned(3720, 12), 671 => to_unsigned(2821, 12), 672 => to_unsigned(1249, 12), 673 => to_unsigned(342, 12), 674 => to_unsigned(250, 12), 675 => to_unsigned(3666, 12), 676 => to_unsigned(1802, 12), 677 => to_unsigned(2622, 12), 678 => to_unsigned(1565, 12), 679 => to_unsigned(139, 12), 680 => to_unsigned(2206, 12), 681 => to_unsigned(327, 12), 682 => to_unsigned(3642, 12), 683 => to_unsigned(990, 12), 684 => to_unsigned(2090, 12), 685 => to_unsigned(4053, 12), 686 => to_unsigned(2375, 12), 687 => to_unsigned(665, 12), 688 => to_unsigned(492, 12), 689 => to_unsigned(822, 12), 690 => to_unsigned(1142, 12), 691 => to_unsigned(339, 12), 692 => to_unsigned(2073, 12), 693 => to_unsigned(2221, 12), 694 => to_unsigned(1401, 12), 695 => to_unsigned(490, 12), 696 => to_unsigned(3203, 12), 697 => to_unsigned(884, 12), 698 => to_unsigned(3028, 12), 699 => to_unsigned(4081, 12), 700 => to_unsigned(851, 12), 701 => to_unsigned(2297, 12), 702 => to_unsigned(2597, 12), 703 => to_unsigned(2209, 12), 704 => to_unsigned(2492, 12), 705 => to_unsigned(876, 12), 706 => to_unsigned(3801, 12), 707 => to_unsigned(1543, 12), 708 => to_unsigned(3004, 12), 709 => to_unsigned(2213, 12), 710 => to_unsigned(3668, 12), 711 => to_unsigned(3066, 12), 712 => to_unsigned(354, 12), 713 => to_unsigned(2320, 12), 714 => to_unsigned(1709, 12), 715 => to_unsigned(1512, 12), 716 => to_unsigned(3239, 12), 717 => to_unsigned(3617, 12), 718 => to_unsigned(3937, 12), 719 => to_unsigned(1857, 12), 720 => to_unsigned(2249, 12), 721 => to_unsigned(2135, 12), 722 => to_unsigned(1348, 12), 723 => to_unsigned(2328, 12), 724 => to_unsigned(1030, 12), 725 => to_unsigned(3937, 12), 726 => to_unsigned(1394, 12), 727 => to_unsigned(767, 12), 728 => to_unsigned(3644, 12), 729 => to_unsigned(3288, 12), 730 => to_unsigned(2109, 12), 731 => to_unsigned(3060, 12), 732 => to_unsigned(3259, 12), 733 => to_unsigned(3575, 12), 734 => to_unsigned(3705, 12), 735 => to_unsigned(2506, 12), 736 => to_unsigned(797, 12), 737 => to_unsigned(1263, 12), 738 => to_unsigned(1016, 12), 739 => to_unsigned(28, 12), 740 => to_unsigned(3224, 12), 741 => to_unsigned(3459, 12), 742 => to_unsigned(466, 12), 743 => to_unsigned(1685, 12), 744 => to_unsigned(3334, 12), 745 => to_unsigned(2132, 12), 746 => to_unsigned(1301, 12), 747 => to_unsigned(3703, 12), 748 => to_unsigned(3355, 12), 749 => to_unsigned(2970, 12), 750 => to_unsigned(4057, 12), 751 => to_unsigned(448, 12), 752 => to_unsigned(2414, 12), 753 => to_unsigned(2435, 12), 754 => to_unsigned(1845, 12), 755 => to_unsigned(2853, 12), 756 => to_unsigned(2055, 12), 757 => to_unsigned(1400, 12), 758 => to_unsigned(3408, 12), 759 => to_unsigned(3531, 12), 760 => to_unsigned(2699, 12), 761 => to_unsigned(2028, 12), 762 => to_unsigned(2434, 12), 763 => to_unsigned(3382, 12), 764 => to_unsigned(1541, 12), 765 => to_unsigned(2833, 12), 766 => to_unsigned(3834, 12), 767 => to_unsigned(3965, 12), 768 => to_unsigned(3662, 12), 769 => to_unsigned(1925, 12), 770 => to_unsigned(2894, 12), 771 => to_unsigned(1105, 12), 772 => to_unsigned(1257, 12), 773 => to_unsigned(110, 12), 774 => to_unsigned(2668, 12), 775 => to_unsigned(1054, 12), 776 => to_unsigned(3938, 12), 777 => to_unsigned(1795, 12), 778 => to_unsigned(128, 12), 779 => to_unsigned(1885, 12), 780 => to_unsigned(2348, 12), 781 => to_unsigned(2732, 12), 782 => to_unsigned(1260, 12), 783 => to_unsigned(3967, 12), 784 => to_unsigned(2675, 12), 785 => to_unsigned(3005, 12), 786 => to_unsigned(2302, 12), 787 => to_unsigned(3072, 12), 788 => to_unsigned(3857, 12), 789 => to_unsigned(2461, 12), 790 => to_unsigned(1627, 12), 791 => to_unsigned(930, 12), 792 => to_unsigned(1010, 12), 793 => to_unsigned(3059, 12), 794 => to_unsigned(1252, 12), 795 => to_unsigned(1211, 12), 796 => to_unsigned(1045, 12), 797 => to_unsigned(63, 12), 798 => to_unsigned(1758, 12), 799 => to_unsigned(3576, 12), 800 => to_unsigned(1637, 12), 801 => to_unsigned(2705, 12), 802 => to_unsigned(3110, 12), 803 => to_unsigned(1743, 12), 804 => to_unsigned(2945, 12), 805 => to_unsigned(2191, 12), 806 => to_unsigned(3049, 12), 807 => to_unsigned(2774, 12), 808 => to_unsigned(1773, 12), 809 => to_unsigned(3601, 12), 810 => to_unsigned(1260, 12), 811 => to_unsigned(1973, 12), 812 => to_unsigned(3478, 12), 813 => to_unsigned(1485, 12), 814 => to_unsigned(2674, 12), 815 => to_unsigned(3247, 12), 816 => to_unsigned(1730, 12), 817 => to_unsigned(267, 12), 818 => to_unsigned(1929, 12), 819 => to_unsigned(2546, 12), 820 => to_unsigned(2856, 12), 821 => to_unsigned(4022, 12), 822 => to_unsigned(947, 12), 823 => to_unsigned(47, 12), 824 => to_unsigned(772, 12), 825 => to_unsigned(1930, 12), 826 => to_unsigned(3569, 12), 827 => to_unsigned(2302, 12), 828 => to_unsigned(646, 12), 829 => to_unsigned(3446, 12), 830 => to_unsigned(3500, 12), 831 => to_unsigned(3400, 12), 832 => to_unsigned(3464, 12), 833 => to_unsigned(2248, 12), 834 => to_unsigned(492, 12), 835 => to_unsigned(3813, 12), 836 => to_unsigned(18, 12), 837 => to_unsigned(1026, 12), 838 => to_unsigned(2245, 12), 839 => to_unsigned(3293, 12), 840 => to_unsigned(505, 12), 841 => to_unsigned(1253, 12), 842 => to_unsigned(1636, 12), 843 => to_unsigned(362, 12), 844 => to_unsigned(2205, 12), 845 => to_unsigned(1179, 12), 846 => to_unsigned(2705, 12), 847 => to_unsigned(442, 12), 848 => to_unsigned(395, 12), 849 => to_unsigned(3377, 12), 850 => to_unsigned(1352, 12), 851 => to_unsigned(344, 12), 852 => to_unsigned(1539, 12), 853 => to_unsigned(1648, 12), 854 => to_unsigned(2059, 12), 855 => to_unsigned(3897, 12), 856 => to_unsigned(3506, 12), 857 => to_unsigned(3727, 12), 858 => to_unsigned(4025, 12), 859 => to_unsigned(131, 12), 860 => to_unsigned(3958, 12), 861 => to_unsigned(3044, 12), 862 => to_unsigned(1980, 12), 863 => to_unsigned(1959, 12), 864 => to_unsigned(1534, 12), 865 => to_unsigned(2005, 12), 866 => to_unsigned(157, 12), 867 => to_unsigned(2997, 12), 868 => to_unsigned(67, 12), 869 => to_unsigned(1592, 12), 870 => to_unsigned(2251, 12), 871 => to_unsigned(3447, 12), 872 => to_unsigned(1103, 12), 873 => to_unsigned(2349, 12), 874 => to_unsigned(602, 12), 875 => to_unsigned(2127, 12), 876 => to_unsigned(3297, 12), 877 => to_unsigned(1035, 12), 878 => to_unsigned(3575, 12), 879 => to_unsigned(2181, 12), 880 => to_unsigned(926, 12), 881 => to_unsigned(3258, 12), 882 => to_unsigned(1604, 12), 883 => to_unsigned(315, 12), 884 => to_unsigned(544, 12), 885 => to_unsigned(3877, 12), 886 => to_unsigned(3243, 12), 887 => to_unsigned(637, 12), 888 => to_unsigned(3388, 12), 889 => to_unsigned(557, 12), 890 => to_unsigned(2333, 12), 891 => to_unsigned(250, 12), 892 => to_unsigned(1179, 12), 893 => to_unsigned(3815, 12), 894 => to_unsigned(795, 12), 895 => to_unsigned(1053, 12), 896 => to_unsigned(126, 12), 897 => to_unsigned(2120, 12), 898 => to_unsigned(1099, 12), 899 => to_unsigned(2145, 12), 900 => to_unsigned(3278, 12), 901 => to_unsigned(3622, 12), 902 => to_unsigned(3339, 12), 903 => to_unsigned(3530, 12), 904 => to_unsigned(1782, 12), 905 => to_unsigned(3929, 12), 906 => to_unsigned(2080, 12), 907 => to_unsigned(1714, 12), 908 => to_unsigned(3112, 12), 909 => to_unsigned(1222, 12), 910 => to_unsigned(2334, 12), 911 => to_unsigned(1686, 12), 912 => to_unsigned(1147, 12), 913 => to_unsigned(3659, 12), 914 => to_unsigned(1315, 12), 915 => to_unsigned(468, 12), 916 => to_unsigned(3012, 12), 917 => to_unsigned(1599, 12), 918 => to_unsigned(772, 12), 919 => to_unsigned(689, 12), 920 => to_unsigned(884, 12), 921 => to_unsigned(1181, 12), 922 => to_unsigned(1727, 12), 923 => to_unsigned(2877, 12), 924 => to_unsigned(603, 12), 925 => to_unsigned(3695, 12), 926 => to_unsigned(3283, 12), 927 => to_unsigned(360, 12), 928 => to_unsigned(2138, 12), 929 => to_unsigned(3610, 12), 930 => to_unsigned(585, 12), 931 => to_unsigned(1970, 12), 932 => to_unsigned(2271, 12), 933 => to_unsigned(3934, 12), 934 => to_unsigned(1809, 12), 935 => to_unsigned(1735, 12), 936 => to_unsigned(3896, 12), 937 => to_unsigned(3059, 12), 938 => to_unsigned(2851, 12), 939 => to_unsigned(201, 12), 940 => to_unsigned(1756, 12), 941 => to_unsigned(3887, 12), 942 => to_unsigned(2096, 12), 943 => to_unsigned(375, 12), 944 => to_unsigned(3015, 12), 945 => to_unsigned(2677, 12), 946 => to_unsigned(2627, 12), 947 => to_unsigned(3707, 12), 948 => to_unsigned(3783, 12), 949 => to_unsigned(2366, 12), 950 => to_unsigned(3016, 12), 951 => to_unsigned(2341, 12), 952 => to_unsigned(3077, 12), 953 => to_unsigned(3681, 12), 954 => to_unsigned(55, 12), 955 => to_unsigned(3548, 12), 956 => to_unsigned(1454, 12), 957 => to_unsigned(2086, 12), 958 => to_unsigned(561, 12), 959 => to_unsigned(2312, 12), 960 => to_unsigned(3706, 12), 961 => to_unsigned(1217, 12), 962 => to_unsigned(1346, 12), 963 => to_unsigned(1086, 12), 964 => to_unsigned(2064, 12), 965 => to_unsigned(1213, 12), 966 => to_unsigned(194, 12), 967 => to_unsigned(3339, 12), 968 => to_unsigned(2463, 12), 969 => to_unsigned(3466, 12), 970 => to_unsigned(20, 12), 971 => to_unsigned(1124, 12), 972 => to_unsigned(1806, 12), 973 => to_unsigned(3704, 12), 974 => to_unsigned(52, 12), 975 => to_unsigned(455, 12), 976 => to_unsigned(3741, 12), 977 => to_unsigned(1925, 12), 978 => to_unsigned(3342, 12), 979 => to_unsigned(1650, 12), 980 => to_unsigned(750, 12), 981 => to_unsigned(3023, 12), 982 => to_unsigned(819, 12), 983 => to_unsigned(3104, 12), 984 => to_unsigned(407, 12), 985 => to_unsigned(1785, 12), 986 => to_unsigned(859, 12), 987 => to_unsigned(774, 12), 988 => to_unsigned(1737, 12), 989 => to_unsigned(2168, 12), 990 => to_unsigned(1089, 12), 991 => to_unsigned(1099, 12), 992 => to_unsigned(855, 12), 993 => to_unsigned(2556, 12), 994 => to_unsigned(1734, 12), 995 => to_unsigned(2856, 12), 996 => to_unsigned(3772, 12), 997 => to_unsigned(1060, 12), 998 => to_unsigned(908, 12), 999 => to_unsigned(931, 12), 1000 => to_unsigned(62, 12), 1001 => to_unsigned(1477, 12), 1002 => to_unsigned(1854, 12), 1003 => to_unsigned(442, 12), 1004 => to_unsigned(588, 12), 1005 => to_unsigned(3602, 12), 1006 => to_unsigned(2432, 12), 1007 => to_unsigned(1025, 12), 1008 => to_unsigned(1748, 12), 1009 => to_unsigned(717, 12), 1010 => to_unsigned(1626, 12), 1011 => to_unsigned(1136, 12), 1012 => to_unsigned(3179, 12), 1013 => to_unsigned(1173, 12), 1014 => to_unsigned(1614, 12), 1015 => to_unsigned(1293, 12), 1016 => to_unsigned(1000, 12), 1017 => to_unsigned(3139, 12), 1018 => to_unsigned(1897, 12), 1019 => to_unsigned(2449, 12), 1020 => to_unsigned(2309, 12), 1021 => to_unsigned(26, 12), 1022 => to_unsigned(2751, 12), 1023 => to_unsigned(1435, 12), 1024 => to_unsigned(4075, 12), 1025 => to_unsigned(1773, 12), 1026 => to_unsigned(4009, 12), 1027 => to_unsigned(525, 12), 1028 => to_unsigned(2861, 12), 1029 => to_unsigned(3504, 12), 1030 => to_unsigned(568, 12), 1031 => to_unsigned(58, 12), 1032 => to_unsigned(3089, 12), 1033 => to_unsigned(1238, 12), 1034 => to_unsigned(2911, 12), 1035 => to_unsigned(3033, 12), 1036 => to_unsigned(2268, 12), 1037 => to_unsigned(3277, 12), 1038 => to_unsigned(391, 12), 1039 => to_unsigned(2330, 12), 1040 => to_unsigned(2321, 12), 1041 => to_unsigned(2756, 12), 1042 => to_unsigned(1579, 12), 1043 => to_unsigned(2479, 12), 1044 => to_unsigned(3806, 12), 1045 => to_unsigned(2173, 12), 1046 => to_unsigned(1372, 12), 1047 => to_unsigned(3577, 12), 1048 => to_unsigned(3912, 12), 1049 => to_unsigned(3770, 12), 1050 => to_unsigned(3867, 12), 1051 => to_unsigned(2054, 12), 1052 => to_unsigned(903, 12), 1053 => to_unsigned(2741, 12), 1054 => to_unsigned(3959, 12), 1055 => to_unsigned(1528, 12), 1056 => to_unsigned(2074, 12), 1057 => to_unsigned(3707, 12), 1058 => to_unsigned(715, 12), 1059 => to_unsigned(3877, 12), 1060 => to_unsigned(1117, 12), 1061 => to_unsigned(433, 12), 1062 => to_unsigned(3604, 12), 1063 => to_unsigned(477, 12), 1064 => to_unsigned(2935, 12), 1065 => to_unsigned(2488, 12), 1066 => to_unsigned(4029, 12), 1067 => to_unsigned(439, 12), 1068 => to_unsigned(732, 12), 1069 => to_unsigned(151, 12), 1070 => to_unsigned(2745, 12), 1071 => to_unsigned(1673, 12), 1072 => to_unsigned(2688, 12), 1073 => to_unsigned(3686, 12), 1074 => to_unsigned(403, 12), 1075 => to_unsigned(2503, 12), 1076 => to_unsigned(3122, 12), 1077 => to_unsigned(2598, 12), 1078 => to_unsigned(3011, 12), 1079 => to_unsigned(1788, 12), 1080 => to_unsigned(3486, 12), 1081 => to_unsigned(3621, 12), 1082 => to_unsigned(1976, 12), 1083 => to_unsigned(1918, 12), 1084 => to_unsigned(4073, 12), 1085 => to_unsigned(645, 12), 1086 => to_unsigned(59, 12), 1087 => to_unsigned(4048, 12), 1088 => to_unsigned(1498, 12), 1089 => to_unsigned(445, 12), 1090 => to_unsigned(1823, 12), 1091 => to_unsigned(966, 12), 1092 => to_unsigned(2393, 12), 1093 => to_unsigned(3275, 12), 1094 => to_unsigned(1681, 12), 1095 => to_unsigned(3103, 12), 1096 => to_unsigned(671, 12), 1097 => to_unsigned(84, 12), 1098 => to_unsigned(90, 12), 1099 => to_unsigned(1063, 12), 1100 => to_unsigned(757, 12), 1101 => to_unsigned(2226, 12), 1102 => to_unsigned(1610, 12), 1103 => to_unsigned(2342, 12), 1104 => to_unsigned(2628, 12), 1105 => to_unsigned(2427, 12), 1106 => to_unsigned(551, 12), 1107 => to_unsigned(127, 12), 1108 => to_unsigned(3279, 12), 1109 => to_unsigned(13, 12), 1110 => to_unsigned(1187, 12), 1111 => to_unsigned(486, 12), 1112 => to_unsigned(1915, 12), 1113 => to_unsigned(3467, 12), 1114 => to_unsigned(359, 12), 1115 => to_unsigned(331, 12), 1116 => to_unsigned(2032, 12), 1117 => to_unsigned(1846, 12), 1118 => to_unsigned(1444, 12), 1119 => to_unsigned(1106, 12), 1120 => to_unsigned(2251, 12), 1121 => to_unsigned(2739, 12), 1122 => to_unsigned(2210, 12), 1123 => to_unsigned(1978, 12), 1124 => to_unsigned(80, 12), 1125 => to_unsigned(540, 12), 1126 => to_unsigned(2441, 12), 1127 => to_unsigned(1893, 12), 1128 => to_unsigned(8, 12), 1129 => to_unsigned(145, 12), 1130 => to_unsigned(1776, 12), 1131 => to_unsigned(236, 12), 1132 => to_unsigned(1244, 12), 1133 => to_unsigned(1689, 12), 1134 => to_unsigned(3422, 12), 1135 => to_unsigned(3195, 12), 1136 => to_unsigned(101, 12), 1137 => to_unsigned(1723, 12), 1138 => to_unsigned(1403, 12), 1139 => to_unsigned(4062, 12), 1140 => to_unsigned(1017, 12), 1141 => to_unsigned(1083, 12), 1142 => to_unsigned(1210, 12), 1143 => to_unsigned(3346, 12), 1144 => to_unsigned(2572, 12), 1145 => to_unsigned(2945, 12), 1146 => to_unsigned(1307, 12), 1147 => to_unsigned(522, 12), 1148 => to_unsigned(1987, 12), 1149 => to_unsigned(1981, 12), 1150 => to_unsigned(784, 12), 1151 => to_unsigned(3355, 12), 1152 => to_unsigned(2684, 12), 1153 => to_unsigned(3846, 12), 1154 => to_unsigned(2560, 12), 1155 => to_unsigned(2055, 12), 1156 => to_unsigned(2713, 12), 1157 => to_unsigned(2115, 12), 1158 => to_unsigned(1851, 12), 1159 => to_unsigned(3832, 12), 1160 => to_unsigned(2420, 12), 1161 => to_unsigned(511, 12), 1162 => to_unsigned(2468, 12), 1163 => to_unsigned(2476, 12), 1164 => to_unsigned(3797, 12), 1165 => to_unsigned(2673, 12), 1166 => to_unsigned(1782, 12), 1167 => to_unsigned(2559, 12), 1168 => to_unsigned(3272, 12), 1169 => to_unsigned(2671, 12), 1170 => to_unsigned(3238, 12), 1171 => to_unsigned(1962, 12), 1172 => to_unsigned(3041, 12), 1173 => to_unsigned(3748, 12), 1174 => to_unsigned(2116, 12), 1175 => to_unsigned(91, 12), 1176 => to_unsigned(781, 12), 1177 => to_unsigned(3725, 12), 1178 => to_unsigned(2985, 12), 1179 => to_unsigned(328, 12), 1180 => to_unsigned(2694, 12), 1181 => to_unsigned(1374, 12), 1182 => to_unsigned(1164, 12), 1183 => to_unsigned(610, 12), 1184 => to_unsigned(1923, 12), 1185 => to_unsigned(2280, 12), 1186 => to_unsigned(3600, 12), 1187 => to_unsigned(2309, 12), 1188 => to_unsigned(3624, 12), 1189 => to_unsigned(1463, 12), 1190 => to_unsigned(2973, 12), 1191 => to_unsigned(1717, 12), 1192 => to_unsigned(278, 12), 1193 => to_unsigned(357, 12), 1194 => to_unsigned(2583, 12), 1195 => to_unsigned(251, 12), 1196 => to_unsigned(3962, 12), 1197 => to_unsigned(932, 12), 1198 => to_unsigned(3819, 12), 1199 => to_unsigned(187, 12), 1200 => to_unsigned(3106, 12), 1201 => to_unsigned(3014, 12), 1202 => to_unsigned(2438, 12), 1203 => to_unsigned(344, 12), 1204 => to_unsigned(1612, 12), 1205 => to_unsigned(1041, 12), 1206 => to_unsigned(1631, 12), 1207 => to_unsigned(1584, 12), 1208 => to_unsigned(3877, 12), 1209 => to_unsigned(3072, 12), 1210 => to_unsigned(3530, 12), 1211 => to_unsigned(2673, 12), 1212 => to_unsigned(2924, 12), 1213 => to_unsigned(3076, 12), 1214 => to_unsigned(3679, 12), 1215 => to_unsigned(956, 12), 1216 => to_unsigned(1663, 12), 1217 => to_unsigned(2570, 12), 1218 => to_unsigned(797, 12), 1219 => to_unsigned(865, 12), 1220 => to_unsigned(1897, 12), 1221 => to_unsigned(1264, 12), 1222 => to_unsigned(1549, 12), 1223 => to_unsigned(275, 12), 1224 => to_unsigned(41, 12), 1225 => to_unsigned(1228, 12), 1226 => to_unsigned(3500, 12), 1227 => to_unsigned(2099, 12), 1228 => to_unsigned(1131, 12), 1229 => to_unsigned(2192, 12), 1230 => to_unsigned(3576, 12), 1231 => to_unsigned(4094, 12), 1232 => to_unsigned(2802, 12), 1233 => to_unsigned(4005, 12), 1234 => to_unsigned(1550, 12), 1235 => to_unsigned(676, 12), 1236 => to_unsigned(3186, 12), 1237 => to_unsigned(1156, 12), 1238 => to_unsigned(4082, 12), 1239 => to_unsigned(303, 12), 1240 => to_unsigned(1920, 12), 1241 => to_unsigned(3889, 12), 1242 => to_unsigned(2981, 12), 1243 => to_unsigned(254, 12), 1244 => to_unsigned(459, 12), 1245 => to_unsigned(2860, 12), 1246 => to_unsigned(1605, 12), 1247 => to_unsigned(360, 12), 1248 => to_unsigned(494, 12), 1249 => to_unsigned(1808, 12), 1250 => to_unsigned(1296, 12), 1251 => to_unsigned(1802, 12), 1252 => to_unsigned(3589, 12), 1253 => to_unsigned(2967, 12), 1254 => to_unsigned(2991, 12), 1255 => to_unsigned(1603, 12), 1256 => to_unsigned(3238, 12), 1257 => to_unsigned(3056, 12), 1258 => to_unsigned(2322, 12), 1259 => to_unsigned(2142, 12), 1260 => to_unsigned(3536, 12), 1261 => to_unsigned(1823, 12), 1262 => to_unsigned(2474, 12), 1263 => to_unsigned(2095, 12), 1264 => to_unsigned(3349, 12), 1265 => to_unsigned(993, 12), 1266 => to_unsigned(3127, 12), 1267 => to_unsigned(1354, 12), 1268 => to_unsigned(2156, 12), 1269 => to_unsigned(1055, 12), 1270 => to_unsigned(595, 12), 1271 => to_unsigned(3138, 12), 1272 => to_unsigned(147, 12), 1273 => to_unsigned(3231, 12), 1274 => to_unsigned(3954, 12), 1275 => to_unsigned(2835, 12), 1276 => to_unsigned(2855, 12), 1277 => to_unsigned(1959, 12), 1278 => to_unsigned(2621, 12), 1279 => to_unsigned(609, 12), 1280 => to_unsigned(4012, 12), 1281 => to_unsigned(2292, 12), 1282 => to_unsigned(3820, 12), 1283 => to_unsigned(438, 12), 1284 => to_unsigned(3806, 12), 1285 => to_unsigned(1146, 12), 1286 => to_unsigned(2535, 12), 1287 => to_unsigned(2238, 12), 1288 => to_unsigned(2252, 12), 1289 => to_unsigned(912, 12), 1290 => to_unsigned(80, 12), 1291 => to_unsigned(2558, 12), 1292 => to_unsigned(1158, 12), 1293 => to_unsigned(1476, 12), 1294 => to_unsigned(813, 12), 1295 => to_unsigned(3028, 12), 1296 => to_unsigned(2554, 12), 1297 => to_unsigned(1694, 12), 1298 => to_unsigned(588, 12), 1299 => to_unsigned(1915, 12), 1300 => to_unsigned(693, 12), 1301 => to_unsigned(3489, 12), 1302 => to_unsigned(602, 12), 1303 => to_unsigned(1426, 12), 1304 => to_unsigned(3206, 12), 1305 => to_unsigned(632, 12), 1306 => to_unsigned(1154, 12), 1307 => to_unsigned(3226, 12), 1308 => to_unsigned(2286, 12), 1309 => to_unsigned(281, 12), 1310 => to_unsigned(2573, 12), 1311 => to_unsigned(1983, 12), 1312 => to_unsigned(2779, 12), 1313 => to_unsigned(2622, 12), 1314 => to_unsigned(3129, 12), 1315 => to_unsigned(2341, 12), 1316 => to_unsigned(941, 12), 1317 => to_unsigned(3477, 12), 1318 => to_unsigned(107, 12), 1319 => to_unsigned(504, 12), 1320 => to_unsigned(837, 12), 1321 => to_unsigned(1017, 12), 1322 => to_unsigned(1841, 12), 1323 => to_unsigned(1049, 12), 1324 => to_unsigned(268, 12), 1325 => to_unsigned(3636, 12), 1326 => to_unsigned(2886, 12), 1327 => to_unsigned(2991, 12), 1328 => to_unsigned(765, 12), 1329 => to_unsigned(73, 12), 1330 => to_unsigned(2954, 12), 1331 => to_unsigned(2632, 12), 1332 => to_unsigned(474, 12), 1333 => to_unsigned(1168, 12), 1334 => to_unsigned(1375, 12), 1335 => to_unsigned(3934, 12), 1336 => to_unsigned(766, 12), 1337 => to_unsigned(3301, 12), 1338 => to_unsigned(2342, 12), 1339 => to_unsigned(1200, 12), 1340 => to_unsigned(1724, 12), 1341 => to_unsigned(518, 12), 1342 => to_unsigned(3056, 12), 1343 => to_unsigned(966, 12), 1344 => to_unsigned(631, 12), 1345 => to_unsigned(513, 12), 1346 => to_unsigned(2415, 12), 1347 => to_unsigned(1215, 12), 1348 => to_unsigned(3265, 12), 1349 => to_unsigned(1661, 12), 1350 => to_unsigned(1301, 12), 1351 => to_unsigned(814, 12), 1352 => to_unsigned(1792, 12), 1353 => to_unsigned(3798, 12), 1354 => to_unsigned(3236, 12), 1355 => to_unsigned(3738, 12), 1356 => to_unsigned(1684, 12), 1357 => to_unsigned(340, 12), 1358 => to_unsigned(3303, 12), 1359 => to_unsigned(1570, 12), 1360 => to_unsigned(2289, 12), 1361 => to_unsigned(2926, 12), 1362 => to_unsigned(3133, 12), 1363 => to_unsigned(1950, 12), 1364 => to_unsigned(2715, 12), 1365 => to_unsigned(2788, 12), 1366 => to_unsigned(1609, 12), 1367 => to_unsigned(3400, 12), 1368 => to_unsigned(1588, 12), 1369 => to_unsigned(3668, 12), 1370 => to_unsigned(919, 12), 1371 => to_unsigned(318, 12), 1372 => to_unsigned(48, 12), 1373 => to_unsigned(2023, 12), 1374 => to_unsigned(1467, 12), 1375 => to_unsigned(1323, 12), 1376 => to_unsigned(4010, 12), 1377 => to_unsigned(653, 12), 1378 => to_unsigned(504, 12), 1379 => to_unsigned(367, 12), 1380 => to_unsigned(1017, 12), 1381 => to_unsigned(777, 12), 1382 => to_unsigned(3227, 12), 1383 => to_unsigned(3674, 12), 1384 => to_unsigned(997, 12), 1385 => to_unsigned(1570, 12), 1386 => to_unsigned(1862, 12), 1387 => to_unsigned(1449, 12), 1388 => to_unsigned(4077, 12), 1389 => to_unsigned(1061, 12), 1390 => to_unsigned(6, 12), 1391 => to_unsigned(3386, 12), 1392 => to_unsigned(597, 12), 1393 => to_unsigned(1027, 12), 1394 => to_unsigned(2123, 12), 1395 => to_unsigned(3818, 12), 1396 => to_unsigned(3339, 12), 1397 => to_unsigned(2461, 12), 1398 => to_unsigned(2126, 12), 1399 => to_unsigned(723, 12), 1400 => to_unsigned(1306, 12), 1401 => to_unsigned(2411, 12), 1402 => to_unsigned(2815, 12), 1403 => to_unsigned(80, 12), 1404 => to_unsigned(1187, 12), 1405 => to_unsigned(1588, 12), 1406 => to_unsigned(913, 12), 1407 => to_unsigned(3664, 12), 1408 => to_unsigned(2442, 12), 1409 => to_unsigned(4089, 12), 1410 => to_unsigned(1212, 12), 1411 => to_unsigned(969, 12), 1412 => to_unsigned(99, 12), 1413 => to_unsigned(921, 12), 1414 => to_unsigned(1663, 12), 1415 => to_unsigned(3226, 12), 1416 => to_unsigned(563, 12), 1417 => to_unsigned(335, 12), 1418 => to_unsigned(2331, 12), 1419 => to_unsigned(2180, 12), 1420 => to_unsigned(3430, 12), 1421 => to_unsigned(3797, 12), 1422 => to_unsigned(2151, 12), 1423 => to_unsigned(2289, 12), 1424 => to_unsigned(2485, 12), 1425 => to_unsigned(3863, 12), 1426 => to_unsigned(1004, 12), 1427 => to_unsigned(4070, 12), 1428 => to_unsigned(3435, 12), 1429 => to_unsigned(2667, 12), 1430 => to_unsigned(1558, 12), 1431 => to_unsigned(1372, 12), 1432 => to_unsigned(4078, 12), 1433 => to_unsigned(3115, 12), 1434 => to_unsigned(1030, 12), 1435 => to_unsigned(909, 12), 1436 => to_unsigned(1229, 12), 1437 => to_unsigned(145, 12), 1438 => to_unsigned(3496, 12), 1439 => to_unsigned(2685, 12), 1440 => to_unsigned(478, 12), 1441 => to_unsigned(1476, 12), 1442 => to_unsigned(1810, 12), 1443 => to_unsigned(752, 12), 1444 => to_unsigned(1154, 12), 1445 => to_unsigned(27, 12), 1446 => to_unsigned(392, 12), 1447 => to_unsigned(3819, 12), 1448 => to_unsigned(1231, 12), 1449 => to_unsigned(1587, 12), 1450 => to_unsigned(215, 12), 1451 => to_unsigned(1967, 12), 1452 => to_unsigned(2879, 12), 1453 => to_unsigned(3230, 12), 1454 => to_unsigned(2573, 12), 1455 => to_unsigned(2908, 12), 1456 => to_unsigned(2990, 12), 1457 => to_unsigned(3982, 12), 1458 => to_unsigned(3826, 12), 1459 => to_unsigned(3246, 12), 1460 => to_unsigned(3245, 12), 1461 => to_unsigned(1633, 12), 1462 => to_unsigned(260, 12), 1463 => to_unsigned(884, 12), 1464 => to_unsigned(650, 12), 1465 => to_unsigned(1396, 12), 1466 => to_unsigned(63, 12), 1467 => to_unsigned(274, 12), 1468 => to_unsigned(3556, 12), 1469 => to_unsigned(2248, 12), 1470 => to_unsigned(119, 12), 1471 => to_unsigned(2362, 12), 1472 => to_unsigned(3785, 12), 1473 => to_unsigned(2798, 12), 1474 => to_unsigned(3469, 12), 1475 => to_unsigned(3596, 12), 1476 => to_unsigned(669, 12), 1477 => to_unsigned(2638, 12), 1478 => to_unsigned(2408, 12), 1479 => to_unsigned(77, 12), 1480 => to_unsigned(3721, 12), 1481 => to_unsigned(4014, 12), 1482 => to_unsigned(700, 12), 1483 => to_unsigned(588, 12), 1484 => to_unsigned(1253, 12), 1485 => to_unsigned(3741, 12), 1486 => to_unsigned(3181, 12), 1487 => to_unsigned(75, 12), 1488 => to_unsigned(3564, 12), 1489 => to_unsigned(2025, 12), 1490 => to_unsigned(1905, 12), 1491 => to_unsigned(1944, 12), 1492 => to_unsigned(3899, 12), 1493 => to_unsigned(4040, 12), 1494 => to_unsigned(2703, 12), 1495 => to_unsigned(2486, 12), 1496 => to_unsigned(672, 12), 1497 => to_unsigned(492, 12), 1498 => to_unsigned(1278, 12), 1499 => to_unsigned(3792, 12), 1500 => to_unsigned(1010, 12), 1501 => to_unsigned(2419, 12), 1502 => to_unsigned(3692, 12), 1503 => to_unsigned(1138, 12), 1504 => to_unsigned(3441, 12), 1505 => to_unsigned(11, 12), 1506 => to_unsigned(2319, 12), 1507 => to_unsigned(1305, 12), 1508 => to_unsigned(789, 12), 1509 => to_unsigned(2198, 12), 1510 => to_unsigned(2001, 12), 1511 => to_unsigned(3036, 12), 1512 => to_unsigned(762, 12), 1513 => to_unsigned(1883, 12), 1514 => to_unsigned(108, 12), 1515 => to_unsigned(456, 12), 1516 => to_unsigned(859, 12), 1517 => to_unsigned(476, 12), 1518 => to_unsigned(2791, 12), 1519 => to_unsigned(2667, 12), 1520 => to_unsigned(103, 12), 1521 => to_unsigned(99, 12), 1522 => to_unsigned(2462, 12), 1523 => to_unsigned(1780, 12), 1524 => to_unsigned(4009, 12), 1525 => to_unsigned(1782, 12), 1526 => to_unsigned(393, 12), 1527 => to_unsigned(886, 12), 1528 => to_unsigned(820, 12), 1529 => to_unsigned(3371, 12), 1530 => to_unsigned(2897, 12), 1531 => to_unsigned(1970, 12), 1532 => to_unsigned(1424, 12), 1533 => to_unsigned(3136, 12), 1534 => to_unsigned(1818, 12), 1535 => to_unsigned(2183, 12), 1536 => to_unsigned(1462, 12), 1537 => to_unsigned(2898, 12), 1538 => to_unsigned(4026, 12), 1539 => to_unsigned(1355, 12), 1540 => to_unsigned(2361, 12), 1541 => to_unsigned(3770, 12), 1542 => to_unsigned(3020, 12), 1543 => to_unsigned(2317, 12), 1544 => to_unsigned(968, 12), 1545 => to_unsigned(232, 12), 1546 => to_unsigned(3858, 12), 1547 => to_unsigned(3217, 12), 1548 => to_unsigned(1194, 12), 1549 => to_unsigned(3372, 12), 1550 => to_unsigned(3298, 12), 1551 => to_unsigned(1739, 12), 1552 => to_unsigned(2903, 12), 1553 => to_unsigned(838, 12), 1554 => to_unsigned(2254, 12), 1555 => to_unsigned(3630, 12), 1556 => to_unsigned(3638, 12), 1557 => to_unsigned(3762, 12), 1558 => to_unsigned(43, 12), 1559 => to_unsigned(577, 12), 1560 => to_unsigned(3022, 12), 1561 => to_unsigned(357, 12), 1562 => to_unsigned(2310, 12), 1563 => to_unsigned(2169, 12), 1564 => to_unsigned(1199, 12), 1565 => to_unsigned(3244, 12), 1566 => to_unsigned(2825, 12), 1567 => to_unsigned(515, 12), 1568 => to_unsigned(1417, 12), 1569 => to_unsigned(123, 12), 1570 => to_unsigned(3828, 12), 1571 => to_unsigned(2555, 12), 1572 => to_unsigned(1058, 12), 1573 => to_unsigned(3550, 12), 1574 => to_unsigned(2561, 12), 1575 => to_unsigned(1318, 12), 1576 => to_unsigned(2254, 12), 1577 => to_unsigned(2000, 12), 1578 => to_unsigned(2910, 12), 1579 => to_unsigned(3506, 12), 1580 => to_unsigned(141, 12), 1581 => to_unsigned(1878, 12), 1582 => to_unsigned(2094, 12), 1583 => to_unsigned(3043, 12), 1584 => to_unsigned(855, 12), 1585 => to_unsigned(805, 12), 1586 => to_unsigned(3933, 12), 1587 => to_unsigned(3821, 12), 1588 => to_unsigned(2794, 12), 1589 => to_unsigned(3418, 12), 1590 => to_unsigned(82, 12), 1591 => to_unsigned(4054, 12), 1592 => to_unsigned(518, 12), 1593 => to_unsigned(1610, 12), 1594 => to_unsigned(3499, 12), 1595 => to_unsigned(2561, 12), 1596 => to_unsigned(3529, 12), 1597 => to_unsigned(2522, 12), 1598 => to_unsigned(176, 12), 1599 => to_unsigned(2895, 12), 1600 => to_unsigned(1425, 12), 1601 => to_unsigned(3347, 12), 1602 => to_unsigned(254, 12), 1603 => to_unsigned(1171, 12), 1604 => to_unsigned(2881, 12), 1605 => to_unsigned(1435, 12), 1606 => to_unsigned(2035, 12), 1607 => to_unsigned(1764, 12), 1608 => to_unsigned(931, 12), 1609 => to_unsigned(2313, 12), 1610 => to_unsigned(745, 12), 1611 => to_unsigned(13, 12), 1612 => to_unsigned(437, 12), 1613 => to_unsigned(3398, 12), 1614 => to_unsigned(984, 12), 1615 => to_unsigned(778, 12), 1616 => to_unsigned(121, 12), 1617 => to_unsigned(1323, 12), 1618 => to_unsigned(3685, 12), 1619 => to_unsigned(1413, 12), 1620 => to_unsigned(168, 12), 1621 => to_unsigned(1268, 12), 1622 => to_unsigned(783, 12), 1623 => to_unsigned(1038, 12), 1624 => to_unsigned(2517, 12), 1625 => to_unsigned(0, 12), 1626 => to_unsigned(1315, 12), 1627 => to_unsigned(1633, 12), 1628 => to_unsigned(3470, 12), 1629 => to_unsigned(1798, 12), 1630 => to_unsigned(600, 12), 1631 => to_unsigned(3574, 12), 1632 => to_unsigned(1027, 12), 1633 => to_unsigned(1348, 12), 1634 => to_unsigned(1125, 12), 1635 => to_unsigned(3560, 12), 1636 => to_unsigned(2911, 12), 1637 => to_unsigned(1947, 12), 1638 => to_unsigned(626, 12), 1639 => to_unsigned(2025, 12), 1640 => to_unsigned(2627, 12), 1641 => to_unsigned(3874, 12), 1642 => to_unsigned(425, 12), 1643 => to_unsigned(781, 12), 1644 => to_unsigned(3967, 12), 1645 => to_unsigned(1137, 12), 1646 => to_unsigned(2449, 12), 1647 => to_unsigned(362, 12), 1648 => to_unsigned(2728, 12), 1649 => to_unsigned(3565, 12), 1650 => to_unsigned(970, 12), 1651 => to_unsigned(2854, 12), 1652 => to_unsigned(3626, 12), 1653 => to_unsigned(323, 12), 1654 => to_unsigned(1307, 12), 1655 => to_unsigned(4028, 12), 1656 => to_unsigned(655, 12), 1657 => to_unsigned(2802, 12), 1658 => to_unsigned(1954, 12), 1659 => to_unsigned(3556, 12), 1660 => to_unsigned(746, 12), 1661 => to_unsigned(3687, 12), 1662 => to_unsigned(3762, 12), 1663 => to_unsigned(2092, 12), 1664 => to_unsigned(340, 12), 1665 => to_unsigned(564, 12), 1666 => to_unsigned(1945, 12), 1667 => to_unsigned(3787, 12), 1668 => to_unsigned(172, 12), 1669 => to_unsigned(81, 12), 1670 => to_unsigned(4095, 12), 1671 => to_unsigned(645, 12), 1672 => to_unsigned(1619, 12), 1673 => to_unsigned(711, 12), 1674 => to_unsigned(255, 12), 1675 => to_unsigned(1860, 12), 1676 => to_unsigned(3679, 12), 1677 => to_unsigned(3421, 12), 1678 => to_unsigned(106, 12), 1679 => to_unsigned(754, 12), 1680 => to_unsigned(1627, 12), 1681 => to_unsigned(1184, 12), 1682 => to_unsigned(3563, 12), 1683 => to_unsigned(937, 12), 1684 => to_unsigned(3282, 12), 1685 => to_unsigned(413, 12), 1686 => to_unsigned(3981, 12), 1687 => to_unsigned(4082, 12), 1688 => to_unsigned(1388, 12), 1689 => to_unsigned(2697, 12), 1690 => to_unsigned(54, 12), 1691 => to_unsigned(2952, 12), 1692 => to_unsigned(3097, 12), 1693 => to_unsigned(2209, 12), 1694 => to_unsigned(529, 12), 1695 => to_unsigned(497, 12), 1696 => to_unsigned(2479, 12), 1697 => to_unsigned(3600, 12), 1698 => to_unsigned(1585, 12), 1699 => to_unsigned(3134, 12), 1700 => to_unsigned(839, 12), 1701 => to_unsigned(3934, 12), 1702 => to_unsigned(4094, 12), 1703 => to_unsigned(3024, 12), 1704 => to_unsigned(1110, 12), 1705 => to_unsigned(2555, 12), 1706 => to_unsigned(2213, 12), 1707 => to_unsigned(1289, 12), 1708 => to_unsigned(4014, 12), 1709 => to_unsigned(652, 12), 1710 => to_unsigned(1112, 12), 1711 => to_unsigned(1405, 12), 1712 => to_unsigned(1397, 12), 1713 => to_unsigned(2454, 12), 1714 => to_unsigned(3256, 12), 1715 => to_unsigned(3662, 12), 1716 => to_unsigned(2605, 12), 1717 => to_unsigned(1825, 12), 1718 => to_unsigned(702, 12), 1719 => to_unsigned(2564, 12), 1720 => to_unsigned(2885, 12), 1721 => to_unsigned(637, 12), 1722 => to_unsigned(1100, 12), 1723 => to_unsigned(681, 12), 1724 => to_unsigned(2444, 12), 1725 => to_unsigned(3840, 12), 1726 => to_unsigned(3781, 12), 1727 => to_unsigned(2198, 12), 1728 => to_unsigned(1769, 12), 1729 => to_unsigned(3425, 12), 1730 => to_unsigned(2737, 12), 1731 => to_unsigned(3699, 12), 1732 => to_unsigned(3905, 12), 1733 => to_unsigned(2442, 12), 1734 => to_unsigned(198, 12), 1735 => to_unsigned(2170, 12), 1736 => to_unsigned(2064, 12), 1737 => to_unsigned(2759, 12), 1738 => to_unsigned(2459, 12), 1739 => to_unsigned(3366, 12), 1740 => to_unsigned(2155, 12), 1741 => to_unsigned(3156, 12), 1742 => to_unsigned(1449, 12), 1743 => to_unsigned(722, 12), 1744 => to_unsigned(627, 12), 1745 => to_unsigned(4074, 12), 1746 => to_unsigned(454, 12), 1747 => to_unsigned(2982, 12), 1748 => to_unsigned(3746, 12), 1749 => to_unsigned(2161, 12), 1750 => to_unsigned(714, 12), 1751 => to_unsigned(3839, 12), 1752 => to_unsigned(359, 12), 1753 => to_unsigned(1832, 12), 1754 => to_unsigned(40, 12), 1755 => to_unsigned(3995, 12), 1756 => to_unsigned(94, 12), 1757 => to_unsigned(4091, 12), 1758 => to_unsigned(3236, 12), 1759 => to_unsigned(2146, 12), 1760 => to_unsigned(571, 12), 1761 => to_unsigned(2649, 12), 1762 => to_unsigned(1947, 12), 1763 => to_unsigned(696, 12), 1764 => to_unsigned(3199, 12), 1765 => to_unsigned(954, 12), 1766 => to_unsigned(1311, 12), 1767 => to_unsigned(2864, 12), 1768 => to_unsigned(3051, 12), 1769 => to_unsigned(2174, 12), 1770 => to_unsigned(387, 12), 1771 => to_unsigned(320, 12), 1772 => to_unsigned(3621, 12), 1773 => to_unsigned(503, 12), 1774 => to_unsigned(1703, 12), 1775 => to_unsigned(1036, 12), 1776 => to_unsigned(2900, 12), 1777 => to_unsigned(3531, 12), 1778 => to_unsigned(2380, 12), 1779 => to_unsigned(1656, 12), 1780 => to_unsigned(370, 12), 1781 => to_unsigned(4059, 12), 1782 => to_unsigned(943, 12), 1783 => to_unsigned(313, 12), 1784 => to_unsigned(2197, 12), 1785 => to_unsigned(3948, 12), 1786 => to_unsigned(524, 12), 1787 => to_unsigned(2031, 12), 1788 => to_unsigned(657, 12), 1789 => to_unsigned(2471, 12), 1790 => to_unsigned(3999, 12), 1791 => to_unsigned(1647, 12), 1792 => to_unsigned(1693, 12), 1793 => to_unsigned(2487, 12), 1794 => to_unsigned(2497, 12), 1795 => to_unsigned(1317, 12), 1796 => to_unsigned(2560, 12), 1797 => to_unsigned(791, 12), 1798 => to_unsigned(909, 12), 1799 => to_unsigned(136, 12), 1800 => to_unsigned(2516, 12), 1801 => to_unsigned(2101, 12), 1802 => to_unsigned(2258, 12), 1803 => to_unsigned(2384, 12), 1804 => to_unsigned(3853, 12), 1805 => to_unsigned(2440, 12), 1806 => to_unsigned(3462, 12), 1807 => to_unsigned(411, 12), 1808 => to_unsigned(3237, 12), 1809 => to_unsigned(419, 12), 1810 => to_unsigned(3624, 12), 1811 => to_unsigned(3738, 12), 1812 => to_unsigned(2398, 12), 1813 => to_unsigned(972, 12), 1814 => to_unsigned(3513, 12), 1815 => to_unsigned(2349, 12), 1816 => to_unsigned(3920, 12), 1817 => to_unsigned(3386, 12), 1818 => to_unsigned(3223, 12), 1819 => to_unsigned(2814, 12), 1820 => to_unsigned(3314, 12), 1821 => to_unsigned(746, 12), 1822 => to_unsigned(968, 12), 1823 => to_unsigned(4087, 12), 1824 => to_unsigned(3062, 12), 1825 => to_unsigned(2512, 12), 1826 => to_unsigned(3317, 12), 1827 => to_unsigned(2941, 12), 1828 => to_unsigned(1554, 12), 1829 => to_unsigned(970, 12), 1830 => to_unsigned(1935, 12), 1831 => to_unsigned(486, 12), 1832 => to_unsigned(1917, 12), 1833 => to_unsigned(856, 12), 1834 => to_unsigned(2020, 12), 1835 => to_unsigned(1775, 12), 1836 => to_unsigned(2880, 12), 1837 => to_unsigned(3459, 12), 1838 => to_unsigned(4058, 12), 1839 => to_unsigned(2964, 12), 1840 => to_unsigned(1007, 12), 1841 => to_unsigned(3247, 12), 1842 => to_unsigned(2494, 12), 1843 => to_unsigned(353, 12), 1844 => to_unsigned(3096, 12), 1845 => to_unsigned(2770, 12), 1846 => to_unsigned(1832, 12), 1847 => to_unsigned(2185, 12), 1848 => to_unsigned(1352, 12), 1849 => to_unsigned(3271, 12), 1850 => to_unsigned(3548, 12), 1851 => to_unsigned(2031, 12), 1852 => to_unsigned(297, 12), 1853 => to_unsigned(1811, 12), 1854 => to_unsigned(2774, 12), 1855 => to_unsigned(1347, 12), 1856 => to_unsigned(2039, 12), 1857 => to_unsigned(1998, 12), 1858 => to_unsigned(3199, 12), 1859 => to_unsigned(3703, 12), 1860 => to_unsigned(3906, 12), 1861 => to_unsigned(1751, 12), 1862 => to_unsigned(235, 12), 1863 => to_unsigned(1048, 12), 1864 => to_unsigned(3668, 12), 1865 => to_unsigned(1699, 12), 1866 => to_unsigned(1914, 12), 1867 => to_unsigned(3502, 12), 1868 => to_unsigned(544, 12), 1869 => to_unsigned(802, 12), 1870 => to_unsigned(1578, 12), 1871 => to_unsigned(860, 12), 1872 => to_unsigned(2085, 12), 1873 => to_unsigned(228, 12), 1874 => to_unsigned(850, 12), 1875 => to_unsigned(1079, 12), 1876 => to_unsigned(1898, 12), 1877 => to_unsigned(2595, 12), 1878 => to_unsigned(4071, 12), 1879 => to_unsigned(355, 12), 1880 => to_unsigned(3137, 12), 1881 => to_unsigned(2397, 12), 1882 => to_unsigned(1684, 12), 1883 => to_unsigned(1253, 12), 1884 => to_unsigned(2403, 12), 1885 => to_unsigned(814, 12), 1886 => to_unsigned(3426, 12), 1887 => to_unsigned(91, 12), 1888 => to_unsigned(2110, 12), 1889 => to_unsigned(2110, 12), 1890 => to_unsigned(497, 12), 1891 => to_unsigned(2299, 12), 1892 => to_unsigned(2638, 12), 1893 => to_unsigned(874, 12), 1894 => to_unsigned(2206, 12), 1895 => to_unsigned(3419, 12), 1896 => to_unsigned(51, 12), 1897 => to_unsigned(2564, 12), 1898 => to_unsigned(1732, 12), 1899 => to_unsigned(902, 12), 1900 => to_unsigned(3817, 12), 1901 => to_unsigned(3881, 12), 1902 => to_unsigned(3331, 12), 1903 => to_unsigned(2727, 12), 1904 => to_unsigned(2540, 12), 1905 => to_unsigned(3172, 12), 1906 => to_unsigned(2459, 12), 1907 => to_unsigned(3725, 12), 1908 => to_unsigned(300, 12), 1909 => to_unsigned(2304, 12), 1910 => to_unsigned(1866, 12), 1911 => to_unsigned(2781, 12), 1912 => to_unsigned(846, 12), 1913 => to_unsigned(1152, 12), 1914 => to_unsigned(3328, 12), 1915 => to_unsigned(2144, 12), 1916 => to_unsigned(1908, 12), 1917 => to_unsigned(3851, 12), 1918 => to_unsigned(2077, 12), 1919 => to_unsigned(3461, 12), 1920 => to_unsigned(2117, 12), 1921 => to_unsigned(697, 12), 1922 => to_unsigned(1310, 12), 1923 => to_unsigned(2834, 12), 1924 => to_unsigned(618, 12), 1925 => to_unsigned(16, 12), 1926 => to_unsigned(1911, 12), 1927 => to_unsigned(3409, 12), 1928 => to_unsigned(1227, 12), 1929 => to_unsigned(2057, 12), 1930 => to_unsigned(1929, 12), 1931 => to_unsigned(2778, 12), 1932 => to_unsigned(1100, 12), 1933 => to_unsigned(1728, 12), 1934 => to_unsigned(1255, 12), 1935 => to_unsigned(1948, 12), 1936 => to_unsigned(1782, 12), 1937 => to_unsigned(2893, 12), 1938 => to_unsigned(855, 12), 1939 => to_unsigned(3002, 12), 1940 => to_unsigned(2681, 12), 1941 => to_unsigned(3504, 12), 1942 => to_unsigned(3483, 12), 1943 => to_unsigned(1899, 12), 1944 => to_unsigned(153, 12), 1945 => to_unsigned(2004, 12), 1946 => to_unsigned(2159, 12), 1947 => to_unsigned(1612, 12), 1948 => to_unsigned(1560, 12), 1949 => to_unsigned(3845, 12), 1950 => to_unsigned(1058, 12), 1951 => to_unsigned(76, 12), 1952 => to_unsigned(3259, 12), 1953 => to_unsigned(3627, 12), 1954 => to_unsigned(975, 12), 1955 => to_unsigned(827, 12), 1956 => to_unsigned(3349, 12), 1957 => to_unsigned(3556, 12), 1958 => to_unsigned(3569, 12), 1959 => to_unsigned(2558, 12), 1960 => to_unsigned(2412, 12), 1961 => to_unsigned(1548, 12), 1962 => to_unsigned(2928, 12), 1963 => to_unsigned(3170, 12), 1964 => to_unsigned(645, 12), 1965 => to_unsigned(3860, 12), 1966 => to_unsigned(1660, 12), 1967 => to_unsigned(2719, 12), 1968 => to_unsigned(1890, 12), 1969 => to_unsigned(2327, 12), 1970 => to_unsigned(1555, 12), 1971 => to_unsigned(2645, 12), 1972 => to_unsigned(2863, 12), 1973 => to_unsigned(2042, 12), 1974 => to_unsigned(3846, 12), 1975 => to_unsigned(68, 12), 1976 => to_unsigned(1225, 12), 1977 => to_unsigned(3608, 12), 1978 => to_unsigned(943, 12), 1979 => to_unsigned(4000, 12), 1980 => to_unsigned(1994, 12), 1981 => to_unsigned(2778, 12), 1982 => to_unsigned(475, 12), 1983 => to_unsigned(1296, 12), 1984 => to_unsigned(1762, 12), 1985 => to_unsigned(3222, 12), 1986 => to_unsigned(1149, 12), 1987 => to_unsigned(1052, 12), 1988 => to_unsigned(284, 12), 1989 => to_unsigned(2673, 12), 1990 => to_unsigned(4046, 12), 1991 => to_unsigned(2917, 12), 1992 => to_unsigned(2649, 12), 1993 => to_unsigned(1157, 12), 1994 => to_unsigned(1602, 12), 1995 => to_unsigned(1443, 12), 1996 => to_unsigned(715, 12), 1997 => to_unsigned(2995, 12), 1998 => to_unsigned(2637, 12), 1999 => to_unsigned(2019, 12), 2000 => to_unsigned(2744, 12), 2001 => to_unsigned(3551, 12), 2002 => to_unsigned(1502, 12), 2003 => to_unsigned(3333, 12), 2004 => to_unsigned(2077, 12), 2005 => to_unsigned(2139, 12), 2006 => to_unsigned(2041, 12), 2007 => to_unsigned(4021, 12), 2008 => to_unsigned(449, 12), 2009 => to_unsigned(1341, 12), 2010 => to_unsigned(488, 12), 2011 => to_unsigned(3226, 12), 2012 => to_unsigned(3356, 12), 2013 => to_unsigned(999, 12), 2014 => to_unsigned(2471, 12), 2015 => to_unsigned(3681, 12), 2016 => to_unsigned(105, 12), 2017 => to_unsigned(2735, 12), 2018 => to_unsigned(2157, 12), 2019 => to_unsigned(1952, 12), 2020 => to_unsigned(377, 12), 2021 => to_unsigned(260, 12), 2022 => to_unsigned(1462, 12), 2023 => to_unsigned(2432, 12), 2024 => to_unsigned(267, 12), 2025 => to_unsigned(179, 12), 2026 => to_unsigned(611, 12), 2027 => to_unsigned(964, 12), 2028 => to_unsigned(3866, 12), 2029 => to_unsigned(3599, 12), 2030 => to_unsigned(2545, 12), 2031 => to_unsigned(732, 12), 2032 => to_unsigned(2922, 12), 2033 => to_unsigned(912, 12), 2034 => to_unsigned(884, 12), 2035 => to_unsigned(1094, 12), 2036 => to_unsigned(2808, 12), 2037 => to_unsigned(2143, 12), 2038 => to_unsigned(1026, 12), 2039 => to_unsigned(508, 12), 2040 => to_unsigned(3345, 12), 2041 => to_unsigned(3314, 12), 2042 => to_unsigned(3905, 12), 2043 => to_unsigned(2208, 12), 2044 => to_unsigned(2273, 12), 2045 => to_unsigned(1446, 12), 2046 => to_unsigned(2628, 12), 2047 => to_unsigned(1886, 12)),
            2 => (0 => to_unsigned(3332, 12), 1 => to_unsigned(1019, 12), 2 => to_unsigned(2383, 12), 3 => to_unsigned(1151, 12), 4 => to_unsigned(277, 12), 5 => to_unsigned(3961, 12), 6 => to_unsigned(1395, 12), 7 => to_unsigned(1126, 12), 8 => to_unsigned(1802, 12), 9 => to_unsigned(272, 12), 10 => to_unsigned(2050, 12), 11 => to_unsigned(1838, 12), 12 => to_unsigned(701, 12), 13 => to_unsigned(2222, 12), 14 => to_unsigned(1134, 12), 15 => to_unsigned(2336, 12), 16 => to_unsigned(231, 12), 17 => to_unsigned(1943, 12), 18 => to_unsigned(3773, 12), 19 => to_unsigned(385, 12), 20 => to_unsigned(3364, 12), 21 => to_unsigned(3929, 12), 22 => to_unsigned(264, 12), 23 => to_unsigned(1583, 12), 24 => to_unsigned(2907, 12), 25 => to_unsigned(1024, 12), 26 => to_unsigned(163, 12), 27 => to_unsigned(3098, 12), 28 => to_unsigned(1214, 12), 29 => to_unsigned(1903, 12), 30 => to_unsigned(2996, 12), 31 => to_unsigned(4074, 12), 32 => to_unsigned(1686, 12), 33 => to_unsigned(2719, 12), 34 => to_unsigned(3713, 12), 35 => to_unsigned(1885, 12), 36 => to_unsigned(2307, 12), 37 => to_unsigned(259, 12), 38 => to_unsigned(1378, 12), 39 => to_unsigned(1140, 12), 40 => to_unsigned(164, 12), 41 => to_unsigned(2474, 12), 42 => to_unsigned(366, 12), 43 => to_unsigned(1044, 12), 44 => to_unsigned(1257, 12), 45 => to_unsigned(2181, 12), 46 => to_unsigned(2776, 12), 47 => to_unsigned(1023, 12), 48 => to_unsigned(3155, 12), 49 => to_unsigned(694, 12), 50 => to_unsigned(741, 12), 51 => to_unsigned(3331, 12), 52 => to_unsigned(3923, 12), 53 => to_unsigned(1175, 12), 54 => to_unsigned(3120, 12), 55 => to_unsigned(2910, 12), 56 => to_unsigned(670, 12), 57 => to_unsigned(1241, 12), 58 => to_unsigned(1927, 12), 59 => to_unsigned(4010, 12), 60 => to_unsigned(652, 12), 61 => to_unsigned(3588, 12), 62 => to_unsigned(240, 12), 63 => to_unsigned(923, 12), 64 => to_unsigned(204, 12), 65 => to_unsigned(3695, 12), 66 => to_unsigned(714, 12), 67 => to_unsigned(3836, 12), 68 => to_unsigned(427, 12), 69 => to_unsigned(3765, 12), 70 => to_unsigned(238, 12), 71 => to_unsigned(3722, 12), 72 => to_unsigned(2803, 12), 73 => to_unsigned(43, 12), 74 => to_unsigned(1798, 12), 75 => to_unsigned(711, 12), 76 => to_unsigned(2560, 12), 77 => to_unsigned(563, 12), 78 => to_unsigned(674, 12), 79 => to_unsigned(2912, 12), 80 => to_unsigned(3095, 12), 81 => to_unsigned(1472, 12), 82 => to_unsigned(1735, 12), 83 => to_unsigned(3998, 12), 84 => to_unsigned(786, 12), 85 => to_unsigned(800, 12), 86 => to_unsigned(2, 12), 87 => to_unsigned(3750, 12), 88 => to_unsigned(3340, 12), 89 => to_unsigned(1600, 12), 90 => to_unsigned(894, 12), 91 => to_unsigned(764, 12), 92 => to_unsigned(3144, 12), 93 => to_unsigned(1795, 12), 94 => to_unsigned(3469, 12), 95 => to_unsigned(894, 12), 96 => to_unsigned(2010, 12), 97 => to_unsigned(131, 12), 98 => to_unsigned(1254, 12), 99 => to_unsigned(2502, 12), 100 => to_unsigned(3718, 12), 101 => to_unsigned(2452, 12), 102 => to_unsigned(826, 12), 103 => to_unsigned(2050, 12), 104 => to_unsigned(981, 12), 105 => to_unsigned(175, 12), 106 => to_unsigned(1535, 12), 107 => to_unsigned(3764, 12), 108 => to_unsigned(3642, 12), 109 => to_unsigned(110, 12), 110 => to_unsigned(1618, 12), 111 => to_unsigned(254, 12), 112 => to_unsigned(1616, 12), 113 => to_unsigned(2361, 12), 114 => to_unsigned(3755, 12), 115 => to_unsigned(1313, 12), 116 => to_unsigned(3562, 12), 117 => to_unsigned(69, 12), 118 => to_unsigned(3293, 12), 119 => to_unsigned(1103, 12), 120 => to_unsigned(3161, 12), 121 => to_unsigned(493, 12), 122 => to_unsigned(3061, 12), 123 => to_unsigned(1304, 12), 124 => to_unsigned(356, 12), 125 => to_unsigned(2748, 12), 126 => to_unsigned(889, 12), 127 => to_unsigned(2880, 12), 128 => to_unsigned(1469, 12), 129 => to_unsigned(1101, 12), 130 => to_unsigned(1548, 12), 131 => to_unsigned(710, 12), 132 => to_unsigned(1137, 12), 133 => to_unsigned(2609, 12), 134 => to_unsigned(131, 12), 135 => to_unsigned(928, 12), 136 => to_unsigned(3187, 12), 137 => to_unsigned(1713, 12), 138 => to_unsigned(3811, 12), 139 => to_unsigned(2445, 12), 140 => to_unsigned(75, 12), 141 => to_unsigned(3089, 12), 142 => to_unsigned(68, 12), 143 => to_unsigned(3543, 12), 144 => to_unsigned(2351, 12), 145 => to_unsigned(330, 12), 146 => to_unsigned(2470, 12), 147 => to_unsigned(2676, 12), 148 => to_unsigned(3317, 12), 149 => to_unsigned(870, 12), 150 => to_unsigned(2480, 12), 151 => to_unsigned(1572, 12), 152 => to_unsigned(1501, 12), 153 => to_unsigned(793, 12), 154 => to_unsigned(547, 12), 155 => to_unsigned(3527, 12), 156 => to_unsigned(960, 12), 157 => to_unsigned(1856, 12), 158 => to_unsigned(1032, 12), 159 => to_unsigned(3011, 12), 160 => to_unsigned(2822, 12), 161 => to_unsigned(3173, 12), 162 => to_unsigned(3068, 12), 163 => to_unsigned(3463, 12), 164 => to_unsigned(947, 12), 165 => to_unsigned(3533, 12), 166 => to_unsigned(82, 12), 167 => to_unsigned(2424, 12), 168 => to_unsigned(1553, 12), 169 => to_unsigned(3843, 12), 170 => to_unsigned(3198, 12), 171 => to_unsigned(3336, 12), 172 => to_unsigned(47, 12), 173 => to_unsigned(1579, 12), 174 => to_unsigned(3773, 12), 175 => to_unsigned(1795, 12), 176 => to_unsigned(300, 12), 177 => to_unsigned(2123, 12), 178 => to_unsigned(4085, 12), 179 => to_unsigned(2353, 12), 180 => to_unsigned(1074, 12), 181 => to_unsigned(3210, 12), 182 => to_unsigned(1195, 12), 183 => to_unsigned(719, 12), 184 => to_unsigned(987, 12), 185 => to_unsigned(3174, 12), 186 => to_unsigned(574, 12), 187 => to_unsigned(3555, 12), 188 => to_unsigned(2386, 12), 189 => to_unsigned(3837, 12), 190 => to_unsigned(3390, 12), 191 => to_unsigned(1397, 12), 192 => to_unsigned(2467, 12), 193 => to_unsigned(341, 12), 194 => to_unsigned(924, 12), 195 => to_unsigned(955, 12), 196 => to_unsigned(2273, 12), 197 => to_unsigned(1113, 12), 198 => to_unsigned(458, 12), 199 => to_unsigned(1537, 12), 200 => to_unsigned(506, 12), 201 => to_unsigned(3477, 12), 202 => to_unsigned(921, 12), 203 => to_unsigned(3722, 12), 204 => to_unsigned(2680, 12), 205 => to_unsigned(1449, 12), 206 => to_unsigned(1037, 12), 207 => to_unsigned(3763, 12), 208 => to_unsigned(3394, 12), 209 => to_unsigned(2258, 12), 210 => to_unsigned(1236, 12), 211 => to_unsigned(1671, 12), 212 => to_unsigned(2856, 12), 213 => to_unsigned(312, 12), 214 => to_unsigned(341, 12), 215 => to_unsigned(2085, 12), 216 => to_unsigned(1454, 12), 217 => to_unsigned(1235, 12), 218 => to_unsigned(1498, 12), 219 => to_unsigned(1719, 12), 220 => to_unsigned(3462, 12), 221 => to_unsigned(3584, 12), 222 => to_unsigned(1416, 12), 223 => to_unsigned(3068, 12), 224 => to_unsigned(2773, 12), 225 => to_unsigned(3451, 12), 226 => to_unsigned(239, 12), 227 => to_unsigned(677, 12), 228 => to_unsigned(963, 12), 229 => to_unsigned(686, 12), 230 => to_unsigned(744, 12), 231 => to_unsigned(425, 12), 232 => to_unsigned(860, 12), 233 => to_unsigned(3135, 12), 234 => to_unsigned(1081, 12), 235 => to_unsigned(1015, 12), 236 => to_unsigned(3684, 12), 237 => to_unsigned(2599, 12), 238 => to_unsigned(705, 12), 239 => to_unsigned(1459, 12), 240 => to_unsigned(701, 12), 241 => to_unsigned(365, 12), 242 => to_unsigned(1733, 12), 243 => to_unsigned(954, 12), 244 => to_unsigned(3931, 12), 245 => to_unsigned(351, 12), 246 => to_unsigned(936, 12), 247 => to_unsigned(2121, 12), 248 => to_unsigned(2741, 12), 249 => to_unsigned(3960, 12), 250 => to_unsigned(2567, 12), 251 => to_unsigned(355, 12), 252 => to_unsigned(2991, 12), 253 => to_unsigned(709, 12), 254 => to_unsigned(681, 12), 255 => to_unsigned(796, 12), 256 => to_unsigned(3318, 12), 257 => to_unsigned(2938, 12), 258 => to_unsigned(2901, 12), 259 => to_unsigned(779, 12), 260 => to_unsigned(515, 12), 261 => to_unsigned(2322, 12), 262 => to_unsigned(1955, 12), 263 => to_unsigned(46, 12), 264 => to_unsigned(2409, 12), 265 => to_unsigned(3217, 12), 266 => to_unsigned(1135, 12), 267 => to_unsigned(2203, 12), 268 => to_unsigned(1078, 12), 269 => to_unsigned(2671, 12), 270 => to_unsigned(713, 12), 271 => to_unsigned(2451, 12), 272 => to_unsigned(199, 12), 273 => to_unsigned(3655, 12), 274 => to_unsigned(3941, 12), 275 => to_unsigned(3499, 12), 276 => to_unsigned(2046, 12), 277 => to_unsigned(940, 12), 278 => to_unsigned(1646, 12), 279 => to_unsigned(3758, 12), 280 => to_unsigned(2722, 12), 281 => to_unsigned(673, 12), 282 => to_unsigned(2122, 12), 283 => to_unsigned(375, 12), 284 => to_unsigned(2885, 12), 285 => to_unsigned(2524, 12), 286 => to_unsigned(1838, 12), 287 => to_unsigned(928, 12), 288 => to_unsigned(211, 12), 289 => to_unsigned(1447, 12), 290 => to_unsigned(414, 12), 291 => to_unsigned(3295, 12), 292 => to_unsigned(1903, 12), 293 => to_unsigned(1199, 12), 294 => to_unsigned(3969, 12), 295 => to_unsigned(4000, 12), 296 => to_unsigned(894, 12), 297 => to_unsigned(1128, 12), 298 => to_unsigned(2417, 12), 299 => to_unsigned(703, 12), 300 => to_unsigned(1143, 12), 301 => to_unsigned(3373, 12), 302 => to_unsigned(2231, 12), 303 => to_unsigned(1134, 12), 304 => to_unsigned(3958, 12), 305 => to_unsigned(3392, 12), 306 => to_unsigned(869, 12), 307 => to_unsigned(3541, 12), 308 => to_unsigned(3734, 12), 309 => to_unsigned(1435, 12), 310 => to_unsigned(2053, 12), 311 => to_unsigned(3949, 12), 312 => to_unsigned(1059, 12), 313 => to_unsigned(877, 12), 314 => to_unsigned(3875, 12), 315 => to_unsigned(1660, 12), 316 => to_unsigned(616, 12), 317 => to_unsigned(3267, 12), 318 => to_unsigned(3228, 12), 319 => to_unsigned(3675, 12), 320 => to_unsigned(3835, 12), 321 => to_unsigned(2185, 12), 322 => to_unsigned(299, 12), 323 => to_unsigned(1667, 12), 324 => to_unsigned(107, 12), 325 => to_unsigned(3979, 12), 326 => to_unsigned(4019, 12), 327 => to_unsigned(1494, 12), 328 => to_unsigned(2666, 12), 329 => to_unsigned(1770, 12), 330 => to_unsigned(132, 12), 331 => to_unsigned(1693, 12), 332 => to_unsigned(316, 12), 333 => to_unsigned(2476, 12), 334 => to_unsigned(2, 12), 335 => to_unsigned(3038, 12), 336 => to_unsigned(1093, 12), 337 => to_unsigned(1583, 12), 338 => to_unsigned(1228, 12), 339 => to_unsigned(1681, 12), 340 => to_unsigned(2127, 12), 341 => to_unsigned(2744, 12), 342 => to_unsigned(1577, 12), 343 => to_unsigned(920, 12), 344 => to_unsigned(2773, 12), 345 => to_unsigned(3688, 12), 346 => to_unsigned(1539, 12), 347 => to_unsigned(3772, 12), 348 => to_unsigned(3886, 12), 349 => to_unsigned(2416, 12), 350 => to_unsigned(1183, 12), 351 => to_unsigned(454, 12), 352 => to_unsigned(2047, 12), 353 => to_unsigned(3891, 12), 354 => to_unsigned(97, 12), 355 => to_unsigned(3247, 12), 356 => to_unsigned(3339, 12), 357 => to_unsigned(1895, 12), 358 => to_unsigned(1342, 12), 359 => to_unsigned(3720, 12), 360 => to_unsigned(2238, 12), 361 => to_unsigned(3203, 12), 362 => to_unsigned(951, 12), 363 => to_unsigned(2155, 12), 364 => to_unsigned(1846, 12), 365 => to_unsigned(2791, 12), 366 => to_unsigned(169, 12), 367 => to_unsigned(1334, 12), 368 => to_unsigned(281, 12), 369 => to_unsigned(3949, 12), 370 => to_unsigned(2438, 12), 371 => to_unsigned(71, 12), 372 => to_unsigned(3816, 12), 373 => to_unsigned(959, 12), 374 => to_unsigned(1373, 12), 375 => to_unsigned(766, 12), 376 => to_unsigned(4037, 12), 377 => to_unsigned(1574, 12), 378 => to_unsigned(1987, 12), 379 => to_unsigned(1287, 12), 380 => to_unsigned(370, 12), 381 => to_unsigned(4011, 12), 382 => to_unsigned(919, 12), 383 => to_unsigned(3288, 12), 384 => to_unsigned(4082, 12), 385 => to_unsigned(797, 12), 386 => to_unsigned(1331, 12), 387 => to_unsigned(3985, 12), 388 => to_unsigned(1720, 12), 389 => to_unsigned(1323, 12), 390 => to_unsigned(2977, 12), 391 => to_unsigned(2864, 12), 392 => to_unsigned(2766, 12), 393 => to_unsigned(2922, 12), 394 => to_unsigned(426, 12), 395 => to_unsigned(3792, 12), 396 => to_unsigned(239, 12), 397 => to_unsigned(2037, 12), 398 => to_unsigned(3201, 12), 399 => to_unsigned(3434, 12), 400 => to_unsigned(2613, 12), 401 => to_unsigned(1472, 12), 402 => to_unsigned(2803, 12), 403 => to_unsigned(1407, 12), 404 => to_unsigned(1080, 12), 405 => to_unsigned(1167, 12), 406 => to_unsigned(336, 12), 407 => to_unsigned(200, 12), 408 => to_unsigned(361, 12), 409 => to_unsigned(1684, 12), 410 => to_unsigned(1725, 12), 411 => to_unsigned(191, 12), 412 => to_unsigned(2870, 12), 413 => to_unsigned(1451, 12), 414 => to_unsigned(409, 12), 415 => to_unsigned(128, 12), 416 => to_unsigned(2171, 12), 417 => to_unsigned(2353, 12), 418 => to_unsigned(2471, 12), 419 => to_unsigned(386, 12), 420 => to_unsigned(1222, 12), 421 => to_unsigned(2947, 12), 422 => to_unsigned(3870, 12), 423 => to_unsigned(781, 12), 424 => to_unsigned(1812, 12), 425 => to_unsigned(884, 12), 426 => to_unsigned(3403, 12), 427 => to_unsigned(3339, 12), 428 => to_unsigned(2693, 12), 429 => to_unsigned(3952, 12), 430 => to_unsigned(656, 12), 431 => to_unsigned(2509, 12), 432 => to_unsigned(1214, 12), 433 => to_unsigned(3464, 12), 434 => to_unsigned(27, 12), 435 => to_unsigned(902, 12), 436 => to_unsigned(2412, 12), 437 => to_unsigned(3830, 12), 438 => to_unsigned(554, 12), 439 => to_unsigned(2692, 12), 440 => to_unsigned(3048, 12), 441 => to_unsigned(3817, 12), 442 => to_unsigned(399, 12), 443 => to_unsigned(1980, 12), 444 => to_unsigned(3456, 12), 445 => to_unsigned(3239, 12), 446 => to_unsigned(3621, 12), 447 => to_unsigned(518, 12), 448 => to_unsigned(3827, 12), 449 => to_unsigned(605, 12), 450 => to_unsigned(2874, 12), 451 => to_unsigned(1903, 12), 452 => to_unsigned(1945, 12), 453 => to_unsigned(1612, 12), 454 => to_unsigned(2112, 12), 455 => to_unsigned(958, 12), 456 => to_unsigned(4020, 12), 457 => to_unsigned(50, 12), 458 => to_unsigned(177, 12), 459 => to_unsigned(1436, 12), 460 => to_unsigned(1018, 12), 461 => to_unsigned(3015, 12), 462 => to_unsigned(2497, 12), 463 => to_unsigned(3692, 12), 464 => to_unsigned(3824, 12), 465 => to_unsigned(1074, 12), 466 => to_unsigned(2439, 12), 467 => to_unsigned(2024, 12), 468 => to_unsigned(3866, 12), 469 => to_unsigned(3752, 12), 470 => to_unsigned(2365, 12), 471 => to_unsigned(2736, 12), 472 => to_unsigned(494, 12), 473 => to_unsigned(1174, 12), 474 => to_unsigned(782, 12), 475 => to_unsigned(319, 12), 476 => to_unsigned(1503, 12), 477 => to_unsigned(1877, 12), 478 => to_unsigned(564, 12), 479 => to_unsigned(391, 12), 480 => to_unsigned(3108, 12), 481 => to_unsigned(3536, 12), 482 => to_unsigned(3782, 12), 483 => to_unsigned(3306, 12), 484 => to_unsigned(2452, 12), 485 => to_unsigned(2598, 12), 486 => to_unsigned(2436, 12), 487 => to_unsigned(2192, 12), 488 => to_unsigned(1762, 12), 489 => to_unsigned(3183, 12), 490 => to_unsigned(3256, 12), 491 => to_unsigned(251, 12), 492 => to_unsigned(879, 12), 493 => to_unsigned(782, 12), 494 => to_unsigned(1007, 12), 495 => to_unsigned(743, 12), 496 => to_unsigned(3199, 12), 497 => to_unsigned(2063, 12), 498 => to_unsigned(3544, 12), 499 => to_unsigned(654, 12), 500 => to_unsigned(1930, 12), 501 => to_unsigned(758, 12), 502 => to_unsigned(3332, 12), 503 => to_unsigned(596, 12), 504 => to_unsigned(1129, 12), 505 => to_unsigned(2792, 12), 506 => to_unsigned(564, 12), 507 => to_unsigned(3787, 12), 508 => to_unsigned(3324, 12), 509 => to_unsigned(3893, 12), 510 => to_unsigned(1501, 12), 511 => to_unsigned(835, 12), 512 => to_unsigned(2292, 12), 513 => to_unsigned(1836, 12), 514 => to_unsigned(1242, 12), 515 => to_unsigned(3452, 12), 516 => to_unsigned(219, 12), 517 => to_unsigned(1794, 12), 518 => to_unsigned(2236, 12), 519 => to_unsigned(2114, 12), 520 => to_unsigned(2557, 12), 521 => to_unsigned(2583, 12), 522 => to_unsigned(749, 12), 523 => to_unsigned(2076, 12), 524 => to_unsigned(2297, 12), 525 => to_unsigned(2869, 12), 526 => to_unsigned(2962, 12), 527 => to_unsigned(1903, 12), 528 => to_unsigned(4027, 12), 529 => to_unsigned(3649, 12), 530 => to_unsigned(1092, 12), 531 => to_unsigned(1060, 12), 532 => to_unsigned(1873, 12), 533 => to_unsigned(1048, 12), 534 => to_unsigned(2777, 12), 535 => to_unsigned(3947, 12), 536 => to_unsigned(3404, 12), 537 => to_unsigned(290, 12), 538 => to_unsigned(3413, 12), 539 => to_unsigned(2872, 12), 540 => to_unsigned(2034, 12), 541 => to_unsigned(3647, 12), 542 => to_unsigned(1993, 12), 543 => to_unsigned(1316, 12), 544 => to_unsigned(3947, 12), 545 => to_unsigned(2473, 12), 546 => to_unsigned(262, 12), 547 => to_unsigned(2961, 12), 548 => to_unsigned(2335, 12), 549 => to_unsigned(506, 12), 550 => to_unsigned(1650, 12), 551 => to_unsigned(2287, 12), 552 => to_unsigned(1004, 12), 553 => to_unsigned(3590, 12), 554 => to_unsigned(178, 12), 555 => to_unsigned(784, 12), 556 => to_unsigned(3870, 12), 557 => to_unsigned(3868, 12), 558 => to_unsigned(3199, 12), 559 => to_unsigned(459, 12), 560 => to_unsigned(160, 12), 561 => to_unsigned(1894, 12), 562 => to_unsigned(473, 12), 563 => to_unsigned(550, 12), 564 => to_unsigned(2333, 12), 565 => to_unsigned(3330, 12), 566 => to_unsigned(1619, 12), 567 => to_unsigned(332, 12), 568 => to_unsigned(1938, 12), 569 => to_unsigned(1088, 12), 570 => to_unsigned(2473, 12), 571 => to_unsigned(1174, 12), 572 => to_unsigned(2577, 12), 573 => to_unsigned(682, 12), 574 => to_unsigned(2052, 12), 575 => to_unsigned(2180, 12), 576 => to_unsigned(1426, 12), 577 => to_unsigned(2757, 12), 578 => to_unsigned(2062, 12), 579 => to_unsigned(10, 12), 580 => to_unsigned(306, 12), 581 => to_unsigned(989, 12), 582 => to_unsigned(2771, 12), 583 => to_unsigned(2850, 12), 584 => to_unsigned(3, 12), 585 => to_unsigned(3080, 12), 586 => to_unsigned(3034, 12), 587 => to_unsigned(1618, 12), 588 => to_unsigned(3652, 12), 589 => to_unsigned(2695, 12), 590 => to_unsigned(2410, 12), 591 => to_unsigned(3421, 12), 592 => to_unsigned(3107, 12), 593 => to_unsigned(3791, 12), 594 => to_unsigned(1070, 12), 595 => to_unsigned(3245, 12), 596 => to_unsigned(2499, 12), 597 => to_unsigned(570, 12), 598 => to_unsigned(643, 12), 599 => to_unsigned(2246, 12), 600 => to_unsigned(3138, 12), 601 => to_unsigned(3045, 12), 602 => to_unsigned(664, 12), 603 => to_unsigned(1719, 12), 604 => to_unsigned(2491, 12), 605 => to_unsigned(1699, 12), 606 => to_unsigned(1283, 12), 607 => to_unsigned(3655, 12), 608 => to_unsigned(3995, 12), 609 => to_unsigned(3058, 12), 610 => to_unsigned(2882, 12), 611 => to_unsigned(1534, 12), 612 => to_unsigned(2416, 12), 613 => to_unsigned(583, 12), 614 => to_unsigned(3082, 12), 615 => to_unsigned(2157, 12), 616 => to_unsigned(1215, 12), 617 => to_unsigned(3451, 12), 618 => to_unsigned(2160, 12), 619 => to_unsigned(1401, 12), 620 => to_unsigned(5, 12), 621 => to_unsigned(3572, 12), 622 => to_unsigned(3368, 12), 623 => to_unsigned(4054, 12), 624 => to_unsigned(436, 12), 625 => to_unsigned(1963, 12), 626 => to_unsigned(3521, 12), 627 => to_unsigned(902, 12), 628 => to_unsigned(3868, 12), 629 => to_unsigned(389, 12), 630 => to_unsigned(232, 12), 631 => to_unsigned(1610, 12), 632 => to_unsigned(647, 12), 633 => to_unsigned(1821, 12), 634 => to_unsigned(2916, 12), 635 => to_unsigned(338, 12), 636 => to_unsigned(47, 12), 637 => to_unsigned(2492, 12), 638 => to_unsigned(2367, 12), 639 => to_unsigned(2683, 12), 640 => to_unsigned(2498, 12), 641 => to_unsigned(297, 12), 642 => to_unsigned(1565, 12), 643 => to_unsigned(1120, 12), 644 => to_unsigned(3633, 12), 645 => to_unsigned(2748, 12), 646 => to_unsigned(820, 12), 647 => to_unsigned(537, 12), 648 => to_unsigned(3620, 12), 649 => to_unsigned(659, 12), 650 => to_unsigned(3936, 12), 651 => to_unsigned(1269, 12), 652 => to_unsigned(603, 12), 653 => to_unsigned(3226, 12), 654 => to_unsigned(3640, 12), 655 => to_unsigned(3384, 12), 656 => to_unsigned(3868, 12), 657 => to_unsigned(4013, 12), 658 => to_unsigned(3031, 12), 659 => to_unsigned(466, 12), 660 => to_unsigned(3333, 12), 661 => to_unsigned(961, 12), 662 => to_unsigned(2645, 12), 663 => to_unsigned(3362, 12), 664 => to_unsigned(897, 12), 665 => to_unsigned(605, 12), 666 => to_unsigned(1773, 12), 667 => to_unsigned(2018, 12), 668 => to_unsigned(2318, 12), 669 => to_unsigned(234, 12), 670 => to_unsigned(1566, 12), 671 => to_unsigned(1929, 12), 672 => to_unsigned(2486, 12), 673 => to_unsigned(3867, 12), 674 => to_unsigned(391, 12), 675 => to_unsigned(4044, 12), 676 => to_unsigned(3421, 12), 677 => to_unsigned(3748, 12), 678 => to_unsigned(166, 12), 679 => to_unsigned(92, 12), 680 => to_unsigned(3697, 12), 681 => to_unsigned(1621, 12), 682 => to_unsigned(2263, 12), 683 => to_unsigned(1445, 12), 684 => to_unsigned(3988, 12), 685 => to_unsigned(781, 12), 686 => to_unsigned(109, 12), 687 => to_unsigned(1704, 12), 688 => to_unsigned(3506, 12), 689 => to_unsigned(3561, 12), 690 => to_unsigned(2358, 12), 691 => to_unsigned(3198, 12), 692 => to_unsigned(1473, 12), 693 => to_unsigned(2888, 12), 694 => to_unsigned(58, 12), 695 => to_unsigned(2151, 12), 696 => to_unsigned(876, 12), 697 => to_unsigned(1097, 12), 698 => to_unsigned(2609, 12), 699 => to_unsigned(273, 12), 700 => to_unsigned(305, 12), 701 => to_unsigned(1113, 12), 702 => to_unsigned(2519, 12), 703 => to_unsigned(3001, 12), 704 => to_unsigned(3048, 12), 705 => to_unsigned(249, 12), 706 => to_unsigned(115, 12), 707 => to_unsigned(714, 12), 708 => to_unsigned(2906, 12), 709 => to_unsigned(3341, 12), 710 => to_unsigned(2335, 12), 711 => to_unsigned(3196, 12), 712 => to_unsigned(3605, 12), 713 => to_unsigned(865, 12), 714 => to_unsigned(2541, 12), 715 => to_unsigned(2305, 12), 716 => to_unsigned(1504, 12), 717 => to_unsigned(2219, 12), 718 => to_unsigned(2743, 12), 719 => to_unsigned(838, 12), 720 => to_unsigned(3362, 12), 721 => to_unsigned(990, 12), 722 => to_unsigned(2606, 12), 723 => to_unsigned(2394, 12), 724 => to_unsigned(1510, 12), 725 => to_unsigned(3044, 12), 726 => to_unsigned(657, 12), 727 => to_unsigned(2928, 12), 728 => to_unsigned(1292, 12), 729 => to_unsigned(3636, 12), 730 => to_unsigned(2863, 12), 731 => to_unsigned(1396, 12), 732 => to_unsigned(935, 12), 733 => to_unsigned(1904, 12), 734 => to_unsigned(2992, 12), 735 => to_unsigned(4023, 12), 736 => to_unsigned(2713, 12), 737 => to_unsigned(2880, 12), 738 => to_unsigned(316, 12), 739 => to_unsigned(998, 12), 740 => to_unsigned(1182, 12), 741 => to_unsigned(2281, 12), 742 => to_unsigned(1775, 12), 743 => to_unsigned(3172, 12), 744 => to_unsigned(3686, 12), 745 => to_unsigned(2908, 12), 746 => to_unsigned(2538, 12), 747 => to_unsigned(3799, 12), 748 => to_unsigned(2639, 12), 749 => to_unsigned(422, 12), 750 => to_unsigned(3430, 12), 751 => to_unsigned(4054, 12), 752 => to_unsigned(3888, 12), 753 => to_unsigned(1287, 12), 754 => to_unsigned(2597, 12), 755 => to_unsigned(2290, 12), 756 => to_unsigned(1858, 12), 757 => to_unsigned(2125, 12), 758 => to_unsigned(1300, 12), 759 => to_unsigned(2862, 12), 760 => to_unsigned(477, 12), 761 => to_unsigned(288, 12), 762 => to_unsigned(1844, 12), 763 => to_unsigned(2487, 12), 764 => to_unsigned(3475, 12), 765 => to_unsigned(2028, 12), 766 => to_unsigned(3052, 12), 767 => to_unsigned(2488, 12), 768 => to_unsigned(3606, 12), 769 => to_unsigned(86, 12), 770 => to_unsigned(2540, 12), 771 => to_unsigned(2277, 12), 772 => to_unsigned(2620, 12), 773 => to_unsigned(2722, 12), 774 => to_unsigned(573, 12), 775 => to_unsigned(950, 12), 776 => to_unsigned(1062, 12), 777 => to_unsigned(3797, 12), 778 => to_unsigned(988, 12), 779 => to_unsigned(688, 12), 780 => to_unsigned(418, 12), 781 => to_unsigned(3005, 12), 782 => to_unsigned(1729, 12), 783 => to_unsigned(3254, 12), 784 => to_unsigned(2925, 12), 785 => to_unsigned(2286, 12), 786 => to_unsigned(145, 12), 787 => to_unsigned(2612, 12), 788 => to_unsigned(2338, 12), 789 => to_unsigned(4011, 12), 790 => to_unsigned(141, 12), 791 => to_unsigned(17, 12), 792 => to_unsigned(3871, 12), 793 => to_unsigned(1557, 12), 794 => to_unsigned(226, 12), 795 => to_unsigned(3693, 12), 796 => to_unsigned(3713, 12), 797 => to_unsigned(3653, 12), 798 => to_unsigned(943, 12), 799 => to_unsigned(3314, 12), 800 => to_unsigned(1190, 12), 801 => to_unsigned(3903, 12), 802 => to_unsigned(1183, 12), 803 => to_unsigned(860, 12), 804 => to_unsigned(2150, 12), 805 => to_unsigned(2810, 12), 806 => to_unsigned(114, 12), 807 => to_unsigned(1264, 12), 808 => to_unsigned(1860, 12), 809 => to_unsigned(2469, 12), 810 => to_unsigned(3975, 12), 811 => to_unsigned(579, 12), 812 => to_unsigned(3126, 12), 813 => to_unsigned(2069, 12), 814 => to_unsigned(2197, 12), 815 => to_unsigned(3385, 12), 816 => to_unsigned(986, 12), 817 => to_unsigned(2370, 12), 818 => to_unsigned(3804, 12), 819 => to_unsigned(2863, 12), 820 => to_unsigned(1056, 12), 821 => to_unsigned(229, 12), 822 => to_unsigned(1697, 12), 823 => to_unsigned(1251, 12), 824 => to_unsigned(1978, 12), 825 => to_unsigned(928, 12), 826 => to_unsigned(1639, 12), 827 => to_unsigned(1169, 12), 828 => to_unsigned(905, 12), 829 => to_unsigned(2659, 12), 830 => to_unsigned(1964, 12), 831 => to_unsigned(2646, 12), 832 => to_unsigned(2309, 12), 833 => to_unsigned(4054, 12), 834 => to_unsigned(3721, 12), 835 => to_unsigned(2166, 12), 836 => to_unsigned(321, 12), 837 => to_unsigned(2749, 12), 838 => to_unsigned(235, 12), 839 => to_unsigned(133, 12), 840 => to_unsigned(2282, 12), 841 => to_unsigned(196, 12), 842 => to_unsigned(2695, 12), 843 => to_unsigned(950, 12), 844 => to_unsigned(19, 12), 845 => to_unsigned(2034, 12), 846 => to_unsigned(2867, 12), 847 => to_unsigned(2982, 12), 848 => to_unsigned(4085, 12), 849 => to_unsigned(2807, 12), 850 => to_unsigned(653, 12), 851 => to_unsigned(11, 12), 852 => to_unsigned(855, 12), 853 => to_unsigned(1382, 12), 854 => to_unsigned(566, 12), 855 => to_unsigned(3253, 12), 856 => to_unsigned(587, 12), 857 => to_unsigned(2344, 12), 858 => to_unsigned(2037, 12), 859 => to_unsigned(607, 12), 860 => to_unsigned(515, 12), 861 => to_unsigned(503, 12), 862 => to_unsigned(3773, 12), 863 => to_unsigned(1154, 12), 864 => to_unsigned(1991, 12), 865 => to_unsigned(258, 12), 866 => to_unsigned(281, 12), 867 => to_unsigned(3886, 12), 868 => to_unsigned(1413, 12), 869 => to_unsigned(2064, 12), 870 => to_unsigned(1138, 12), 871 => to_unsigned(136, 12), 872 => to_unsigned(721, 12), 873 => to_unsigned(1144, 12), 874 => to_unsigned(3442, 12), 875 => to_unsigned(3676, 12), 876 => to_unsigned(590, 12), 877 => to_unsigned(3512, 12), 878 => to_unsigned(2566, 12), 879 => to_unsigned(589, 12), 880 => to_unsigned(568, 12), 881 => to_unsigned(3036, 12), 882 => to_unsigned(1795, 12), 883 => to_unsigned(3564, 12), 884 => to_unsigned(1339, 12), 885 => to_unsigned(3686, 12), 886 => to_unsigned(2415, 12), 887 => to_unsigned(3076, 12), 888 => to_unsigned(1024, 12), 889 => to_unsigned(3787, 12), 890 => to_unsigned(934, 12), 891 => to_unsigned(3206, 12), 892 => to_unsigned(1907, 12), 893 => to_unsigned(1684, 12), 894 => to_unsigned(2552, 12), 895 => to_unsigned(2758, 12), 896 => to_unsigned(3984, 12), 897 => to_unsigned(832, 12), 898 => to_unsigned(323, 12), 899 => to_unsigned(3195, 12), 900 => to_unsigned(3141, 12), 901 => to_unsigned(367, 12), 902 => to_unsigned(61, 12), 903 => to_unsigned(2343, 12), 904 => to_unsigned(1339, 12), 905 => to_unsigned(208, 12), 906 => to_unsigned(473, 12), 907 => to_unsigned(505, 12), 908 => to_unsigned(4062, 12), 909 => to_unsigned(3355, 12), 910 => to_unsigned(3275, 12), 911 => to_unsigned(3048, 12), 912 => to_unsigned(960, 12), 913 => to_unsigned(289, 12), 914 => to_unsigned(1305, 12), 915 => to_unsigned(692, 12), 916 => to_unsigned(3982, 12), 917 => to_unsigned(688, 12), 918 => to_unsigned(2466, 12), 919 => to_unsigned(1652, 12), 920 => to_unsigned(1576, 12), 921 => to_unsigned(946, 12), 922 => to_unsigned(2750, 12), 923 => to_unsigned(3186, 12), 924 => to_unsigned(3371, 12), 925 => to_unsigned(1655, 12), 926 => to_unsigned(2086, 12), 927 => to_unsigned(2195, 12), 928 => to_unsigned(3882, 12), 929 => to_unsigned(2530, 12), 930 => to_unsigned(3814, 12), 931 => to_unsigned(1173, 12), 932 => to_unsigned(3988, 12), 933 => to_unsigned(3418, 12), 934 => to_unsigned(419, 12), 935 => to_unsigned(3995, 12), 936 => to_unsigned(2691, 12), 937 => to_unsigned(3033, 12), 938 => to_unsigned(2940, 12), 939 => to_unsigned(391, 12), 940 => to_unsigned(3332, 12), 941 => to_unsigned(516, 12), 942 => to_unsigned(2101, 12), 943 => to_unsigned(393, 12), 944 => to_unsigned(964, 12), 945 => to_unsigned(2721, 12), 946 => to_unsigned(2993, 12), 947 => to_unsigned(3786, 12), 948 => to_unsigned(1943, 12), 949 => to_unsigned(3001, 12), 950 => to_unsigned(2800, 12), 951 => to_unsigned(3040, 12), 952 => to_unsigned(3917, 12), 953 => to_unsigned(3477, 12), 954 => to_unsigned(92, 12), 955 => to_unsigned(3095, 12), 956 => to_unsigned(112, 12), 957 => to_unsigned(3461, 12), 958 => to_unsigned(1981, 12), 959 => to_unsigned(2050, 12), 960 => to_unsigned(3328, 12), 961 => to_unsigned(1801, 12), 962 => to_unsigned(1863, 12), 963 => to_unsigned(3997, 12), 964 => to_unsigned(149, 12), 965 => to_unsigned(1488, 12), 966 => to_unsigned(590, 12), 967 => to_unsigned(2003, 12), 968 => to_unsigned(3621, 12), 969 => to_unsigned(3674, 12), 970 => to_unsigned(1100, 12), 971 => to_unsigned(1359, 12), 972 => to_unsigned(723, 12), 973 => to_unsigned(3218, 12), 974 => to_unsigned(3562, 12), 975 => to_unsigned(1602, 12), 976 => to_unsigned(784, 12), 977 => to_unsigned(3064, 12), 978 => to_unsigned(331, 12), 979 => to_unsigned(4067, 12), 980 => to_unsigned(3593, 12), 981 => to_unsigned(377, 12), 982 => to_unsigned(1353, 12), 983 => to_unsigned(3870, 12), 984 => to_unsigned(1046, 12), 985 => to_unsigned(3690, 12), 986 => to_unsigned(2324, 12), 987 => to_unsigned(617, 12), 988 => to_unsigned(2515, 12), 989 => to_unsigned(1348, 12), 990 => to_unsigned(3438, 12), 991 => to_unsigned(1103, 12), 992 => to_unsigned(1441, 12), 993 => to_unsigned(3008, 12), 994 => to_unsigned(879, 12), 995 => to_unsigned(3983, 12), 996 => to_unsigned(3405, 12), 997 => to_unsigned(905, 12), 998 => to_unsigned(3121, 12), 999 => to_unsigned(2794, 12), 1000 => to_unsigned(3210, 12), 1001 => to_unsigned(369, 12), 1002 => to_unsigned(615, 12), 1003 => to_unsigned(2594, 12), 1004 => to_unsigned(1959, 12), 1005 => to_unsigned(1968, 12), 1006 => to_unsigned(1324, 12), 1007 => to_unsigned(3820, 12), 1008 => to_unsigned(618, 12), 1009 => to_unsigned(2305, 12), 1010 => to_unsigned(1992, 12), 1011 => to_unsigned(1280, 12), 1012 => to_unsigned(2187, 12), 1013 => to_unsigned(2970, 12), 1014 => to_unsigned(478, 12), 1015 => to_unsigned(1899, 12), 1016 => to_unsigned(4010, 12), 1017 => to_unsigned(2835, 12), 1018 => to_unsigned(853, 12), 1019 => to_unsigned(3951, 12), 1020 => to_unsigned(1793, 12), 1021 => to_unsigned(1530, 12), 1022 => to_unsigned(956, 12), 1023 => to_unsigned(594, 12), 1024 => to_unsigned(3548, 12), 1025 => to_unsigned(3646, 12), 1026 => to_unsigned(3979, 12), 1027 => to_unsigned(3067, 12), 1028 => to_unsigned(2737, 12), 1029 => to_unsigned(3263, 12), 1030 => to_unsigned(884, 12), 1031 => to_unsigned(615, 12), 1032 => to_unsigned(3721, 12), 1033 => to_unsigned(1048, 12), 1034 => to_unsigned(2116, 12), 1035 => to_unsigned(2842, 12), 1036 => to_unsigned(3892, 12), 1037 => to_unsigned(3179, 12), 1038 => to_unsigned(2614, 12), 1039 => to_unsigned(2517, 12), 1040 => to_unsigned(3790, 12), 1041 => to_unsigned(3229, 12), 1042 => to_unsigned(3969, 12), 1043 => to_unsigned(1230, 12), 1044 => to_unsigned(2304, 12), 1045 => to_unsigned(2575, 12), 1046 => to_unsigned(3489, 12), 1047 => to_unsigned(672, 12), 1048 => to_unsigned(765, 12), 1049 => to_unsigned(755, 12), 1050 => to_unsigned(2789, 12), 1051 => to_unsigned(197, 12), 1052 => to_unsigned(1950, 12), 1053 => to_unsigned(3574, 12), 1054 => to_unsigned(3177, 12), 1055 => to_unsigned(687, 12), 1056 => to_unsigned(1522, 12), 1057 => to_unsigned(3642, 12), 1058 => to_unsigned(4041, 12), 1059 => to_unsigned(373, 12), 1060 => to_unsigned(2951, 12), 1061 => to_unsigned(2046, 12), 1062 => to_unsigned(2974, 12), 1063 => to_unsigned(3413, 12), 1064 => to_unsigned(1054, 12), 1065 => to_unsigned(2473, 12), 1066 => to_unsigned(3080, 12), 1067 => to_unsigned(2113, 12), 1068 => to_unsigned(3693, 12), 1069 => to_unsigned(3541, 12), 1070 => to_unsigned(3336, 12), 1071 => to_unsigned(3321, 12), 1072 => to_unsigned(749, 12), 1073 => to_unsigned(1073, 12), 1074 => to_unsigned(372, 12), 1075 => to_unsigned(2112, 12), 1076 => to_unsigned(2651, 12), 1077 => to_unsigned(2098, 12), 1078 => to_unsigned(3248, 12), 1079 => to_unsigned(3545, 12), 1080 => to_unsigned(2717, 12), 1081 => to_unsigned(583, 12), 1082 => to_unsigned(1562, 12), 1083 => to_unsigned(1503, 12), 1084 => to_unsigned(3470, 12), 1085 => to_unsigned(2937, 12), 1086 => to_unsigned(2835, 12), 1087 => to_unsigned(1150, 12), 1088 => to_unsigned(2184, 12), 1089 => to_unsigned(3111, 12), 1090 => to_unsigned(925, 12), 1091 => to_unsigned(3351, 12), 1092 => to_unsigned(3917, 12), 1093 => to_unsigned(40, 12), 1094 => to_unsigned(3201, 12), 1095 => to_unsigned(857, 12), 1096 => to_unsigned(1496, 12), 1097 => to_unsigned(798, 12), 1098 => to_unsigned(1449, 12), 1099 => to_unsigned(2896, 12), 1100 => to_unsigned(1404, 12), 1101 => to_unsigned(2878, 12), 1102 => to_unsigned(3915, 12), 1103 => to_unsigned(1895, 12), 1104 => to_unsigned(1863, 12), 1105 => to_unsigned(1638, 12), 1106 => to_unsigned(3541, 12), 1107 => to_unsigned(4056, 12), 1108 => to_unsigned(1317, 12), 1109 => to_unsigned(2859, 12), 1110 => to_unsigned(2491, 12), 1111 => to_unsigned(3748, 12), 1112 => to_unsigned(672, 12), 1113 => to_unsigned(2889, 12), 1114 => to_unsigned(753, 12), 1115 => to_unsigned(767, 12), 1116 => to_unsigned(2024, 12), 1117 => to_unsigned(2960, 12), 1118 => to_unsigned(3491, 12), 1119 => to_unsigned(3831, 12), 1120 => to_unsigned(387, 12), 1121 => to_unsigned(1575, 12), 1122 => to_unsigned(421, 12), 1123 => to_unsigned(1530, 12), 1124 => to_unsigned(3331, 12), 1125 => to_unsigned(3496, 12), 1126 => to_unsigned(2618, 12), 1127 => to_unsigned(3555, 12), 1128 => to_unsigned(3713, 12), 1129 => to_unsigned(515, 12), 1130 => to_unsigned(523, 12), 1131 => to_unsigned(3459, 12), 1132 => to_unsigned(1134, 12), 1133 => to_unsigned(3582, 12), 1134 => to_unsigned(2747, 12), 1135 => to_unsigned(1164, 12), 1136 => to_unsigned(1888, 12), 1137 => to_unsigned(1959, 12), 1138 => to_unsigned(2866, 12), 1139 => to_unsigned(2816, 12), 1140 => to_unsigned(566, 12), 1141 => to_unsigned(1078, 12), 1142 => to_unsigned(3695, 12), 1143 => to_unsigned(1879, 12), 1144 => to_unsigned(711, 12), 1145 => to_unsigned(1723, 12), 1146 => to_unsigned(3393, 12), 1147 => to_unsigned(482, 12), 1148 => to_unsigned(1805, 12), 1149 => to_unsigned(4024, 12), 1150 => to_unsigned(1054, 12), 1151 => to_unsigned(3413, 12), 1152 => to_unsigned(3665, 12), 1153 => to_unsigned(663, 12), 1154 => to_unsigned(2979, 12), 1155 => to_unsigned(929, 12), 1156 => to_unsigned(902, 12), 1157 => to_unsigned(2072, 12), 1158 => to_unsigned(1058, 12), 1159 => to_unsigned(3063, 12), 1160 => to_unsigned(1640, 12), 1161 => to_unsigned(441, 12), 1162 => to_unsigned(358, 12), 1163 => to_unsigned(457, 12), 1164 => to_unsigned(664, 12), 1165 => to_unsigned(1757, 12), 1166 => to_unsigned(1541, 12), 1167 => to_unsigned(1264, 12), 1168 => to_unsigned(2992, 12), 1169 => to_unsigned(2969, 12), 1170 => to_unsigned(1476, 12), 1171 => to_unsigned(1774, 12), 1172 => to_unsigned(2086, 12), 1173 => to_unsigned(2432, 12), 1174 => to_unsigned(3387, 12), 1175 => to_unsigned(2254, 12), 1176 => to_unsigned(3145, 12), 1177 => to_unsigned(2276, 12), 1178 => to_unsigned(3567, 12), 1179 => to_unsigned(1970, 12), 1180 => to_unsigned(28, 12), 1181 => to_unsigned(1423, 12), 1182 => to_unsigned(706, 12), 1183 => to_unsigned(3108, 12), 1184 => to_unsigned(647, 12), 1185 => to_unsigned(2001, 12), 1186 => to_unsigned(1695, 12), 1187 => to_unsigned(3243, 12), 1188 => to_unsigned(41, 12), 1189 => to_unsigned(1487, 12), 1190 => to_unsigned(2844, 12), 1191 => to_unsigned(382, 12), 1192 => to_unsigned(182, 12), 1193 => to_unsigned(1844, 12), 1194 => to_unsigned(2166, 12), 1195 => to_unsigned(2730, 12), 1196 => to_unsigned(1784, 12), 1197 => to_unsigned(1439, 12), 1198 => to_unsigned(86, 12), 1199 => to_unsigned(2617, 12), 1200 => to_unsigned(2546, 12), 1201 => to_unsigned(3095, 12), 1202 => to_unsigned(1148, 12), 1203 => to_unsigned(836, 12), 1204 => to_unsigned(2624, 12), 1205 => to_unsigned(3985, 12), 1206 => to_unsigned(2246, 12), 1207 => to_unsigned(2116, 12), 1208 => to_unsigned(3275, 12), 1209 => to_unsigned(2016, 12), 1210 => to_unsigned(1232, 12), 1211 => to_unsigned(3970, 12), 1212 => to_unsigned(3578, 12), 1213 => to_unsigned(2762, 12), 1214 => to_unsigned(3495, 12), 1215 => to_unsigned(510, 12), 1216 => to_unsigned(3238, 12), 1217 => to_unsigned(1462, 12), 1218 => to_unsigned(3836, 12), 1219 => to_unsigned(1639, 12), 1220 => to_unsigned(1021, 12), 1221 => to_unsigned(1271, 12), 1222 => to_unsigned(128, 12), 1223 => to_unsigned(2825, 12), 1224 => to_unsigned(1611, 12), 1225 => to_unsigned(3500, 12), 1226 => to_unsigned(1076, 12), 1227 => to_unsigned(1233, 12), 1228 => to_unsigned(3428, 12), 1229 => to_unsigned(1385, 12), 1230 => to_unsigned(687, 12), 1231 => to_unsigned(2757, 12), 1232 => to_unsigned(3561, 12), 1233 => to_unsigned(3632, 12), 1234 => to_unsigned(3494, 12), 1235 => to_unsigned(2084, 12), 1236 => to_unsigned(1412, 12), 1237 => to_unsigned(1787, 12), 1238 => to_unsigned(1009, 12), 1239 => to_unsigned(2251, 12), 1240 => to_unsigned(3111, 12), 1241 => to_unsigned(221, 12), 1242 => to_unsigned(747, 12), 1243 => to_unsigned(190, 12), 1244 => to_unsigned(685, 12), 1245 => to_unsigned(2507, 12), 1246 => to_unsigned(1834, 12), 1247 => to_unsigned(2208, 12), 1248 => to_unsigned(897, 12), 1249 => to_unsigned(748, 12), 1250 => to_unsigned(1199, 12), 1251 => to_unsigned(3746, 12), 1252 => to_unsigned(3370, 12), 1253 => to_unsigned(1322, 12), 1254 => to_unsigned(364, 12), 1255 => to_unsigned(3274, 12), 1256 => to_unsigned(426, 12), 1257 => to_unsigned(3836, 12), 1258 => to_unsigned(1768, 12), 1259 => to_unsigned(3630, 12), 1260 => to_unsigned(999, 12), 1261 => to_unsigned(3535, 12), 1262 => to_unsigned(2669, 12), 1263 => to_unsigned(3802, 12), 1264 => to_unsigned(1641, 12), 1265 => to_unsigned(1576, 12), 1266 => to_unsigned(2668, 12), 1267 => to_unsigned(368, 12), 1268 => to_unsigned(1872, 12), 1269 => to_unsigned(3499, 12), 1270 => to_unsigned(2908, 12), 1271 => to_unsigned(448, 12), 1272 => to_unsigned(1599, 12), 1273 => to_unsigned(1068, 12), 1274 => to_unsigned(2941, 12), 1275 => to_unsigned(2690, 12), 1276 => to_unsigned(3606, 12), 1277 => to_unsigned(3452, 12), 1278 => to_unsigned(1944, 12), 1279 => to_unsigned(4012, 12), 1280 => to_unsigned(3923, 12), 1281 => to_unsigned(3806, 12), 1282 => to_unsigned(1997, 12), 1283 => to_unsigned(1415, 12), 1284 => to_unsigned(3283, 12), 1285 => to_unsigned(2275, 12), 1286 => to_unsigned(309, 12), 1287 => to_unsigned(501, 12), 1288 => to_unsigned(3390, 12), 1289 => to_unsigned(1437, 12), 1290 => to_unsigned(724, 12), 1291 => to_unsigned(3592, 12), 1292 => to_unsigned(970, 12), 1293 => to_unsigned(809, 12), 1294 => to_unsigned(930, 12), 1295 => to_unsigned(1198, 12), 1296 => to_unsigned(3005, 12), 1297 => to_unsigned(2763, 12), 1298 => to_unsigned(3325, 12), 1299 => to_unsigned(712, 12), 1300 => to_unsigned(1653, 12), 1301 => to_unsigned(1335, 12), 1302 => to_unsigned(4053, 12), 1303 => to_unsigned(1780, 12), 1304 => to_unsigned(2628, 12), 1305 => to_unsigned(303, 12), 1306 => to_unsigned(2567, 12), 1307 => to_unsigned(248, 12), 1308 => to_unsigned(312, 12), 1309 => to_unsigned(85, 12), 1310 => to_unsigned(1110, 12), 1311 => to_unsigned(3398, 12), 1312 => to_unsigned(19, 12), 1313 => to_unsigned(3755, 12), 1314 => to_unsigned(1350, 12), 1315 => to_unsigned(1376, 12), 1316 => to_unsigned(3579, 12), 1317 => to_unsigned(357, 12), 1318 => to_unsigned(1366, 12), 1319 => to_unsigned(2409, 12), 1320 => to_unsigned(3861, 12), 1321 => to_unsigned(1780, 12), 1322 => to_unsigned(3211, 12), 1323 => to_unsigned(1195, 12), 1324 => to_unsigned(67, 12), 1325 => to_unsigned(1760, 12), 1326 => to_unsigned(925, 12), 1327 => to_unsigned(2965, 12), 1328 => to_unsigned(1233, 12), 1329 => to_unsigned(3397, 12), 1330 => to_unsigned(3823, 12), 1331 => to_unsigned(2523, 12), 1332 => to_unsigned(2305, 12), 1333 => to_unsigned(2721, 12), 1334 => to_unsigned(3496, 12), 1335 => to_unsigned(1387, 12), 1336 => to_unsigned(1127, 12), 1337 => to_unsigned(2809, 12), 1338 => to_unsigned(1707, 12), 1339 => to_unsigned(2099, 12), 1340 => to_unsigned(3045, 12), 1341 => to_unsigned(3422, 12), 1342 => to_unsigned(466, 12), 1343 => to_unsigned(2486, 12), 1344 => to_unsigned(1999, 12), 1345 => to_unsigned(3836, 12), 1346 => to_unsigned(307, 12), 1347 => to_unsigned(2477, 12), 1348 => to_unsigned(1256, 12), 1349 => to_unsigned(3421, 12), 1350 => to_unsigned(132, 12), 1351 => to_unsigned(2744, 12), 1352 => to_unsigned(3504, 12), 1353 => to_unsigned(1912, 12), 1354 => to_unsigned(490, 12), 1355 => to_unsigned(2452, 12), 1356 => to_unsigned(784, 12), 1357 => to_unsigned(1077, 12), 1358 => to_unsigned(2005, 12), 1359 => to_unsigned(706, 12), 1360 => to_unsigned(1428, 12), 1361 => to_unsigned(4077, 12), 1362 => to_unsigned(952, 12), 1363 => to_unsigned(408, 12), 1364 => to_unsigned(3883, 12), 1365 => to_unsigned(3412, 12), 1366 => to_unsigned(749, 12), 1367 => to_unsigned(1727, 12), 1368 => to_unsigned(1039, 12), 1369 => to_unsigned(3425, 12), 1370 => to_unsigned(2328, 12), 1371 => to_unsigned(3416, 12), 1372 => to_unsigned(2408, 12), 1373 => to_unsigned(3675, 12), 1374 => to_unsigned(3389, 12), 1375 => to_unsigned(643, 12), 1376 => to_unsigned(2451, 12), 1377 => to_unsigned(652, 12), 1378 => to_unsigned(114, 12), 1379 => to_unsigned(3372, 12), 1380 => to_unsigned(1866, 12), 1381 => to_unsigned(2441, 12), 1382 => to_unsigned(2751, 12), 1383 => to_unsigned(988, 12), 1384 => to_unsigned(373, 12), 1385 => to_unsigned(3758, 12), 1386 => to_unsigned(1759, 12), 1387 => to_unsigned(3543, 12), 1388 => to_unsigned(3981, 12), 1389 => to_unsigned(3653, 12), 1390 => to_unsigned(3757, 12), 1391 => to_unsigned(2024, 12), 1392 => to_unsigned(3207, 12), 1393 => to_unsigned(1321, 12), 1394 => to_unsigned(622, 12), 1395 => to_unsigned(400, 12), 1396 => to_unsigned(1202, 12), 1397 => to_unsigned(2855, 12), 1398 => to_unsigned(2083, 12), 1399 => to_unsigned(1898, 12), 1400 => to_unsigned(2332, 12), 1401 => to_unsigned(1653, 12), 1402 => to_unsigned(1105, 12), 1403 => to_unsigned(2085, 12), 1404 => to_unsigned(513, 12), 1405 => to_unsigned(2513, 12), 1406 => to_unsigned(2334, 12), 1407 => to_unsigned(3106, 12), 1408 => to_unsigned(3956, 12), 1409 => to_unsigned(1027, 12), 1410 => to_unsigned(3489, 12), 1411 => to_unsigned(2219, 12), 1412 => to_unsigned(3417, 12), 1413 => to_unsigned(1537, 12), 1414 => to_unsigned(354, 12), 1415 => to_unsigned(3512, 12), 1416 => to_unsigned(1841, 12), 1417 => to_unsigned(3175, 12), 1418 => to_unsigned(808, 12), 1419 => to_unsigned(3154, 12), 1420 => to_unsigned(553, 12), 1421 => to_unsigned(310, 12), 1422 => to_unsigned(3029, 12), 1423 => to_unsigned(1711, 12), 1424 => to_unsigned(1628, 12), 1425 => to_unsigned(1919, 12), 1426 => to_unsigned(4033, 12), 1427 => to_unsigned(2857, 12), 1428 => to_unsigned(3878, 12), 1429 => to_unsigned(1420, 12), 1430 => to_unsigned(2255, 12), 1431 => to_unsigned(924, 12), 1432 => to_unsigned(1305, 12), 1433 => to_unsigned(2299, 12), 1434 => to_unsigned(1266, 12), 1435 => to_unsigned(53, 12), 1436 => to_unsigned(3542, 12), 1437 => to_unsigned(3775, 12), 1438 => to_unsigned(3419, 12), 1439 => to_unsigned(1101, 12), 1440 => to_unsigned(1697, 12), 1441 => to_unsigned(2510, 12), 1442 => to_unsigned(2421, 12), 1443 => to_unsigned(904, 12), 1444 => to_unsigned(3268, 12), 1445 => to_unsigned(2094, 12), 1446 => to_unsigned(3702, 12), 1447 => to_unsigned(853, 12), 1448 => to_unsigned(3757, 12), 1449 => to_unsigned(3548, 12), 1450 => to_unsigned(1814, 12), 1451 => to_unsigned(270, 12), 1452 => to_unsigned(2304, 12), 1453 => to_unsigned(434, 12), 1454 => to_unsigned(485, 12), 1455 => to_unsigned(2230, 12), 1456 => to_unsigned(1202, 12), 1457 => to_unsigned(2953, 12), 1458 => to_unsigned(1825, 12), 1459 => to_unsigned(3316, 12), 1460 => to_unsigned(1576, 12), 1461 => to_unsigned(680, 12), 1462 => to_unsigned(2803, 12), 1463 => to_unsigned(1927, 12), 1464 => to_unsigned(922, 12), 1465 => to_unsigned(3741, 12), 1466 => to_unsigned(1970, 12), 1467 => to_unsigned(185, 12), 1468 => to_unsigned(1553, 12), 1469 => to_unsigned(638, 12), 1470 => to_unsigned(2314, 12), 1471 => to_unsigned(2347, 12), 1472 => to_unsigned(3006, 12), 1473 => to_unsigned(225, 12), 1474 => to_unsigned(4033, 12), 1475 => to_unsigned(742, 12), 1476 => to_unsigned(3965, 12), 1477 => to_unsigned(787, 12), 1478 => to_unsigned(3293, 12), 1479 => to_unsigned(390, 12), 1480 => to_unsigned(3077, 12), 1481 => to_unsigned(3268, 12), 1482 => to_unsigned(1474, 12), 1483 => to_unsigned(3831, 12), 1484 => to_unsigned(3496, 12), 1485 => to_unsigned(2536, 12), 1486 => to_unsigned(4048, 12), 1487 => to_unsigned(839, 12), 1488 => to_unsigned(1960, 12), 1489 => to_unsigned(2840, 12), 1490 => to_unsigned(1239, 12), 1491 => to_unsigned(1716, 12), 1492 => to_unsigned(3450, 12), 1493 => to_unsigned(2710, 12), 1494 => to_unsigned(1577, 12), 1495 => to_unsigned(774, 12), 1496 => to_unsigned(2168, 12), 1497 => to_unsigned(3278, 12), 1498 => to_unsigned(563, 12), 1499 => to_unsigned(679, 12), 1500 => to_unsigned(3071, 12), 1501 => to_unsigned(536, 12), 1502 => to_unsigned(3103, 12), 1503 => to_unsigned(3732, 12), 1504 => to_unsigned(3730, 12), 1505 => to_unsigned(803, 12), 1506 => to_unsigned(3552, 12), 1507 => to_unsigned(2772, 12), 1508 => to_unsigned(1112, 12), 1509 => to_unsigned(2528, 12), 1510 => to_unsigned(1627, 12), 1511 => to_unsigned(3884, 12), 1512 => to_unsigned(4090, 12), 1513 => to_unsigned(868, 12), 1514 => to_unsigned(1490, 12), 1515 => to_unsigned(150, 12), 1516 => to_unsigned(1506, 12), 1517 => to_unsigned(927, 12), 1518 => to_unsigned(3762, 12), 1519 => to_unsigned(3858, 12), 1520 => to_unsigned(2556, 12), 1521 => to_unsigned(3150, 12), 1522 => to_unsigned(3591, 12), 1523 => to_unsigned(523, 12), 1524 => to_unsigned(1727, 12), 1525 => to_unsigned(1738, 12), 1526 => to_unsigned(3001, 12), 1527 => to_unsigned(1338, 12), 1528 => to_unsigned(2598, 12), 1529 => to_unsigned(1193, 12), 1530 => to_unsigned(3030, 12), 1531 => to_unsigned(4032, 12), 1532 => to_unsigned(1058, 12), 1533 => to_unsigned(209, 12), 1534 => to_unsigned(426, 12), 1535 => to_unsigned(4020, 12), 1536 => to_unsigned(3142, 12), 1537 => to_unsigned(3203, 12), 1538 => to_unsigned(2984, 12), 1539 => to_unsigned(3963, 12), 1540 => to_unsigned(91, 12), 1541 => to_unsigned(3020, 12), 1542 => to_unsigned(1703, 12), 1543 => to_unsigned(213, 12), 1544 => to_unsigned(793, 12), 1545 => to_unsigned(3840, 12), 1546 => to_unsigned(107, 12), 1547 => to_unsigned(4002, 12), 1548 => to_unsigned(1405, 12), 1549 => to_unsigned(3009, 12), 1550 => to_unsigned(1904, 12), 1551 => to_unsigned(2603, 12), 1552 => to_unsigned(2725, 12), 1553 => to_unsigned(4078, 12), 1554 => to_unsigned(107, 12), 1555 => to_unsigned(1497, 12), 1556 => to_unsigned(983, 12), 1557 => to_unsigned(3882, 12), 1558 => to_unsigned(3571, 12), 1559 => to_unsigned(708, 12), 1560 => to_unsigned(3764, 12), 1561 => to_unsigned(455, 12), 1562 => to_unsigned(1117, 12), 1563 => to_unsigned(2049, 12), 1564 => to_unsigned(23, 12), 1565 => to_unsigned(2263, 12), 1566 => to_unsigned(344, 12), 1567 => to_unsigned(2393, 12), 1568 => to_unsigned(2373, 12), 1569 => to_unsigned(1942, 12), 1570 => to_unsigned(4081, 12), 1571 => to_unsigned(1104, 12), 1572 => to_unsigned(2399, 12), 1573 => to_unsigned(3312, 12), 1574 => to_unsigned(1728, 12), 1575 => to_unsigned(498, 12), 1576 => to_unsigned(1987, 12), 1577 => to_unsigned(353, 12), 1578 => to_unsigned(3871, 12), 1579 => to_unsigned(1478, 12), 1580 => to_unsigned(1076, 12), 1581 => to_unsigned(3648, 12), 1582 => to_unsigned(1800, 12), 1583 => to_unsigned(2840, 12), 1584 => to_unsigned(1094, 12), 1585 => to_unsigned(1355, 12), 1586 => to_unsigned(4036, 12), 1587 => to_unsigned(3902, 12), 1588 => to_unsigned(1269, 12), 1589 => to_unsigned(1125, 12), 1590 => to_unsigned(3911, 12), 1591 => to_unsigned(1527, 12), 1592 => to_unsigned(1561, 12), 1593 => to_unsigned(2483, 12), 1594 => to_unsigned(2858, 12), 1595 => to_unsigned(2693, 12), 1596 => to_unsigned(4005, 12), 1597 => to_unsigned(900, 12), 1598 => to_unsigned(764, 12), 1599 => to_unsigned(1791, 12), 1600 => to_unsigned(3006, 12), 1601 => to_unsigned(1834, 12), 1602 => to_unsigned(3065, 12), 1603 => to_unsigned(3084, 12), 1604 => to_unsigned(2832, 12), 1605 => to_unsigned(3257, 12), 1606 => to_unsigned(3653, 12), 1607 => to_unsigned(13, 12), 1608 => to_unsigned(1803, 12), 1609 => to_unsigned(4054, 12), 1610 => to_unsigned(2410, 12), 1611 => to_unsigned(3367, 12), 1612 => to_unsigned(1280, 12), 1613 => to_unsigned(408, 12), 1614 => to_unsigned(2928, 12), 1615 => to_unsigned(2715, 12), 1616 => to_unsigned(887, 12), 1617 => to_unsigned(2718, 12), 1618 => to_unsigned(1240, 12), 1619 => to_unsigned(3036, 12), 1620 => to_unsigned(1432, 12), 1621 => to_unsigned(1791, 12), 1622 => to_unsigned(2942, 12), 1623 => to_unsigned(1118, 12), 1624 => to_unsigned(2681, 12), 1625 => to_unsigned(1972, 12), 1626 => to_unsigned(366, 12), 1627 => to_unsigned(2720, 12), 1628 => to_unsigned(4030, 12), 1629 => to_unsigned(3901, 12), 1630 => to_unsigned(1518, 12), 1631 => to_unsigned(995, 12), 1632 => to_unsigned(3158, 12), 1633 => to_unsigned(2863, 12), 1634 => to_unsigned(648, 12), 1635 => to_unsigned(3587, 12), 1636 => to_unsigned(612, 12), 1637 => to_unsigned(2740, 12), 1638 => to_unsigned(2254, 12), 1639 => to_unsigned(1852, 12), 1640 => to_unsigned(1764, 12), 1641 => to_unsigned(827, 12), 1642 => to_unsigned(1489, 12), 1643 => to_unsigned(955, 12), 1644 => to_unsigned(2003, 12), 1645 => to_unsigned(1368, 12), 1646 => to_unsigned(2136, 12), 1647 => to_unsigned(99, 12), 1648 => to_unsigned(1266, 12), 1649 => to_unsigned(3905, 12), 1650 => to_unsigned(204, 12), 1651 => to_unsigned(2388, 12), 1652 => to_unsigned(3079, 12), 1653 => to_unsigned(1110, 12), 1654 => to_unsigned(1836, 12), 1655 => to_unsigned(760, 12), 1656 => to_unsigned(207, 12), 1657 => to_unsigned(3104, 12), 1658 => to_unsigned(1057, 12), 1659 => to_unsigned(3405, 12), 1660 => to_unsigned(1665, 12), 1661 => to_unsigned(3587, 12), 1662 => to_unsigned(423, 12), 1663 => to_unsigned(248, 12), 1664 => to_unsigned(1470, 12), 1665 => to_unsigned(62, 12), 1666 => to_unsigned(3684, 12), 1667 => to_unsigned(3046, 12), 1668 => to_unsigned(2331, 12), 1669 => to_unsigned(954, 12), 1670 => to_unsigned(1634, 12), 1671 => to_unsigned(1389, 12), 1672 => to_unsigned(230, 12), 1673 => to_unsigned(3503, 12), 1674 => to_unsigned(1945, 12), 1675 => to_unsigned(1360, 12), 1676 => to_unsigned(3312, 12), 1677 => to_unsigned(3186, 12), 1678 => to_unsigned(1535, 12), 1679 => to_unsigned(3273, 12), 1680 => to_unsigned(2713, 12), 1681 => to_unsigned(3520, 12), 1682 => to_unsigned(1807, 12), 1683 => to_unsigned(3573, 12), 1684 => to_unsigned(1104, 12), 1685 => to_unsigned(3818, 12), 1686 => to_unsigned(2557, 12), 1687 => to_unsigned(1636, 12), 1688 => to_unsigned(7, 12), 1689 => to_unsigned(3479, 12), 1690 => to_unsigned(1265, 12), 1691 => to_unsigned(2344, 12), 1692 => to_unsigned(550, 12), 1693 => to_unsigned(3949, 12), 1694 => to_unsigned(2597, 12), 1695 => to_unsigned(1649, 12), 1696 => to_unsigned(1637, 12), 1697 => to_unsigned(1476, 12), 1698 => to_unsigned(3298, 12), 1699 => to_unsigned(3926, 12), 1700 => to_unsigned(4028, 12), 1701 => to_unsigned(3322, 12), 1702 => to_unsigned(3377, 12), 1703 => to_unsigned(542, 12), 1704 => to_unsigned(3835, 12), 1705 => to_unsigned(1761, 12), 1706 => to_unsigned(1499, 12), 1707 => to_unsigned(3399, 12), 1708 => to_unsigned(3789, 12), 1709 => to_unsigned(1753, 12), 1710 => to_unsigned(1445, 12), 1711 => to_unsigned(1951, 12), 1712 => to_unsigned(740, 12), 1713 => to_unsigned(1274, 12), 1714 => to_unsigned(2993, 12), 1715 => to_unsigned(1967, 12), 1716 => to_unsigned(2357, 12), 1717 => to_unsigned(615, 12), 1718 => to_unsigned(1672, 12), 1719 => to_unsigned(1810, 12), 1720 => to_unsigned(3028, 12), 1721 => to_unsigned(3097, 12), 1722 => to_unsigned(423, 12), 1723 => to_unsigned(2013, 12), 1724 => to_unsigned(258, 12), 1725 => to_unsigned(3560, 12), 1726 => to_unsigned(1714, 12), 1727 => to_unsigned(1233, 12), 1728 => to_unsigned(616, 12), 1729 => to_unsigned(3687, 12), 1730 => to_unsigned(609, 12), 1731 => to_unsigned(1027, 12), 1732 => to_unsigned(2074, 12), 1733 => to_unsigned(437, 12), 1734 => to_unsigned(3183, 12), 1735 => to_unsigned(2008, 12), 1736 => to_unsigned(2239, 12), 1737 => to_unsigned(1279, 12), 1738 => to_unsigned(4095, 12), 1739 => to_unsigned(369, 12), 1740 => to_unsigned(478, 12), 1741 => to_unsigned(627, 12), 1742 => to_unsigned(441, 12), 1743 => to_unsigned(1089, 12), 1744 => to_unsigned(3690, 12), 1745 => to_unsigned(850, 12), 1746 => to_unsigned(2375, 12), 1747 => to_unsigned(1707, 12), 1748 => to_unsigned(2629, 12), 1749 => to_unsigned(2874, 12), 1750 => to_unsigned(2472, 12), 1751 => to_unsigned(1637, 12), 1752 => to_unsigned(1683, 12), 1753 => to_unsigned(3106, 12), 1754 => to_unsigned(3285, 12), 1755 => to_unsigned(3044, 12), 1756 => to_unsigned(2136, 12), 1757 => to_unsigned(606, 12), 1758 => to_unsigned(3777, 12), 1759 => to_unsigned(640, 12), 1760 => to_unsigned(216, 12), 1761 => to_unsigned(365, 12), 1762 => to_unsigned(1839, 12), 1763 => to_unsigned(2936, 12), 1764 => to_unsigned(516, 12), 1765 => to_unsigned(2112, 12), 1766 => to_unsigned(1444, 12), 1767 => to_unsigned(3644, 12), 1768 => to_unsigned(3762, 12), 1769 => to_unsigned(3255, 12), 1770 => to_unsigned(468, 12), 1771 => to_unsigned(3908, 12), 1772 => to_unsigned(1797, 12), 1773 => to_unsigned(1725, 12), 1774 => to_unsigned(3534, 12), 1775 => to_unsigned(1046, 12), 1776 => to_unsigned(4047, 12), 1777 => to_unsigned(83, 12), 1778 => to_unsigned(844, 12), 1779 => to_unsigned(2365, 12), 1780 => to_unsigned(2215, 12), 1781 => to_unsigned(2848, 12), 1782 => to_unsigned(3769, 12), 1783 => to_unsigned(3102, 12), 1784 => to_unsigned(3412, 12), 1785 => to_unsigned(404, 12), 1786 => to_unsigned(2490, 12), 1787 => to_unsigned(581, 12), 1788 => to_unsigned(458, 12), 1789 => to_unsigned(344, 12), 1790 => to_unsigned(3275, 12), 1791 => to_unsigned(2965, 12), 1792 => to_unsigned(2300, 12), 1793 => to_unsigned(2374, 12), 1794 => to_unsigned(705, 12), 1795 => to_unsigned(3508, 12), 1796 => to_unsigned(525, 12), 1797 => to_unsigned(3919, 12), 1798 => to_unsigned(3695, 12), 1799 => to_unsigned(3883, 12), 1800 => to_unsigned(2005, 12), 1801 => to_unsigned(835, 12), 1802 => to_unsigned(2269, 12), 1803 => to_unsigned(1033, 12), 1804 => to_unsigned(566, 12), 1805 => to_unsigned(856, 12), 1806 => to_unsigned(2743, 12), 1807 => to_unsigned(2532, 12), 1808 => to_unsigned(3068, 12), 1809 => to_unsigned(1658, 12), 1810 => to_unsigned(823, 12), 1811 => to_unsigned(184, 12), 1812 => to_unsigned(3377, 12), 1813 => to_unsigned(2324, 12), 1814 => to_unsigned(3493, 12), 1815 => to_unsigned(4021, 12), 1816 => to_unsigned(3901, 12), 1817 => to_unsigned(4078, 12), 1818 => to_unsigned(1491, 12), 1819 => to_unsigned(3880, 12), 1820 => to_unsigned(1406, 12), 1821 => to_unsigned(579, 12), 1822 => to_unsigned(293, 12), 1823 => to_unsigned(1667, 12), 1824 => to_unsigned(3540, 12), 1825 => to_unsigned(2982, 12), 1826 => to_unsigned(734, 12), 1827 => to_unsigned(2849, 12), 1828 => to_unsigned(1113, 12), 1829 => to_unsigned(3241, 12), 1830 => to_unsigned(3820, 12), 1831 => to_unsigned(3575, 12), 1832 => to_unsigned(22, 12), 1833 => to_unsigned(1509, 12), 1834 => to_unsigned(2370, 12), 1835 => to_unsigned(569, 12), 1836 => to_unsigned(3739, 12), 1837 => to_unsigned(494, 12), 1838 => to_unsigned(243, 12), 1839 => to_unsigned(3301, 12), 1840 => to_unsigned(3130, 12), 1841 => to_unsigned(1144, 12), 1842 => to_unsigned(2204, 12), 1843 => to_unsigned(956, 12), 1844 => to_unsigned(2275, 12), 1845 => to_unsigned(2863, 12), 1846 => to_unsigned(1313, 12), 1847 => to_unsigned(2969, 12), 1848 => to_unsigned(3702, 12), 1849 => to_unsigned(2506, 12), 1850 => to_unsigned(231, 12), 1851 => to_unsigned(1480, 12), 1852 => to_unsigned(1489, 12), 1853 => to_unsigned(3289, 12), 1854 => to_unsigned(775, 12), 1855 => to_unsigned(4019, 12), 1856 => to_unsigned(1309, 12), 1857 => to_unsigned(2215, 12), 1858 => to_unsigned(425, 12), 1859 => to_unsigned(3860, 12), 1860 => to_unsigned(1313, 12), 1861 => to_unsigned(1649, 12), 1862 => to_unsigned(120, 12), 1863 => to_unsigned(1276, 12), 1864 => to_unsigned(1546, 12), 1865 => to_unsigned(3660, 12), 1866 => to_unsigned(1583, 12), 1867 => to_unsigned(1410, 12), 1868 => to_unsigned(736, 12), 1869 => to_unsigned(984, 12), 1870 => to_unsigned(309, 12), 1871 => to_unsigned(1349, 12), 1872 => to_unsigned(2451, 12), 1873 => to_unsigned(1408, 12), 1874 => to_unsigned(2449, 12), 1875 => to_unsigned(471, 12), 1876 => to_unsigned(3694, 12), 1877 => to_unsigned(3028, 12), 1878 => to_unsigned(58, 12), 1879 => to_unsigned(3044, 12), 1880 => to_unsigned(3748, 12), 1881 => to_unsigned(1420, 12), 1882 => to_unsigned(1708, 12), 1883 => to_unsigned(1764, 12), 1884 => to_unsigned(2895, 12), 1885 => to_unsigned(2469, 12), 1886 => to_unsigned(118, 12), 1887 => to_unsigned(408, 12), 1888 => to_unsigned(1709, 12), 1889 => to_unsigned(180, 12), 1890 => to_unsigned(3924, 12), 1891 => to_unsigned(890, 12), 1892 => to_unsigned(2748, 12), 1893 => to_unsigned(391, 12), 1894 => to_unsigned(1902, 12), 1895 => to_unsigned(1047, 12), 1896 => to_unsigned(2836, 12), 1897 => to_unsigned(2117, 12), 1898 => to_unsigned(2311, 12), 1899 => to_unsigned(804, 12), 1900 => to_unsigned(3183, 12), 1901 => to_unsigned(1673, 12), 1902 => to_unsigned(1221, 12), 1903 => to_unsigned(1305, 12), 1904 => to_unsigned(545, 12), 1905 => to_unsigned(1492, 12), 1906 => to_unsigned(2624, 12), 1907 => to_unsigned(2209, 12), 1908 => to_unsigned(3155, 12), 1909 => to_unsigned(3529, 12), 1910 => to_unsigned(258, 12), 1911 => to_unsigned(1552, 12), 1912 => to_unsigned(3198, 12), 1913 => to_unsigned(3159, 12), 1914 => to_unsigned(1853, 12), 1915 => to_unsigned(3898, 12), 1916 => to_unsigned(1650, 12), 1917 => to_unsigned(3097, 12), 1918 => to_unsigned(122, 12), 1919 => to_unsigned(2986, 12), 1920 => to_unsigned(720, 12), 1921 => to_unsigned(913, 12), 1922 => to_unsigned(40, 12), 1923 => to_unsigned(3388, 12), 1924 => to_unsigned(3409, 12), 1925 => to_unsigned(3578, 12), 1926 => to_unsigned(3325, 12), 1927 => to_unsigned(497, 12), 1928 => to_unsigned(1765, 12), 1929 => to_unsigned(425, 12), 1930 => to_unsigned(1446, 12), 1931 => to_unsigned(3276, 12), 1932 => to_unsigned(1222, 12), 1933 => to_unsigned(367, 12), 1934 => to_unsigned(1304, 12), 1935 => to_unsigned(3361, 12), 1936 => to_unsigned(2510, 12), 1937 => to_unsigned(197, 12), 1938 => to_unsigned(1033, 12), 1939 => to_unsigned(37, 12), 1940 => to_unsigned(1382, 12), 1941 => to_unsigned(1931, 12), 1942 => to_unsigned(921, 12), 1943 => to_unsigned(1808, 12), 1944 => to_unsigned(3155, 12), 1945 => to_unsigned(3901, 12), 1946 => to_unsigned(3450, 12), 1947 => to_unsigned(1943, 12), 1948 => to_unsigned(1458, 12), 1949 => to_unsigned(633, 12), 1950 => to_unsigned(1904, 12), 1951 => to_unsigned(3593, 12), 1952 => to_unsigned(1834, 12), 1953 => to_unsigned(2473, 12), 1954 => to_unsigned(1769, 12), 1955 => to_unsigned(3047, 12), 1956 => to_unsigned(2074, 12), 1957 => to_unsigned(3447, 12), 1958 => to_unsigned(630, 12), 1959 => to_unsigned(810, 12), 1960 => to_unsigned(2110, 12), 1961 => to_unsigned(1803, 12), 1962 => to_unsigned(3015, 12), 1963 => to_unsigned(3035, 12), 1964 => to_unsigned(1184, 12), 1965 => to_unsigned(637, 12), 1966 => to_unsigned(2846, 12), 1967 => to_unsigned(1878, 12), 1968 => to_unsigned(1309, 12), 1969 => to_unsigned(2080, 12), 1970 => to_unsigned(2498, 12), 1971 => to_unsigned(406, 12), 1972 => to_unsigned(1199, 12), 1973 => to_unsigned(2088, 12), 1974 => to_unsigned(2287, 12), 1975 => to_unsigned(408, 12), 1976 => to_unsigned(2422, 12), 1977 => to_unsigned(1011, 12), 1978 => to_unsigned(1678, 12), 1979 => to_unsigned(514, 12), 1980 => to_unsigned(1219, 12), 1981 => to_unsigned(2593, 12), 1982 => to_unsigned(2858, 12), 1983 => to_unsigned(1316, 12), 1984 => to_unsigned(128, 12), 1985 => to_unsigned(920, 12), 1986 => to_unsigned(1074, 12), 1987 => to_unsigned(2342, 12), 1988 => to_unsigned(3895, 12), 1989 => to_unsigned(268, 12), 1990 => to_unsigned(637, 12), 1991 => to_unsigned(1295, 12), 1992 => to_unsigned(26, 12), 1993 => to_unsigned(1943, 12), 1994 => to_unsigned(1720, 12), 1995 => to_unsigned(3037, 12), 1996 => to_unsigned(1808, 12), 1997 => to_unsigned(2386, 12), 1998 => to_unsigned(941, 12), 1999 => to_unsigned(3745, 12), 2000 => to_unsigned(246, 12), 2001 => to_unsigned(2435, 12), 2002 => to_unsigned(3642, 12), 2003 => to_unsigned(2918, 12), 2004 => to_unsigned(71, 12), 2005 => to_unsigned(2105, 12), 2006 => to_unsigned(1684, 12), 2007 => to_unsigned(2416, 12), 2008 => to_unsigned(1496, 12), 2009 => to_unsigned(2882, 12), 2010 => to_unsigned(3582, 12), 2011 => to_unsigned(2108, 12), 2012 => to_unsigned(522, 12), 2013 => to_unsigned(563, 12), 2014 => to_unsigned(3938, 12), 2015 => to_unsigned(3800, 12), 2016 => to_unsigned(1280, 12), 2017 => to_unsigned(2118, 12), 2018 => to_unsigned(2829, 12), 2019 => to_unsigned(2790, 12), 2020 => to_unsigned(1049, 12), 2021 => to_unsigned(1115, 12), 2022 => to_unsigned(2351, 12), 2023 => to_unsigned(2373, 12), 2024 => to_unsigned(3565, 12), 2025 => to_unsigned(2045, 12), 2026 => to_unsigned(1641, 12), 2027 => to_unsigned(2071, 12), 2028 => to_unsigned(4019, 12), 2029 => to_unsigned(2486, 12), 2030 => to_unsigned(3352, 12), 2031 => to_unsigned(1485, 12), 2032 => to_unsigned(1813, 12), 2033 => to_unsigned(1549, 12), 2034 => to_unsigned(3138, 12), 2035 => to_unsigned(3576, 12), 2036 => to_unsigned(2729, 12), 2037 => to_unsigned(2689, 12), 2038 => to_unsigned(2106, 12), 2039 => to_unsigned(4077, 12), 2040 => to_unsigned(2612, 12), 2041 => to_unsigned(3968, 12), 2042 => to_unsigned(3513, 12), 2043 => to_unsigned(1918, 12), 2044 => to_unsigned(2044, 12), 2045 => to_unsigned(2574, 12), 2046 => to_unsigned(3428, 12), 2047 => to_unsigned(3207, 12)),
            3 => (0 => to_unsigned(816, 12), 1 => to_unsigned(73, 12), 2 => to_unsigned(3180, 12), 3 => to_unsigned(2609, 12), 4 => to_unsigned(2564, 12), 5 => to_unsigned(2064, 12), 6 => to_unsigned(3216, 12), 7 => to_unsigned(3321, 12), 8 => to_unsigned(2879, 12), 9 => to_unsigned(3984, 12), 10 => to_unsigned(1475, 12), 11 => to_unsigned(2920, 12), 12 => to_unsigned(3254, 12), 13 => to_unsigned(3330, 12), 14 => to_unsigned(2592, 12), 15 => to_unsigned(1721, 12), 16 => to_unsigned(1350, 12), 17 => to_unsigned(981, 12), 18 => to_unsigned(668, 12), 19 => to_unsigned(790, 12), 20 => to_unsigned(3739, 12), 21 => to_unsigned(1913, 12), 22 => to_unsigned(2225, 12), 23 => to_unsigned(3966, 12), 24 => to_unsigned(3844, 12), 25 => to_unsigned(772, 12), 26 => to_unsigned(4063, 12), 27 => to_unsigned(1986, 12), 28 => to_unsigned(1241, 12), 29 => to_unsigned(1758, 12), 30 => to_unsigned(2379, 12), 31 => to_unsigned(2762, 12), 32 => to_unsigned(1218, 12), 33 => to_unsigned(1355, 12), 34 => to_unsigned(2636, 12), 35 => to_unsigned(3540, 12), 36 => to_unsigned(1673, 12), 37 => to_unsigned(2810, 12), 38 => to_unsigned(2083, 12), 39 => to_unsigned(3507, 12), 40 => to_unsigned(646, 12), 41 => to_unsigned(510, 12), 42 => to_unsigned(1567, 12), 43 => to_unsigned(1307, 12), 44 => to_unsigned(10, 12), 45 => to_unsigned(688, 12), 46 => to_unsigned(968, 12), 47 => to_unsigned(3289, 12), 48 => to_unsigned(1637, 12), 49 => to_unsigned(335, 12), 50 => to_unsigned(1562, 12), 51 => to_unsigned(837, 12), 52 => to_unsigned(2258, 12), 53 => to_unsigned(4032, 12), 54 => to_unsigned(4004, 12), 55 => to_unsigned(1056, 12), 56 => to_unsigned(1061, 12), 57 => to_unsigned(3666, 12), 58 => to_unsigned(2125, 12), 59 => to_unsigned(3795, 12), 60 => to_unsigned(2882, 12), 61 => to_unsigned(2287, 12), 62 => to_unsigned(3833, 12), 63 => to_unsigned(2216, 12), 64 => to_unsigned(1257, 12), 65 => to_unsigned(2176, 12), 66 => to_unsigned(166, 12), 67 => to_unsigned(320, 12), 68 => to_unsigned(905, 12), 69 => to_unsigned(3902, 12), 70 => to_unsigned(1969, 12), 71 => to_unsigned(1539, 12), 72 => to_unsigned(1157, 12), 73 => to_unsigned(2897, 12), 74 => to_unsigned(3836, 12), 75 => to_unsigned(1298, 12), 76 => to_unsigned(2861, 12), 77 => to_unsigned(715, 12), 78 => to_unsigned(576, 12), 79 => to_unsigned(3701, 12), 80 => to_unsigned(1318, 12), 81 => to_unsigned(108, 12), 82 => to_unsigned(1193, 12), 83 => to_unsigned(1553, 12), 84 => to_unsigned(1708, 12), 85 => to_unsigned(2706, 12), 86 => to_unsigned(3519, 12), 87 => to_unsigned(390, 12), 88 => to_unsigned(4047, 12), 89 => to_unsigned(822, 12), 90 => to_unsigned(2748, 12), 91 => to_unsigned(2471, 12), 92 => to_unsigned(384, 12), 93 => to_unsigned(1317, 12), 94 => to_unsigned(3620, 12), 95 => to_unsigned(135, 12), 96 => to_unsigned(3629, 12), 97 => to_unsigned(1535, 12), 98 => to_unsigned(3979, 12), 99 => to_unsigned(2692, 12), 100 => to_unsigned(1734, 12), 101 => to_unsigned(1574, 12), 102 => to_unsigned(892, 12), 103 => to_unsigned(808, 12), 104 => to_unsigned(3902, 12), 105 => to_unsigned(1862, 12), 106 => to_unsigned(3024, 12), 107 => to_unsigned(1698, 12), 108 => to_unsigned(848, 12), 109 => to_unsigned(1760, 12), 110 => to_unsigned(1016, 12), 111 => to_unsigned(1436, 12), 112 => to_unsigned(996, 12), 113 => to_unsigned(2976, 12), 114 => to_unsigned(3889, 12), 115 => to_unsigned(2032, 12), 116 => to_unsigned(264, 12), 117 => to_unsigned(3861, 12), 118 => to_unsigned(2098, 12), 119 => to_unsigned(1432, 12), 120 => to_unsigned(400, 12), 121 => to_unsigned(3157, 12), 122 => to_unsigned(266, 12), 123 => to_unsigned(160, 12), 124 => to_unsigned(2440, 12), 125 => to_unsigned(1211, 12), 126 => to_unsigned(2533, 12), 127 => to_unsigned(2502, 12), 128 => to_unsigned(1498, 12), 129 => to_unsigned(2154, 12), 130 => to_unsigned(1755, 12), 131 => to_unsigned(3834, 12), 132 => to_unsigned(1069, 12), 133 => to_unsigned(985, 12), 134 => to_unsigned(1684, 12), 135 => to_unsigned(468, 12), 136 => to_unsigned(2765, 12), 137 => to_unsigned(2210, 12), 138 => to_unsigned(3332, 12), 139 => to_unsigned(1584, 12), 140 => to_unsigned(1998, 12), 141 => to_unsigned(1560, 12), 142 => to_unsigned(705, 12), 143 => to_unsigned(615, 12), 144 => to_unsigned(2859, 12), 145 => to_unsigned(2253, 12), 146 => to_unsigned(228, 12), 147 => to_unsigned(1505, 12), 148 => to_unsigned(1228, 12), 149 => to_unsigned(1552, 12), 150 => to_unsigned(1081, 12), 151 => to_unsigned(3589, 12), 152 => to_unsigned(3041, 12), 153 => to_unsigned(1403, 12), 154 => to_unsigned(3807, 12), 155 => to_unsigned(3080, 12), 156 => to_unsigned(3105, 12), 157 => to_unsigned(2358, 12), 158 => to_unsigned(1344, 12), 159 => to_unsigned(2464, 12), 160 => to_unsigned(2527, 12), 161 => to_unsigned(3842, 12), 162 => to_unsigned(490, 12), 163 => to_unsigned(2203, 12), 164 => to_unsigned(1744, 12), 165 => to_unsigned(87, 12), 166 => to_unsigned(3906, 12), 167 => to_unsigned(967, 12), 168 => to_unsigned(3813, 12), 169 => to_unsigned(45, 12), 170 => to_unsigned(1684, 12), 171 => to_unsigned(1728, 12), 172 => to_unsigned(647, 12), 173 => to_unsigned(473, 12), 174 => to_unsigned(792, 12), 175 => to_unsigned(193, 12), 176 => to_unsigned(611, 12), 177 => to_unsigned(1342, 12), 178 => to_unsigned(2142, 12), 179 => to_unsigned(2466, 12), 180 => to_unsigned(2268, 12), 181 => to_unsigned(2274, 12), 182 => to_unsigned(3989, 12), 183 => to_unsigned(2391, 12), 184 => to_unsigned(913, 12), 185 => to_unsigned(1349, 12), 186 => to_unsigned(3967, 12), 187 => to_unsigned(2819, 12), 188 => to_unsigned(345, 12), 189 => to_unsigned(2197, 12), 190 => to_unsigned(699, 12), 191 => to_unsigned(646, 12), 192 => to_unsigned(1725, 12), 193 => to_unsigned(723, 12), 194 => to_unsigned(3094, 12), 195 => to_unsigned(1559, 12), 196 => to_unsigned(1109, 12), 197 => to_unsigned(1100, 12), 198 => to_unsigned(2710, 12), 199 => to_unsigned(1084, 12), 200 => to_unsigned(906, 12), 201 => to_unsigned(2766, 12), 202 => to_unsigned(3052, 12), 203 => to_unsigned(2233, 12), 204 => to_unsigned(3113, 12), 205 => to_unsigned(1605, 12), 206 => to_unsigned(1703, 12), 207 => to_unsigned(3829, 12), 208 => to_unsigned(883, 12), 209 => to_unsigned(1482, 12), 210 => to_unsigned(2493, 12), 211 => to_unsigned(2394, 12), 212 => to_unsigned(410, 12), 213 => to_unsigned(3795, 12), 214 => to_unsigned(3246, 12), 215 => to_unsigned(628, 12), 216 => to_unsigned(3216, 12), 217 => to_unsigned(3713, 12), 218 => to_unsigned(211, 12), 219 => to_unsigned(2382, 12), 220 => to_unsigned(3593, 12), 221 => to_unsigned(2879, 12), 222 => to_unsigned(1516, 12), 223 => to_unsigned(2367, 12), 224 => to_unsigned(3516, 12), 225 => to_unsigned(3235, 12), 226 => to_unsigned(3427, 12), 227 => to_unsigned(2184, 12), 228 => to_unsigned(1754, 12), 229 => to_unsigned(3640, 12), 230 => to_unsigned(2419, 12), 231 => to_unsigned(2408, 12), 232 => to_unsigned(173, 12), 233 => to_unsigned(2893, 12), 234 => to_unsigned(3261, 12), 235 => to_unsigned(2777, 12), 236 => to_unsigned(3372, 12), 237 => to_unsigned(2996, 12), 238 => to_unsigned(2574, 12), 239 => to_unsigned(3568, 12), 240 => to_unsigned(1165, 12), 241 => to_unsigned(2618, 12), 242 => to_unsigned(902, 12), 243 => to_unsigned(363, 12), 244 => to_unsigned(2300, 12), 245 => to_unsigned(1608, 12), 246 => to_unsigned(742, 12), 247 => to_unsigned(1075, 12), 248 => to_unsigned(2830, 12), 249 => to_unsigned(622, 12), 250 => to_unsigned(2844, 12), 251 => to_unsigned(157, 12), 252 => to_unsigned(3295, 12), 253 => to_unsigned(94, 12), 254 => to_unsigned(1288, 12), 255 => to_unsigned(619, 12), 256 => to_unsigned(2498, 12), 257 => to_unsigned(2104, 12), 258 => to_unsigned(1359, 12), 259 => to_unsigned(440, 12), 260 => to_unsigned(1976, 12), 261 => to_unsigned(3036, 12), 262 => to_unsigned(3938, 12), 263 => to_unsigned(805, 12), 264 => to_unsigned(1706, 12), 265 => to_unsigned(3174, 12), 266 => to_unsigned(1381, 12), 267 => to_unsigned(2264, 12), 268 => to_unsigned(261, 12), 269 => to_unsigned(1934, 12), 270 => to_unsigned(1720, 12), 271 => to_unsigned(1250, 12), 272 => to_unsigned(1419, 12), 273 => to_unsigned(1936, 12), 274 => to_unsigned(1695, 12), 275 => to_unsigned(1266, 12), 276 => to_unsigned(588, 12), 277 => to_unsigned(3258, 12), 278 => to_unsigned(3003, 12), 279 => to_unsigned(2496, 12), 280 => to_unsigned(1981, 12), 281 => to_unsigned(1890, 12), 282 => to_unsigned(4089, 12), 283 => to_unsigned(576, 12), 284 => to_unsigned(632, 12), 285 => to_unsigned(57, 12), 286 => to_unsigned(1680, 12), 287 => to_unsigned(1919, 12), 288 => to_unsigned(644, 12), 289 => to_unsigned(3428, 12), 290 => to_unsigned(1539, 12), 291 => to_unsigned(3461, 12), 292 => to_unsigned(734, 12), 293 => to_unsigned(3323, 12), 294 => to_unsigned(3122, 12), 295 => to_unsigned(1407, 12), 296 => to_unsigned(3242, 12), 297 => to_unsigned(2772, 12), 298 => to_unsigned(3504, 12), 299 => to_unsigned(813, 12), 300 => to_unsigned(271, 12), 301 => to_unsigned(2277, 12), 302 => to_unsigned(2281, 12), 303 => to_unsigned(1141, 12), 304 => to_unsigned(1756, 12), 305 => to_unsigned(1627, 12), 306 => to_unsigned(183, 12), 307 => to_unsigned(1211, 12), 308 => to_unsigned(3579, 12), 309 => to_unsigned(3565, 12), 310 => to_unsigned(3255, 12), 311 => to_unsigned(2941, 12), 312 => to_unsigned(673, 12), 313 => to_unsigned(2315, 12), 314 => to_unsigned(2687, 12), 315 => to_unsigned(4059, 12), 316 => to_unsigned(2850, 12), 317 => to_unsigned(3544, 12), 318 => to_unsigned(1293, 12), 319 => to_unsigned(2439, 12), 320 => to_unsigned(3480, 12), 321 => to_unsigned(2753, 12), 322 => to_unsigned(1123, 12), 323 => to_unsigned(3666, 12), 324 => to_unsigned(2414, 12), 325 => to_unsigned(2344, 12), 326 => to_unsigned(1719, 12), 327 => to_unsigned(2625, 12), 328 => to_unsigned(1258, 12), 329 => to_unsigned(1307, 12), 330 => to_unsigned(2959, 12), 331 => to_unsigned(3215, 12), 332 => to_unsigned(2345, 12), 333 => to_unsigned(4045, 12), 334 => to_unsigned(1542, 12), 335 => to_unsigned(3710, 12), 336 => to_unsigned(3322, 12), 337 => to_unsigned(3296, 12), 338 => to_unsigned(1500, 12), 339 => to_unsigned(3896, 12), 340 => to_unsigned(180, 12), 341 => to_unsigned(3718, 12), 342 => to_unsigned(1358, 12), 343 => to_unsigned(1439, 12), 344 => to_unsigned(2438, 12), 345 => to_unsigned(545, 12), 346 => to_unsigned(383, 12), 347 => to_unsigned(3258, 12), 348 => to_unsigned(1786, 12), 349 => to_unsigned(1918, 12), 350 => to_unsigned(2094, 12), 351 => to_unsigned(639, 12), 352 => to_unsigned(538, 12), 353 => to_unsigned(1075, 12), 354 => to_unsigned(1184, 12), 355 => to_unsigned(3772, 12), 356 => to_unsigned(1787, 12), 357 => to_unsigned(1838, 12), 358 => to_unsigned(3167, 12), 359 => to_unsigned(647, 12), 360 => to_unsigned(689, 12), 361 => to_unsigned(807, 12), 362 => to_unsigned(3265, 12), 363 => to_unsigned(1285, 12), 364 => to_unsigned(1637, 12), 365 => to_unsigned(2715, 12), 366 => to_unsigned(1958, 12), 367 => to_unsigned(1581, 12), 368 => to_unsigned(663, 12), 369 => to_unsigned(268, 12), 370 => to_unsigned(649, 12), 371 => to_unsigned(2205, 12), 372 => to_unsigned(2205, 12), 373 => to_unsigned(2061, 12), 374 => to_unsigned(599, 12), 375 => to_unsigned(1816, 12), 376 => to_unsigned(649, 12), 377 => to_unsigned(3140, 12), 378 => to_unsigned(1445, 12), 379 => to_unsigned(1464, 12), 380 => to_unsigned(1739, 12), 381 => to_unsigned(2390, 12), 382 => to_unsigned(2236, 12), 383 => to_unsigned(3736, 12), 384 => to_unsigned(1637, 12), 385 => to_unsigned(104, 12), 386 => to_unsigned(488, 12), 387 => to_unsigned(1204, 12), 388 => to_unsigned(565, 12), 389 => to_unsigned(3938, 12), 390 => to_unsigned(942, 12), 391 => to_unsigned(2721, 12), 392 => to_unsigned(3066, 12), 393 => to_unsigned(2701, 12), 394 => to_unsigned(481, 12), 395 => to_unsigned(455, 12), 396 => to_unsigned(1548, 12), 397 => to_unsigned(1225, 12), 398 => to_unsigned(2478, 12), 399 => to_unsigned(285, 12), 400 => to_unsigned(2316, 12), 401 => to_unsigned(1719, 12), 402 => to_unsigned(1072, 12), 403 => to_unsigned(246, 12), 404 => to_unsigned(3875, 12), 405 => to_unsigned(2082, 12), 406 => to_unsigned(3130, 12), 407 => to_unsigned(3772, 12), 408 => to_unsigned(3713, 12), 409 => to_unsigned(2705, 12), 410 => to_unsigned(171, 12), 411 => to_unsigned(1776, 12), 412 => to_unsigned(2487, 12), 413 => to_unsigned(2057, 12), 414 => to_unsigned(2487, 12), 415 => to_unsigned(2809, 12), 416 => to_unsigned(1021, 12), 417 => to_unsigned(1680, 12), 418 => to_unsigned(835, 12), 419 => to_unsigned(2729, 12), 420 => to_unsigned(2518, 12), 421 => to_unsigned(815, 12), 422 => to_unsigned(724, 12), 423 => to_unsigned(2136, 12), 424 => to_unsigned(3297, 12), 425 => to_unsigned(507, 12), 426 => to_unsigned(1850, 12), 427 => to_unsigned(4052, 12), 428 => to_unsigned(3285, 12), 429 => to_unsigned(804, 12), 430 => to_unsigned(3820, 12), 431 => to_unsigned(3340, 12), 432 => to_unsigned(26, 12), 433 => to_unsigned(3074, 12), 434 => to_unsigned(1018, 12), 435 => to_unsigned(3834, 12), 436 => to_unsigned(790, 12), 437 => to_unsigned(1582, 12), 438 => to_unsigned(1875, 12), 439 => to_unsigned(2297, 12), 440 => to_unsigned(2066, 12), 441 => to_unsigned(3106, 12), 442 => to_unsigned(1119, 12), 443 => to_unsigned(3267, 12), 444 => to_unsigned(0, 12), 445 => to_unsigned(1691, 12), 446 => to_unsigned(2096, 12), 447 => to_unsigned(3566, 12), 448 => to_unsigned(726, 12), 449 => to_unsigned(500, 12), 450 => to_unsigned(3971, 12), 451 => to_unsigned(3836, 12), 452 => to_unsigned(2016, 12), 453 => to_unsigned(11, 12), 454 => to_unsigned(2672, 12), 455 => to_unsigned(1752, 12), 456 => to_unsigned(2204, 12), 457 => to_unsigned(2344, 12), 458 => to_unsigned(1225, 12), 459 => to_unsigned(2818, 12), 460 => to_unsigned(1486, 12), 461 => to_unsigned(2619, 12), 462 => to_unsigned(3060, 12), 463 => to_unsigned(778, 12), 464 => to_unsigned(3460, 12), 465 => to_unsigned(1737, 12), 466 => to_unsigned(2413, 12), 467 => to_unsigned(1151, 12), 468 => to_unsigned(1114, 12), 469 => to_unsigned(3691, 12), 470 => to_unsigned(253, 12), 471 => to_unsigned(264, 12), 472 => to_unsigned(3365, 12), 473 => to_unsigned(4072, 12), 474 => to_unsigned(2274, 12), 475 => to_unsigned(3052, 12), 476 => to_unsigned(2806, 12), 477 => to_unsigned(3174, 12), 478 => to_unsigned(1883, 12), 479 => to_unsigned(2800, 12), 480 => to_unsigned(442, 12), 481 => to_unsigned(3002, 12), 482 => to_unsigned(4017, 12), 483 => to_unsigned(245, 12), 484 => to_unsigned(2323, 12), 485 => to_unsigned(3875, 12), 486 => to_unsigned(2468, 12), 487 => to_unsigned(636, 12), 488 => to_unsigned(1354, 12), 489 => to_unsigned(1329, 12), 490 => to_unsigned(658, 12), 491 => to_unsigned(3332, 12), 492 => to_unsigned(1496, 12), 493 => to_unsigned(975, 12), 494 => to_unsigned(817, 12), 495 => to_unsigned(990, 12), 496 => to_unsigned(2317, 12), 497 => to_unsigned(435, 12), 498 => to_unsigned(1424, 12), 499 => to_unsigned(2487, 12), 500 => to_unsigned(104, 12), 501 => to_unsigned(1005, 12), 502 => to_unsigned(3787, 12), 503 => to_unsigned(3133, 12), 504 => to_unsigned(354, 12), 505 => to_unsigned(1297, 12), 506 => to_unsigned(2758, 12), 507 => to_unsigned(3608, 12), 508 => to_unsigned(3677, 12), 509 => to_unsigned(3293, 12), 510 => to_unsigned(2626, 12), 511 => to_unsigned(203, 12), 512 => to_unsigned(4090, 12), 513 => to_unsigned(3118, 12), 514 => to_unsigned(168, 12), 515 => to_unsigned(1745, 12), 516 => to_unsigned(1191, 12), 517 => to_unsigned(2559, 12), 518 => to_unsigned(777, 12), 519 => to_unsigned(363, 12), 520 => to_unsigned(3354, 12), 521 => to_unsigned(788, 12), 522 => to_unsigned(953, 12), 523 => to_unsigned(3012, 12), 524 => to_unsigned(2666, 12), 525 => to_unsigned(1346, 12), 526 => to_unsigned(1076, 12), 527 => to_unsigned(2855, 12), 528 => to_unsigned(851, 12), 529 => to_unsigned(1471, 12), 530 => to_unsigned(1396, 12), 531 => to_unsigned(1671, 12), 532 => to_unsigned(2591, 12), 533 => to_unsigned(3168, 12), 534 => to_unsigned(2244, 12), 535 => to_unsigned(1012, 12), 536 => to_unsigned(2203, 12), 537 => to_unsigned(1176, 12), 538 => to_unsigned(1002, 12), 539 => to_unsigned(2871, 12), 540 => to_unsigned(648, 12), 541 => to_unsigned(556, 12), 542 => to_unsigned(2869, 12), 543 => to_unsigned(1754, 12), 544 => to_unsigned(3622, 12), 545 => to_unsigned(3227, 12), 546 => to_unsigned(2274, 12), 547 => to_unsigned(1067, 12), 548 => to_unsigned(1996, 12), 549 => to_unsigned(3823, 12), 550 => to_unsigned(1544, 12), 551 => to_unsigned(680, 12), 552 => to_unsigned(2680, 12), 553 => to_unsigned(3565, 12), 554 => to_unsigned(288, 12), 555 => to_unsigned(1472, 12), 556 => to_unsigned(4079, 12), 557 => to_unsigned(721, 12), 558 => to_unsigned(1740, 12), 559 => to_unsigned(1552, 12), 560 => to_unsigned(117, 12), 561 => to_unsigned(3832, 12), 562 => to_unsigned(331, 12), 563 => to_unsigned(2639, 12), 564 => to_unsigned(1244, 12), 565 => to_unsigned(1587, 12), 566 => to_unsigned(1472, 12), 567 => to_unsigned(1902, 12), 568 => to_unsigned(732, 12), 569 => to_unsigned(932, 12), 570 => to_unsigned(1084, 12), 571 => to_unsigned(3602, 12), 572 => to_unsigned(721, 12), 573 => to_unsigned(1177, 12), 574 => to_unsigned(2600, 12), 575 => to_unsigned(921, 12), 576 => to_unsigned(1796, 12), 577 => to_unsigned(1930, 12), 578 => to_unsigned(2145, 12), 579 => to_unsigned(3158, 12), 580 => to_unsigned(225, 12), 581 => to_unsigned(2414, 12), 582 => to_unsigned(3282, 12), 583 => to_unsigned(1699, 12), 584 => to_unsigned(1776, 12), 585 => to_unsigned(1620, 12), 586 => to_unsigned(901, 12), 587 => to_unsigned(314, 12), 588 => to_unsigned(3683, 12), 589 => to_unsigned(3503, 12), 590 => to_unsigned(461, 12), 591 => to_unsigned(2536, 12), 592 => to_unsigned(3175, 12), 593 => to_unsigned(2462, 12), 594 => to_unsigned(2443, 12), 595 => to_unsigned(3080, 12), 596 => to_unsigned(2169, 12), 597 => to_unsigned(1050, 12), 598 => to_unsigned(3176, 12), 599 => to_unsigned(95, 12), 600 => to_unsigned(2010, 12), 601 => to_unsigned(562, 12), 602 => to_unsigned(1253, 12), 603 => to_unsigned(3091, 12), 604 => to_unsigned(2487, 12), 605 => to_unsigned(1276, 12), 606 => to_unsigned(799, 12), 607 => to_unsigned(1990, 12), 608 => to_unsigned(947, 12), 609 => to_unsigned(293, 12), 610 => to_unsigned(2699, 12), 611 => to_unsigned(3407, 12), 612 => to_unsigned(940, 12), 613 => to_unsigned(3381, 12), 614 => to_unsigned(132, 12), 615 => to_unsigned(1507, 12), 616 => to_unsigned(242, 12), 617 => to_unsigned(1937, 12), 618 => to_unsigned(492, 12), 619 => to_unsigned(537, 12), 620 => to_unsigned(2998, 12), 621 => to_unsigned(3450, 12), 622 => to_unsigned(3660, 12), 623 => to_unsigned(1792, 12), 624 => to_unsigned(3936, 12), 625 => to_unsigned(1990, 12), 626 => to_unsigned(1763, 12), 627 => to_unsigned(3497, 12), 628 => to_unsigned(2408, 12), 629 => to_unsigned(1107, 12), 630 => to_unsigned(3707, 12), 631 => to_unsigned(2147, 12), 632 => to_unsigned(3421, 12), 633 => to_unsigned(2538, 12), 634 => to_unsigned(727, 12), 635 => to_unsigned(793, 12), 636 => to_unsigned(1236, 12), 637 => to_unsigned(2939, 12), 638 => to_unsigned(428, 12), 639 => to_unsigned(3400, 12), 640 => to_unsigned(3110, 12), 641 => to_unsigned(1494, 12), 642 => to_unsigned(3303, 12), 643 => to_unsigned(306, 12), 644 => to_unsigned(3061, 12), 645 => to_unsigned(655, 12), 646 => to_unsigned(1535, 12), 647 => to_unsigned(3972, 12), 648 => to_unsigned(3787, 12), 649 => to_unsigned(3354, 12), 650 => to_unsigned(1099, 12), 651 => to_unsigned(1818, 12), 652 => to_unsigned(1996, 12), 653 => to_unsigned(2844, 12), 654 => to_unsigned(3968, 12), 655 => to_unsigned(325, 12), 656 => to_unsigned(2105, 12), 657 => to_unsigned(2534, 12), 658 => to_unsigned(525, 12), 659 => to_unsigned(3862, 12), 660 => to_unsigned(763, 12), 661 => to_unsigned(1275, 12), 662 => to_unsigned(4056, 12), 663 => to_unsigned(3389, 12), 664 => to_unsigned(602, 12), 665 => to_unsigned(1598, 12), 666 => to_unsigned(3717, 12), 667 => to_unsigned(2898, 12), 668 => to_unsigned(3884, 12), 669 => to_unsigned(3438, 12), 670 => to_unsigned(2268, 12), 671 => to_unsigned(1603, 12), 672 => to_unsigned(3095, 12), 673 => to_unsigned(2953, 12), 674 => to_unsigned(1459, 12), 675 => to_unsigned(1541, 12), 676 => to_unsigned(218, 12), 677 => to_unsigned(1569, 12), 678 => to_unsigned(2177, 12), 679 => to_unsigned(3135, 12), 680 => to_unsigned(1504, 12), 681 => to_unsigned(2132, 12), 682 => to_unsigned(3577, 12), 683 => to_unsigned(2749, 12), 684 => to_unsigned(1519, 12), 685 => to_unsigned(3419, 12), 686 => to_unsigned(2794, 12), 687 => to_unsigned(204, 12), 688 => to_unsigned(1311, 12), 689 => to_unsigned(3309, 12), 690 => to_unsigned(3547, 12), 691 => to_unsigned(4026, 12), 692 => to_unsigned(2435, 12), 693 => to_unsigned(2291, 12), 694 => to_unsigned(1620, 12), 695 => to_unsigned(1418, 12), 696 => to_unsigned(1203, 12), 697 => to_unsigned(2121, 12), 698 => to_unsigned(1989, 12), 699 => to_unsigned(141, 12), 700 => to_unsigned(3388, 12), 701 => to_unsigned(3688, 12), 702 => to_unsigned(2897, 12), 703 => to_unsigned(1466, 12), 704 => to_unsigned(301, 12), 705 => to_unsigned(2201, 12), 706 => to_unsigned(2947, 12), 707 => to_unsigned(2496, 12), 708 => to_unsigned(3830, 12), 709 => to_unsigned(2766, 12), 710 => to_unsigned(1268, 12), 711 => to_unsigned(3854, 12), 712 => to_unsigned(2263, 12), 713 => to_unsigned(3014, 12), 714 => to_unsigned(271, 12), 715 => to_unsigned(1541, 12), 716 => to_unsigned(822, 12), 717 => to_unsigned(3584, 12), 718 => to_unsigned(1767, 12), 719 => to_unsigned(711, 12), 720 => to_unsigned(1981, 12), 721 => to_unsigned(3409, 12), 722 => to_unsigned(3872, 12), 723 => to_unsigned(3130, 12), 724 => to_unsigned(2589, 12), 725 => to_unsigned(3999, 12), 726 => to_unsigned(463, 12), 727 => to_unsigned(1739, 12), 728 => to_unsigned(3051, 12), 729 => to_unsigned(3487, 12), 730 => to_unsigned(3346, 12), 731 => to_unsigned(3179, 12), 732 => to_unsigned(102, 12), 733 => to_unsigned(3542, 12), 734 => to_unsigned(3399, 12), 735 => to_unsigned(1780, 12), 736 => to_unsigned(3555, 12), 737 => to_unsigned(3774, 12), 738 => to_unsigned(3603, 12), 739 => to_unsigned(3397, 12), 740 => to_unsigned(2737, 12), 741 => to_unsigned(2240, 12), 742 => to_unsigned(491, 12), 743 => to_unsigned(3457, 12), 744 => to_unsigned(3890, 12), 745 => to_unsigned(3765, 12), 746 => to_unsigned(3644, 12), 747 => to_unsigned(2618, 12), 748 => to_unsigned(4046, 12), 749 => to_unsigned(3956, 12), 750 => to_unsigned(3769, 12), 751 => to_unsigned(1682, 12), 752 => to_unsigned(3241, 12), 753 => to_unsigned(1798, 12), 754 => to_unsigned(2276, 12), 755 => to_unsigned(171, 12), 756 => to_unsigned(1777, 12), 757 => to_unsigned(928, 12), 758 => to_unsigned(3915, 12), 759 => to_unsigned(2263, 12), 760 => to_unsigned(2683, 12), 761 => to_unsigned(1816, 12), 762 => to_unsigned(1074, 12), 763 => to_unsigned(1416, 12), 764 => to_unsigned(117, 12), 765 => to_unsigned(1619, 12), 766 => to_unsigned(258, 12), 767 => to_unsigned(3570, 12), 768 => to_unsigned(28, 12), 769 => to_unsigned(3110, 12), 770 => to_unsigned(1272, 12), 771 => to_unsigned(3502, 12), 772 => to_unsigned(2859, 12), 773 => to_unsigned(3937, 12), 774 => to_unsigned(3956, 12), 775 => to_unsigned(2061, 12), 776 => to_unsigned(3373, 12), 777 => to_unsigned(2593, 12), 778 => to_unsigned(1802, 12), 779 => to_unsigned(1907, 12), 780 => to_unsigned(2903, 12), 781 => to_unsigned(3965, 12), 782 => to_unsigned(2893, 12), 783 => to_unsigned(1395, 12), 784 => to_unsigned(494, 12), 785 => to_unsigned(1822, 12), 786 => to_unsigned(64, 12), 787 => to_unsigned(2411, 12), 788 => to_unsigned(1223, 12), 789 => to_unsigned(2371, 12), 790 => to_unsigned(638, 12), 791 => to_unsigned(1390, 12), 792 => to_unsigned(1152, 12), 793 => to_unsigned(3935, 12), 794 => to_unsigned(2440, 12), 795 => to_unsigned(3395, 12), 796 => to_unsigned(2571, 12), 797 => to_unsigned(1431, 12), 798 => to_unsigned(1556, 12), 799 => to_unsigned(769, 12), 800 => to_unsigned(710, 12), 801 => to_unsigned(2286, 12), 802 => to_unsigned(3068, 12), 803 => to_unsigned(324, 12), 804 => to_unsigned(1194, 12), 805 => to_unsigned(355, 12), 806 => to_unsigned(1148, 12), 807 => to_unsigned(1263, 12), 808 => to_unsigned(3350, 12), 809 => to_unsigned(2206, 12), 810 => to_unsigned(2086, 12), 811 => to_unsigned(331, 12), 812 => to_unsigned(3892, 12), 813 => to_unsigned(866, 12), 814 => to_unsigned(1527, 12), 815 => to_unsigned(1731, 12), 816 => to_unsigned(1393, 12), 817 => to_unsigned(490, 12), 818 => to_unsigned(3264, 12), 819 => to_unsigned(1030, 12), 820 => to_unsigned(1569, 12), 821 => to_unsigned(2046, 12), 822 => to_unsigned(285, 12), 823 => to_unsigned(2389, 12), 824 => to_unsigned(3086, 12), 825 => to_unsigned(1844, 12), 826 => to_unsigned(598, 12), 827 => to_unsigned(2139, 12), 828 => to_unsigned(1219, 12), 829 => to_unsigned(1905, 12), 830 => to_unsigned(2047, 12), 831 => to_unsigned(2910, 12), 832 => to_unsigned(2151, 12), 833 => to_unsigned(430, 12), 834 => to_unsigned(1367, 12), 835 => to_unsigned(24, 12), 836 => to_unsigned(3307, 12), 837 => to_unsigned(397, 12), 838 => to_unsigned(2464, 12), 839 => to_unsigned(2080, 12), 840 => to_unsigned(1266, 12), 841 => to_unsigned(3446, 12), 842 => to_unsigned(1521, 12), 843 => to_unsigned(3865, 12), 844 => to_unsigned(2889, 12), 845 => to_unsigned(1381, 12), 846 => to_unsigned(3436, 12), 847 => to_unsigned(2705, 12), 848 => to_unsigned(3735, 12), 849 => to_unsigned(2339, 12), 850 => to_unsigned(3067, 12), 851 => to_unsigned(2425, 12), 852 => to_unsigned(3875, 12), 853 => to_unsigned(3746, 12), 854 => to_unsigned(2132, 12), 855 => to_unsigned(453, 12), 856 => to_unsigned(2836, 12), 857 => to_unsigned(3846, 12), 858 => to_unsigned(904, 12), 859 => to_unsigned(3840, 12), 860 => to_unsigned(829, 12), 861 => to_unsigned(748, 12), 862 => to_unsigned(3673, 12), 863 => to_unsigned(3430, 12), 864 => to_unsigned(71, 12), 865 => to_unsigned(3529, 12), 866 => to_unsigned(2426, 12), 867 => to_unsigned(2822, 12), 868 => to_unsigned(2269, 12), 869 => to_unsigned(3525, 12), 870 => to_unsigned(932, 12), 871 => to_unsigned(669, 12), 872 => to_unsigned(103, 12), 873 => to_unsigned(3603, 12), 874 => to_unsigned(3631, 12), 875 => to_unsigned(1430, 12), 876 => to_unsigned(2115, 12), 877 => to_unsigned(2183, 12), 878 => to_unsigned(3640, 12), 879 => to_unsigned(93, 12), 880 => to_unsigned(212, 12), 881 => to_unsigned(3912, 12), 882 => to_unsigned(2706, 12), 883 => to_unsigned(1430, 12), 884 => to_unsigned(2198, 12), 885 => to_unsigned(1493, 12), 886 => to_unsigned(1582, 12), 887 => to_unsigned(2343, 12), 888 => to_unsigned(2616, 12), 889 => to_unsigned(2210, 12), 890 => to_unsigned(1596, 12), 891 => to_unsigned(3682, 12), 892 => to_unsigned(1023, 12), 893 => to_unsigned(1488, 12), 894 => to_unsigned(909, 12), 895 => to_unsigned(540, 12), 896 => to_unsigned(3320, 12), 897 => to_unsigned(2619, 12), 898 => to_unsigned(13, 12), 899 => to_unsigned(1441, 12), 900 => to_unsigned(1658, 12), 901 => to_unsigned(2714, 12), 902 => to_unsigned(2125, 12), 903 => to_unsigned(3001, 12), 904 => to_unsigned(1149, 12), 905 => to_unsigned(3658, 12), 906 => to_unsigned(3578, 12), 907 => to_unsigned(2647, 12), 908 => to_unsigned(2261, 12), 909 => to_unsigned(1627, 12), 910 => to_unsigned(3565, 12), 911 => to_unsigned(567, 12), 912 => to_unsigned(2556, 12), 913 => to_unsigned(2133, 12), 914 => to_unsigned(3807, 12), 915 => to_unsigned(2534, 12), 916 => to_unsigned(466, 12), 917 => to_unsigned(603, 12), 918 => to_unsigned(1789, 12), 919 => to_unsigned(474, 12), 920 => to_unsigned(1303, 12), 921 => to_unsigned(3271, 12), 922 => to_unsigned(2957, 12), 923 => to_unsigned(788, 12), 924 => to_unsigned(3550, 12), 925 => to_unsigned(3363, 12), 926 => to_unsigned(1994, 12), 927 => to_unsigned(419, 12), 928 => to_unsigned(2757, 12), 929 => to_unsigned(2853, 12), 930 => to_unsigned(1430, 12), 931 => to_unsigned(2721, 12), 932 => to_unsigned(18, 12), 933 => to_unsigned(896, 12), 934 => to_unsigned(3359, 12), 935 => to_unsigned(2540, 12), 936 => to_unsigned(3870, 12), 937 => to_unsigned(1197, 12), 938 => to_unsigned(1154, 12), 939 => to_unsigned(3221, 12), 940 => to_unsigned(1810, 12), 941 => to_unsigned(2384, 12), 942 => to_unsigned(611, 12), 943 => to_unsigned(4095, 12), 944 => to_unsigned(1804, 12), 945 => to_unsigned(3912, 12), 946 => to_unsigned(3452, 12), 947 => to_unsigned(4058, 12), 948 => to_unsigned(2748, 12), 949 => to_unsigned(99, 12), 950 => to_unsigned(2953, 12), 951 => to_unsigned(2079, 12), 952 => to_unsigned(3308, 12), 953 => to_unsigned(1073, 12), 954 => to_unsigned(3391, 12), 955 => to_unsigned(3179, 12), 956 => to_unsigned(3887, 12), 957 => to_unsigned(2944, 12), 958 => to_unsigned(4013, 12), 959 => to_unsigned(892, 12), 960 => to_unsigned(1846, 12), 961 => to_unsigned(4052, 12), 962 => to_unsigned(732, 12), 963 => to_unsigned(2854, 12), 964 => to_unsigned(2084, 12), 965 => to_unsigned(3486, 12), 966 => to_unsigned(3105, 12), 967 => to_unsigned(2147, 12), 968 => to_unsigned(3177, 12), 969 => to_unsigned(2678, 12), 970 => to_unsigned(382, 12), 971 => to_unsigned(538, 12), 972 => to_unsigned(1838, 12), 973 => to_unsigned(2066, 12), 974 => to_unsigned(2776, 12), 975 => to_unsigned(344, 12), 976 => to_unsigned(3534, 12), 977 => to_unsigned(1244, 12), 978 => to_unsigned(498, 12), 979 => to_unsigned(2601, 12), 980 => to_unsigned(1299, 12), 981 => to_unsigned(1794, 12), 982 => to_unsigned(298, 12), 983 => to_unsigned(561, 12), 984 => to_unsigned(3322, 12), 985 => to_unsigned(3741, 12), 986 => to_unsigned(3521, 12), 987 => to_unsigned(789, 12), 988 => to_unsigned(1910, 12), 989 => to_unsigned(1745, 12), 990 => to_unsigned(503, 12), 991 => to_unsigned(2905, 12), 992 => to_unsigned(78, 12), 993 => to_unsigned(1913, 12), 994 => to_unsigned(86, 12), 995 => to_unsigned(1231, 12), 996 => to_unsigned(754, 12), 997 => to_unsigned(466, 12), 998 => to_unsigned(4095, 12), 999 => to_unsigned(395, 12), 1000 => to_unsigned(3382, 12), 1001 => to_unsigned(280, 12), 1002 => to_unsigned(3909, 12), 1003 => to_unsigned(2283, 12), 1004 => to_unsigned(2566, 12), 1005 => to_unsigned(2621, 12), 1006 => to_unsigned(2089, 12), 1007 => to_unsigned(1212, 12), 1008 => to_unsigned(1131, 12), 1009 => to_unsigned(1711, 12), 1010 => to_unsigned(1420, 12), 1011 => to_unsigned(1676, 12), 1012 => to_unsigned(301, 12), 1013 => to_unsigned(549, 12), 1014 => to_unsigned(2386, 12), 1015 => to_unsigned(2505, 12), 1016 => to_unsigned(2248, 12), 1017 => to_unsigned(2357, 12), 1018 => to_unsigned(552, 12), 1019 => to_unsigned(3976, 12), 1020 => to_unsigned(3328, 12), 1021 => to_unsigned(2336, 12), 1022 => to_unsigned(3468, 12), 1023 => to_unsigned(3316, 12), 1024 => to_unsigned(3092, 12), 1025 => to_unsigned(1273, 12), 1026 => to_unsigned(3067, 12), 1027 => to_unsigned(3573, 12), 1028 => to_unsigned(2418, 12), 1029 => to_unsigned(2831, 12), 1030 => to_unsigned(791, 12), 1031 => to_unsigned(446, 12), 1032 => to_unsigned(2102, 12), 1033 => to_unsigned(3436, 12), 1034 => to_unsigned(4049, 12), 1035 => to_unsigned(3415, 12), 1036 => to_unsigned(1033, 12), 1037 => to_unsigned(2669, 12), 1038 => to_unsigned(1506, 12), 1039 => to_unsigned(480, 12), 1040 => to_unsigned(3945, 12), 1041 => to_unsigned(1606, 12), 1042 => to_unsigned(1015, 12), 1043 => to_unsigned(3547, 12), 1044 => to_unsigned(3747, 12), 1045 => to_unsigned(2771, 12), 1046 => to_unsigned(4006, 12), 1047 => to_unsigned(2369, 12), 1048 => to_unsigned(289, 12), 1049 => to_unsigned(2661, 12), 1050 => to_unsigned(3425, 12), 1051 => to_unsigned(929, 12), 1052 => to_unsigned(131, 12), 1053 => to_unsigned(854, 12), 1054 => to_unsigned(357, 12), 1055 => to_unsigned(3194, 12), 1056 => to_unsigned(690, 12), 1057 => to_unsigned(4001, 12), 1058 => to_unsigned(515, 12), 1059 => to_unsigned(333, 12), 1060 => to_unsigned(1442, 12), 1061 => to_unsigned(847, 12), 1062 => to_unsigned(2987, 12), 1063 => to_unsigned(481, 12), 1064 => to_unsigned(3102, 12), 1065 => to_unsigned(4009, 12), 1066 => to_unsigned(3996, 12), 1067 => to_unsigned(2697, 12), 1068 => to_unsigned(3851, 12), 1069 => to_unsigned(3225, 12), 1070 => to_unsigned(1776, 12), 1071 => to_unsigned(1276, 12), 1072 => to_unsigned(2361, 12), 1073 => to_unsigned(585, 12), 1074 => to_unsigned(1532, 12), 1075 => to_unsigned(1342, 12), 1076 => to_unsigned(2144, 12), 1077 => to_unsigned(1941, 12), 1078 => to_unsigned(996, 12), 1079 => to_unsigned(203, 12), 1080 => to_unsigned(1699, 12), 1081 => to_unsigned(1208, 12), 1082 => to_unsigned(2937, 12), 1083 => to_unsigned(1452, 12), 1084 => to_unsigned(1730, 12), 1085 => to_unsigned(2144, 12), 1086 => to_unsigned(2140, 12), 1087 => to_unsigned(1636, 12), 1088 => to_unsigned(2808, 12), 1089 => to_unsigned(2634, 12), 1090 => to_unsigned(2403, 12), 1091 => to_unsigned(2333, 12), 1092 => to_unsigned(1213, 12), 1093 => to_unsigned(3563, 12), 1094 => to_unsigned(41, 12), 1095 => to_unsigned(2007, 12), 1096 => to_unsigned(933, 12), 1097 => to_unsigned(703, 12), 1098 => to_unsigned(1181, 12), 1099 => to_unsigned(3425, 12), 1100 => to_unsigned(2301, 12), 1101 => to_unsigned(3107, 12), 1102 => to_unsigned(3818, 12), 1103 => to_unsigned(2256, 12), 1104 => to_unsigned(2132, 12), 1105 => to_unsigned(3105, 12), 1106 => to_unsigned(643, 12), 1107 => to_unsigned(2399, 12), 1108 => to_unsigned(3309, 12), 1109 => to_unsigned(1124, 12), 1110 => to_unsigned(3016, 12), 1111 => to_unsigned(3416, 12), 1112 => to_unsigned(702, 12), 1113 => to_unsigned(3609, 12), 1114 => to_unsigned(2905, 12), 1115 => to_unsigned(1317, 12), 1116 => to_unsigned(1738, 12), 1117 => to_unsigned(1248, 12), 1118 => to_unsigned(707, 12), 1119 => to_unsigned(3711, 12), 1120 => to_unsigned(2751, 12), 1121 => to_unsigned(1749, 12), 1122 => to_unsigned(1000, 12), 1123 => to_unsigned(589, 12), 1124 => to_unsigned(96, 12), 1125 => to_unsigned(3690, 12), 1126 => to_unsigned(3077, 12), 1127 => to_unsigned(2325, 12), 1128 => to_unsigned(1192, 12), 1129 => to_unsigned(1165, 12), 1130 => to_unsigned(27, 12), 1131 => to_unsigned(546, 12), 1132 => to_unsigned(1408, 12), 1133 => to_unsigned(1591, 12), 1134 => to_unsigned(761, 12), 1135 => to_unsigned(3116, 12), 1136 => to_unsigned(743, 12), 1137 => to_unsigned(1200, 12), 1138 => to_unsigned(367, 12), 1139 => to_unsigned(1331, 12), 1140 => to_unsigned(827, 12), 1141 => to_unsigned(529, 12), 1142 => to_unsigned(352, 12), 1143 => to_unsigned(1528, 12), 1144 => to_unsigned(3808, 12), 1145 => to_unsigned(1803, 12), 1146 => to_unsigned(1450, 12), 1147 => to_unsigned(710, 12), 1148 => to_unsigned(3282, 12), 1149 => to_unsigned(801, 12), 1150 => to_unsigned(3123, 12), 1151 => to_unsigned(2484, 12), 1152 => to_unsigned(3909, 12), 1153 => to_unsigned(81, 12), 1154 => to_unsigned(4022, 12), 1155 => to_unsigned(2314, 12), 1156 => to_unsigned(3276, 12), 1157 => to_unsigned(41, 12), 1158 => to_unsigned(3537, 12), 1159 => to_unsigned(1951, 12), 1160 => to_unsigned(259, 12), 1161 => to_unsigned(744, 12), 1162 => to_unsigned(1250, 12), 1163 => to_unsigned(3498, 12), 1164 => to_unsigned(1886, 12), 1165 => to_unsigned(2694, 12), 1166 => to_unsigned(3904, 12), 1167 => to_unsigned(4, 12), 1168 => to_unsigned(644, 12), 1169 => to_unsigned(575, 12), 1170 => to_unsigned(748, 12), 1171 => to_unsigned(3520, 12), 1172 => to_unsigned(4083, 12), 1173 => to_unsigned(1507, 12), 1174 => to_unsigned(1366, 12), 1175 => to_unsigned(2014, 12), 1176 => to_unsigned(1511, 12), 1177 => to_unsigned(2973, 12), 1178 => to_unsigned(790, 12), 1179 => to_unsigned(2135, 12), 1180 => to_unsigned(1329, 12), 1181 => to_unsigned(2842, 12), 1182 => to_unsigned(2166, 12), 1183 => to_unsigned(1848, 12), 1184 => to_unsigned(1163, 12), 1185 => to_unsigned(2946, 12), 1186 => to_unsigned(3029, 12), 1187 => to_unsigned(1036, 12), 1188 => to_unsigned(2000, 12), 1189 => to_unsigned(2, 12), 1190 => to_unsigned(2139, 12), 1191 => to_unsigned(716, 12), 1192 => to_unsigned(117, 12), 1193 => to_unsigned(2169, 12), 1194 => to_unsigned(2681, 12), 1195 => to_unsigned(1769, 12), 1196 => to_unsigned(3107, 12), 1197 => to_unsigned(3712, 12), 1198 => to_unsigned(1341, 12), 1199 => to_unsigned(3149, 12), 1200 => to_unsigned(511, 12), 1201 => to_unsigned(3685, 12), 1202 => to_unsigned(2450, 12), 1203 => to_unsigned(4003, 12), 1204 => to_unsigned(3594, 12), 1205 => to_unsigned(1299, 12), 1206 => to_unsigned(1772, 12), 1207 => to_unsigned(2715, 12), 1208 => to_unsigned(265, 12), 1209 => to_unsigned(624, 12), 1210 => to_unsigned(3494, 12), 1211 => to_unsigned(3962, 12), 1212 => to_unsigned(780, 12), 1213 => to_unsigned(3823, 12), 1214 => to_unsigned(3302, 12), 1215 => to_unsigned(1521, 12), 1216 => to_unsigned(102, 12), 1217 => to_unsigned(69, 12), 1218 => to_unsigned(342, 12), 1219 => to_unsigned(62, 12), 1220 => to_unsigned(3084, 12), 1221 => to_unsigned(1602, 12), 1222 => to_unsigned(59, 12), 1223 => to_unsigned(1920, 12), 1224 => to_unsigned(497, 12), 1225 => to_unsigned(3096, 12), 1226 => to_unsigned(362, 12), 1227 => to_unsigned(3805, 12), 1228 => to_unsigned(1500, 12), 1229 => to_unsigned(992, 12), 1230 => to_unsigned(3204, 12), 1231 => to_unsigned(4040, 12), 1232 => to_unsigned(1426, 12), 1233 => to_unsigned(813, 12), 1234 => to_unsigned(476, 12), 1235 => to_unsigned(199, 12), 1236 => to_unsigned(584, 12), 1237 => to_unsigned(2960, 12), 1238 => to_unsigned(1622, 12), 1239 => to_unsigned(3946, 12), 1240 => to_unsigned(79, 12), 1241 => to_unsigned(1919, 12), 1242 => to_unsigned(2324, 12), 1243 => to_unsigned(1584, 12), 1244 => to_unsigned(1493, 12), 1245 => to_unsigned(1623, 12), 1246 => to_unsigned(481, 12), 1247 => to_unsigned(2370, 12), 1248 => to_unsigned(1584, 12), 1249 => to_unsigned(1754, 12), 1250 => to_unsigned(2187, 12), 1251 => to_unsigned(2200, 12), 1252 => to_unsigned(2447, 12), 1253 => to_unsigned(2927, 12), 1254 => to_unsigned(1689, 12), 1255 => to_unsigned(1919, 12), 1256 => to_unsigned(1925, 12), 1257 => to_unsigned(2582, 12), 1258 => to_unsigned(310, 12), 1259 => to_unsigned(2867, 12), 1260 => to_unsigned(1186, 12), 1261 => to_unsigned(1181, 12), 1262 => to_unsigned(2188, 12), 1263 => to_unsigned(2348, 12), 1264 => to_unsigned(2874, 12), 1265 => to_unsigned(3964, 12), 1266 => to_unsigned(3348, 12), 1267 => to_unsigned(319, 12), 1268 => to_unsigned(942, 12), 1269 => to_unsigned(353, 12), 1270 => to_unsigned(587, 12), 1271 => to_unsigned(814, 12), 1272 => to_unsigned(2398, 12), 1273 => to_unsigned(1134, 12), 1274 => to_unsigned(2808, 12), 1275 => to_unsigned(1291, 12), 1276 => to_unsigned(3014, 12), 1277 => to_unsigned(1887, 12), 1278 => to_unsigned(1826, 12), 1279 => to_unsigned(3369, 12), 1280 => to_unsigned(149, 12), 1281 => to_unsigned(2762, 12), 1282 => to_unsigned(2139, 12), 1283 => to_unsigned(81, 12), 1284 => to_unsigned(1510, 12), 1285 => to_unsigned(1849, 12), 1286 => to_unsigned(390, 12), 1287 => to_unsigned(2955, 12), 1288 => to_unsigned(189, 12), 1289 => to_unsigned(368, 12), 1290 => to_unsigned(2013, 12), 1291 => to_unsigned(3533, 12), 1292 => to_unsigned(1902, 12), 1293 => to_unsigned(3731, 12), 1294 => to_unsigned(249, 12), 1295 => to_unsigned(1031, 12), 1296 => to_unsigned(1337, 12), 1297 => to_unsigned(656, 12), 1298 => to_unsigned(3910, 12), 1299 => to_unsigned(2216, 12), 1300 => to_unsigned(1999, 12), 1301 => to_unsigned(190, 12), 1302 => to_unsigned(3266, 12), 1303 => to_unsigned(1546, 12), 1304 => to_unsigned(297, 12), 1305 => to_unsigned(4010, 12), 1306 => to_unsigned(2472, 12), 1307 => to_unsigned(2973, 12), 1308 => to_unsigned(3146, 12), 1309 => to_unsigned(1354, 12), 1310 => to_unsigned(2719, 12), 1311 => to_unsigned(3665, 12), 1312 => to_unsigned(1019, 12), 1313 => to_unsigned(2915, 12), 1314 => to_unsigned(1956, 12), 1315 => to_unsigned(1508, 12), 1316 => to_unsigned(3133, 12), 1317 => to_unsigned(849, 12), 1318 => to_unsigned(1905, 12), 1319 => to_unsigned(469, 12), 1320 => to_unsigned(923, 12), 1321 => to_unsigned(3353, 12), 1322 => to_unsigned(1967, 12), 1323 => to_unsigned(1206, 12), 1324 => to_unsigned(3528, 12), 1325 => to_unsigned(4065, 12), 1326 => to_unsigned(1786, 12), 1327 => to_unsigned(3439, 12), 1328 => to_unsigned(3529, 12), 1329 => to_unsigned(1931, 12), 1330 => to_unsigned(2224, 12), 1331 => to_unsigned(3055, 12), 1332 => to_unsigned(604, 12), 1333 => to_unsigned(784, 12), 1334 => to_unsigned(2288, 12), 1335 => to_unsigned(962, 12), 1336 => to_unsigned(1224, 12), 1337 => to_unsigned(417, 12), 1338 => to_unsigned(3707, 12), 1339 => to_unsigned(2736, 12), 1340 => to_unsigned(398, 12), 1341 => to_unsigned(1704, 12), 1342 => to_unsigned(1345, 12), 1343 => to_unsigned(2734, 12), 1344 => to_unsigned(1247, 12), 1345 => to_unsigned(790, 12), 1346 => to_unsigned(3053, 12), 1347 => to_unsigned(192, 12), 1348 => to_unsigned(3788, 12), 1349 => to_unsigned(2216, 12), 1350 => to_unsigned(3832, 12), 1351 => to_unsigned(1535, 12), 1352 => to_unsigned(1472, 12), 1353 => to_unsigned(2012, 12), 1354 => to_unsigned(2207, 12), 1355 => to_unsigned(1084, 12), 1356 => to_unsigned(1406, 12), 1357 => to_unsigned(2332, 12), 1358 => to_unsigned(3196, 12), 1359 => to_unsigned(1528, 12), 1360 => to_unsigned(1721, 12), 1361 => to_unsigned(3155, 12), 1362 => to_unsigned(2035, 12), 1363 => to_unsigned(3168, 12), 1364 => to_unsigned(1130, 12), 1365 => to_unsigned(2347, 12), 1366 => to_unsigned(503, 12), 1367 => to_unsigned(3652, 12), 1368 => to_unsigned(3570, 12), 1369 => to_unsigned(2769, 12), 1370 => to_unsigned(3165, 12), 1371 => to_unsigned(2534, 12), 1372 => to_unsigned(1562, 12), 1373 => to_unsigned(3801, 12), 1374 => to_unsigned(3026, 12), 1375 => to_unsigned(3507, 12), 1376 => to_unsigned(2900, 12), 1377 => to_unsigned(3375, 12), 1378 => to_unsigned(3897, 12), 1379 => to_unsigned(1065, 12), 1380 => to_unsigned(455, 12), 1381 => to_unsigned(3298, 12), 1382 => to_unsigned(412, 12), 1383 => to_unsigned(2720, 12), 1384 => to_unsigned(1521, 12), 1385 => to_unsigned(3558, 12), 1386 => to_unsigned(2700, 12), 1387 => to_unsigned(3672, 12), 1388 => to_unsigned(1134, 12), 1389 => to_unsigned(3566, 12), 1390 => to_unsigned(199, 12), 1391 => to_unsigned(457, 12), 1392 => to_unsigned(4028, 12), 1393 => to_unsigned(1319, 12), 1394 => to_unsigned(3373, 12), 1395 => to_unsigned(161, 12), 1396 => to_unsigned(1118, 12), 1397 => to_unsigned(2019, 12), 1398 => to_unsigned(3132, 12), 1399 => to_unsigned(1954, 12), 1400 => to_unsigned(3047, 12), 1401 => to_unsigned(1474, 12), 1402 => to_unsigned(1181, 12), 1403 => to_unsigned(3960, 12), 1404 => to_unsigned(1191, 12), 1405 => to_unsigned(3903, 12), 1406 => to_unsigned(3734, 12), 1407 => to_unsigned(739, 12), 1408 => to_unsigned(53, 12), 1409 => to_unsigned(2752, 12), 1410 => to_unsigned(2074, 12), 1411 => to_unsigned(2116, 12), 1412 => to_unsigned(1525, 12), 1413 => to_unsigned(2091, 12), 1414 => to_unsigned(3503, 12), 1415 => to_unsigned(2185, 12), 1416 => to_unsigned(582, 12), 1417 => to_unsigned(1949, 12), 1418 => to_unsigned(2053, 12), 1419 => to_unsigned(1537, 12), 1420 => to_unsigned(892, 12), 1421 => to_unsigned(3670, 12), 1422 => to_unsigned(26, 12), 1423 => to_unsigned(3933, 12), 1424 => to_unsigned(3717, 12), 1425 => to_unsigned(2448, 12), 1426 => to_unsigned(3994, 12), 1427 => to_unsigned(300, 12), 1428 => to_unsigned(282, 12), 1429 => to_unsigned(2126, 12), 1430 => to_unsigned(2904, 12), 1431 => to_unsigned(2696, 12), 1432 => to_unsigned(3859, 12), 1433 => to_unsigned(4061, 12), 1434 => to_unsigned(2935, 12), 1435 => to_unsigned(1339, 12), 1436 => to_unsigned(1099, 12), 1437 => to_unsigned(2222, 12), 1438 => to_unsigned(789, 12), 1439 => to_unsigned(450, 12), 1440 => to_unsigned(1213, 12), 1441 => to_unsigned(3129, 12), 1442 => to_unsigned(2458, 12), 1443 => to_unsigned(1077, 12), 1444 => to_unsigned(2416, 12), 1445 => to_unsigned(4075, 12), 1446 => to_unsigned(452, 12), 1447 => to_unsigned(2169, 12), 1448 => to_unsigned(918, 12), 1449 => to_unsigned(2386, 12), 1450 => to_unsigned(2726, 12), 1451 => to_unsigned(449, 12), 1452 => to_unsigned(1668, 12), 1453 => to_unsigned(3197, 12), 1454 => to_unsigned(3303, 12), 1455 => to_unsigned(1427, 12), 1456 => to_unsigned(859, 12), 1457 => to_unsigned(1415, 12), 1458 => to_unsigned(2416, 12), 1459 => to_unsigned(1397, 12), 1460 => to_unsigned(2525, 12), 1461 => to_unsigned(1890, 12), 1462 => to_unsigned(856, 12), 1463 => to_unsigned(825, 12), 1464 => to_unsigned(3532, 12), 1465 => to_unsigned(1349, 12), 1466 => to_unsigned(556, 12), 1467 => to_unsigned(1037, 12), 1468 => to_unsigned(2544, 12), 1469 => to_unsigned(3494, 12), 1470 => to_unsigned(207, 12), 1471 => to_unsigned(1024, 12), 1472 => to_unsigned(2161, 12), 1473 => to_unsigned(1459, 12), 1474 => to_unsigned(1732, 12), 1475 => to_unsigned(3117, 12), 1476 => to_unsigned(662, 12), 1477 => to_unsigned(3870, 12), 1478 => to_unsigned(3581, 12), 1479 => to_unsigned(2592, 12), 1480 => to_unsigned(631, 12), 1481 => to_unsigned(607, 12), 1482 => to_unsigned(3117, 12), 1483 => to_unsigned(2148, 12), 1484 => to_unsigned(1923, 12), 1485 => to_unsigned(2748, 12), 1486 => to_unsigned(2979, 12), 1487 => to_unsigned(19, 12), 1488 => to_unsigned(1634, 12), 1489 => to_unsigned(3729, 12), 1490 => to_unsigned(2284, 12), 1491 => to_unsigned(2307, 12), 1492 => to_unsigned(3772, 12), 1493 => to_unsigned(3528, 12), 1494 => to_unsigned(2113, 12), 1495 => to_unsigned(1679, 12), 1496 => to_unsigned(873, 12), 1497 => to_unsigned(2312, 12), 1498 => to_unsigned(376, 12), 1499 => to_unsigned(2356, 12), 1500 => to_unsigned(2966, 12), 1501 => to_unsigned(2058, 12), 1502 => to_unsigned(1068, 12), 1503 => to_unsigned(2188, 12), 1504 => to_unsigned(3075, 12), 1505 => to_unsigned(1302, 12), 1506 => to_unsigned(652, 12), 1507 => to_unsigned(3737, 12), 1508 => to_unsigned(3765, 12), 1509 => to_unsigned(3162, 12), 1510 => to_unsigned(552, 12), 1511 => to_unsigned(169, 12), 1512 => to_unsigned(1664, 12), 1513 => to_unsigned(3767, 12), 1514 => to_unsigned(1083, 12), 1515 => to_unsigned(3814, 12), 1516 => to_unsigned(1204, 12), 1517 => to_unsigned(2203, 12), 1518 => to_unsigned(3624, 12), 1519 => to_unsigned(3556, 12), 1520 => to_unsigned(2773, 12), 1521 => to_unsigned(1045, 12), 1522 => to_unsigned(3526, 12), 1523 => to_unsigned(1100, 12), 1524 => to_unsigned(2695, 12), 1525 => to_unsigned(1155, 12), 1526 => to_unsigned(2552, 12), 1527 => to_unsigned(970, 12), 1528 => to_unsigned(2075, 12), 1529 => to_unsigned(2745, 12), 1530 => to_unsigned(2289, 12), 1531 => to_unsigned(3569, 12), 1532 => to_unsigned(2392, 12), 1533 => to_unsigned(177, 12), 1534 => to_unsigned(3246, 12), 1535 => to_unsigned(3785, 12), 1536 => to_unsigned(2540, 12), 1537 => to_unsigned(2028, 12), 1538 => to_unsigned(36, 12), 1539 => to_unsigned(520, 12), 1540 => to_unsigned(1417, 12), 1541 => to_unsigned(483, 12), 1542 => to_unsigned(2433, 12), 1543 => to_unsigned(2726, 12), 1544 => to_unsigned(1428, 12), 1545 => to_unsigned(3117, 12), 1546 => to_unsigned(3929, 12), 1547 => to_unsigned(172, 12), 1548 => to_unsigned(2649, 12), 1549 => to_unsigned(965, 12), 1550 => to_unsigned(2368, 12), 1551 => to_unsigned(4094, 12), 1552 => to_unsigned(103, 12), 1553 => to_unsigned(3386, 12), 1554 => to_unsigned(3014, 12), 1555 => to_unsigned(2374, 12), 1556 => to_unsigned(615, 12), 1557 => to_unsigned(2802, 12), 1558 => to_unsigned(529, 12), 1559 => to_unsigned(1803, 12), 1560 => to_unsigned(17, 12), 1561 => to_unsigned(2853, 12), 1562 => to_unsigned(1630, 12), 1563 => to_unsigned(3257, 12), 1564 => to_unsigned(1010, 12), 1565 => to_unsigned(1905, 12), 1566 => to_unsigned(2761, 12), 1567 => to_unsigned(780, 12), 1568 => to_unsigned(3985, 12), 1569 => to_unsigned(2686, 12), 1570 => to_unsigned(1828, 12), 1571 => to_unsigned(672, 12), 1572 => to_unsigned(1407, 12), 1573 => to_unsigned(2947, 12), 1574 => to_unsigned(2553, 12), 1575 => to_unsigned(3958, 12), 1576 => to_unsigned(4044, 12), 1577 => to_unsigned(2165, 12), 1578 => to_unsigned(3311, 12), 1579 => to_unsigned(677, 12), 1580 => to_unsigned(1524, 12), 1581 => to_unsigned(3783, 12), 1582 => to_unsigned(238, 12), 1583 => to_unsigned(1725, 12), 1584 => to_unsigned(1541, 12), 1585 => to_unsigned(145, 12), 1586 => to_unsigned(1298, 12), 1587 => to_unsigned(3602, 12), 1588 => to_unsigned(1873, 12), 1589 => to_unsigned(2593, 12), 1590 => to_unsigned(2698, 12), 1591 => to_unsigned(305, 12), 1592 => to_unsigned(3593, 12), 1593 => to_unsigned(666, 12), 1594 => to_unsigned(2180, 12), 1595 => to_unsigned(872, 12), 1596 => to_unsigned(1625, 12), 1597 => to_unsigned(114, 12), 1598 => to_unsigned(2277, 12), 1599 => to_unsigned(3399, 12), 1600 => to_unsigned(3425, 12), 1601 => to_unsigned(1809, 12), 1602 => to_unsigned(764, 12), 1603 => to_unsigned(1519, 12), 1604 => to_unsigned(1511, 12), 1605 => to_unsigned(2672, 12), 1606 => to_unsigned(1041, 12), 1607 => to_unsigned(1894, 12), 1608 => to_unsigned(1736, 12), 1609 => to_unsigned(614, 12), 1610 => to_unsigned(570, 12), 1611 => to_unsigned(3159, 12), 1612 => to_unsigned(951, 12), 1613 => to_unsigned(2210, 12), 1614 => to_unsigned(3813, 12), 1615 => to_unsigned(4059, 12), 1616 => to_unsigned(3780, 12), 1617 => to_unsigned(2690, 12), 1618 => to_unsigned(2541, 12), 1619 => to_unsigned(3953, 12), 1620 => to_unsigned(793, 12), 1621 => to_unsigned(1350, 12), 1622 => to_unsigned(2186, 12), 1623 => to_unsigned(531, 12), 1624 => to_unsigned(1965, 12), 1625 => to_unsigned(1871, 12), 1626 => to_unsigned(2132, 12), 1627 => to_unsigned(3509, 12), 1628 => to_unsigned(4047, 12), 1629 => to_unsigned(182, 12), 1630 => to_unsigned(3875, 12), 1631 => to_unsigned(1967, 12), 1632 => to_unsigned(1735, 12), 1633 => to_unsigned(2920, 12), 1634 => to_unsigned(828, 12), 1635 => to_unsigned(1572, 12), 1636 => to_unsigned(3697, 12), 1637 => to_unsigned(3996, 12), 1638 => to_unsigned(428, 12), 1639 => to_unsigned(3630, 12), 1640 => to_unsigned(3465, 12), 1641 => to_unsigned(2404, 12), 1642 => to_unsigned(1111, 12), 1643 => to_unsigned(2211, 12), 1644 => to_unsigned(1116, 12), 1645 => to_unsigned(1042, 12), 1646 => to_unsigned(2638, 12), 1647 => to_unsigned(3815, 12), 1648 => to_unsigned(3220, 12), 1649 => to_unsigned(2084, 12), 1650 => to_unsigned(1864, 12), 1651 => to_unsigned(1392, 12), 1652 => to_unsigned(871, 12), 1653 => to_unsigned(525, 12), 1654 => to_unsigned(2039, 12), 1655 => to_unsigned(619, 12), 1656 => to_unsigned(3560, 12), 1657 => to_unsigned(1301, 12), 1658 => to_unsigned(315, 12), 1659 => to_unsigned(1263, 12), 1660 => to_unsigned(3261, 12), 1661 => to_unsigned(3552, 12), 1662 => to_unsigned(2336, 12), 1663 => to_unsigned(30, 12), 1664 => to_unsigned(1609, 12), 1665 => to_unsigned(2139, 12), 1666 => to_unsigned(2493, 12), 1667 => to_unsigned(3996, 12), 1668 => to_unsigned(2872, 12), 1669 => to_unsigned(3051, 12), 1670 => to_unsigned(2839, 12), 1671 => to_unsigned(1372, 12), 1672 => to_unsigned(4024, 12), 1673 => to_unsigned(3394, 12), 1674 => to_unsigned(788, 12), 1675 => to_unsigned(1366, 12), 1676 => to_unsigned(2656, 12), 1677 => to_unsigned(2951, 12), 1678 => to_unsigned(3512, 12), 1679 => to_unsigned(2325, 12), 1680 => to_unsigned(596, 12), 1681 => to_unsigned(2963, 12), 1682 => to_unsigned(857, 12), 1683 => to_unsigned(1199, 12), 1684 => to_unsigned(1445, 12), 1685 => to_unsigned(2136, 12), 1686 => to_unsigned(851, 12), 1687 => to_unsigned(2487, 12), 1688 => to_unsigned(682, 12), 1689 => to_unsigned(1549, 12), 1690 => to_unsigned(3500, 12), 1691 => to_unsigned(2651, 12), 1692 => to_unsigned(1366, 12), 1693 => to_unsigned(1371, 12), 1694 => to_unsigned(2691, 12), 1695 => to_unsigned(1465, 12), 1696 => to_unsigned(161, 12), 1697 => to_unsigned(2845, 12), 1698 => to_unsigned(3413, 12), 1699 => to_unsigned(3138, 12), 1700 => to_unsigned(3110, 12), 1701 => to_unsigned(1432, 12), 1702 => to_unsigned(209, 12), 1703 => to_unsigned(2637, 12), 1704 => to_unsigned(3529, 12), 1705 => to_unsigned(3817, 12), 1706 => to_unsigned(3609, 12), 1707 => to_unsigned(3109, 12), 1708 => to_unsigned(2830, 12), 1709 => to_unsigned(925, 12), 1710 => to_unsigned(2415, 12), 1711 => to_unsigned(903, 12), 1712 => to_unsigned(1338, 12), 1713 => to_unsigned(1947, 12), 1714 => to_unsigned(1948, 12), 1715 => to_unsigned(854, 12), 1716 => to_unsigned(1092, 12), 1717 => to_unsigned(4035, 12), 1718 => to_unsigned(280, 12), 1719 => to_unsigned(3303, 12), 1720 => to_unsigned(3226, 12), 1721 => to_unsigned(1274, 12), 1722 => to_unsigned(3721, 12), 1723 => to_unsigned(3003, 12), 1724 => to_unsigned(873, 12), 1725 => to_unsigned(3316, 12), 1726 => to_unsigned(2231, 12), 1727 => to_unsigned(3911, 12), 1728 => to_unsigned(1620, 12), 1729 => to_unsigned(1419, 12), 1730 => to_unsigned(198, 12), 1731 => to_unsigned(348, 12), 1732 => to_unsigned(2925, 12), 1733 => to_unsigned(258, 12), 1734 => to_unsigned(2215, 12), 1735 => to_unsigned(1593, 12), 1736 => to_unsigned(2298, 12), 1737 => to_unsigned(2971, 12), 1738 => to_unsigned(415, 12), 1739 => to_unsigned(2979, 12), 1740 => to_unsigned(3212, 12), 1741 => to_unsigned(3904, 12), 1742 => to_unsigned(767, 12), 1743 => to_unsigned(663, 12), 1744 => to_unsigned(1669, 12), 1745 => to_unsigned(1719, 12), 1746 => to_unsigned(192, 12), 1747 => to_unsigned(803, 12), 1748 => to_unsigned(1407, 12), 1749 => to_unsigned(2058, 12), 1750 => to_unsigned(3741, 12), 1751 => to_unsigned(2367, 12), 1752 => to_unsigned(4049, 12), 1753 => to_unsigned(1840, 12), 1754 => to_unsigned(2024, 12), 1755 => to_unsigned(2258, 12), 1756 => to_unsigned(2619, 12), 1757 => to_unsigned(116, 12), 1758 => to_unsigned(175, 12), 1759 => to_unsigned(1981, 12), 1760 => to_unsigned(1162, 12), 1761 => to_unsigned(1171, 12), 1762 => to_unsigned(3813, 12), 1763 => to_unsigned(3149, 12), 1764 => to_unsigned(2233, 12), 1765 => to_unsigned(1987, 12), 1766 => to_unsigned(3620, 12), 1767 => to_unsigned(1539, 12), 1768 => to_unsigned(3491, 12), 1769 => to_unsigned(967, 12), 1770 => to_unsigned(2806, 12), 1771 => to_unsigned(3914, 12), 1772 => to_unsigned(3156, 12), 1773 => to_unsigned(2908, 12), 1774 => to_unsigned(3656, 12), 1775 => to_unsigned(1032, 12), 1776 => to_unsigned(465, 12), 1777 => to_unsigned(2001, 12), 1778 => to_unsigned(1404, 12), 1779 => to_unsigned(3781, 12), 1780 => to_unsigned(4063, 12), 1781 => to_unsigned(1245, 12), 1782 => to_unsigned(1979, 12), 1783 => to_unsigned(720, 12), 1784 => to_unsigned(441, 12), 1785 => to_unsigned(3444, 12), 1786 => to_unsigned(854, 12), 1787 => to_unsigned(739, 12), 1788 => to_unsigned(1586, 12), 1789 => to_unsigned(867, 12), 1790 => to_unsigned(592, 12), 1791 => to_unsigned(117, 12), 1792 => to_unsigned(2459, 12), 1793 => to_unsigned(2656, 12), 1794 => to_unsigned(1327, 12), 1795 => to_unsigned(450, 12), 1796 => to_unsigned(11, 12), 1797 => to_unsigned(1106, 12), 1798 => to_unsigned(216, 12), 1799 => to_unsigned(3608, 12), 1800 => to_unsigned(2176, 12), 1801 => to_unsigned(621, 12), 1802 => to_unsigned(3516, 12), 1803 => to_unsigned(1224, 12), 1804 => to_unsigned(2135, 12), 1805 => to_unsigned(513, 12), 1806 => to_unsigned(1275, 12), 1807 => to_unsigned(349, 12), 1808 => to_unsigned(47, 12), 1809 => to_unsigned(3686, 12), 1810 => to_unsigned(2278, 12), 1811 => to_unsigned(1260, 12), 1812 => to_unsigned(3058, 12), 1813 => to_unsigned(434, 12), 1814 => to_unsigned(977, 12), 1815 => to_unsigned(2259, 12), 1816 => to_unsigned(2173, 12), 1817 => to_unsigned(1753, 12), 1818 => to_unsigned(3710, 12), 1819 => to_unsigned(965, 12), 1820 => to_unsigned(507, 12), 1821 => to_unsigned(750, 12), 1822 => to_unsigned(1877, 12), 1823 => to_unsigned(546, 12), 1824 => to_unsigned(3553, 12), 1825 => to_unsigned(2854, 12), 1826 => to_unsigned(1778, 12), 1827 => to_unsigned(2943, 12), 1828 => to_unsigned(3547, 12), 1829 => to_unsigned(361, 12), 1830 => to_unsigned(3045, 12), 1831 => to_unsigned(817, 12), 1832 => to_unsigned(2556, 12), 1833 => to_unsigned(1924, 12), 1834 => to_unsigned(211, 12), 1835 => to_unsigned(2867, 12), 1836 => to_unsigned(801, 12), 1837 => to_unsigned(853, 12), 1838 => to_unsigned(3204, 12), 1839 => to_unsigned(3507, 12), 1840 => to_unsigned(1753, 12), 1841 => to_unsigned(2941, 12), 1842 => to_unsigned(2291, 12), 1843 => to_unsigned(71, 12), 1844 => to_unsigned(1464, 12), 1845 => to_unsigned(1662, 12), 1846 => to_unsigned(1828, 12), 1847 => to_unsigned(2611, 12), 1848 => to_unsigned(223, 12), 1849 => to_unsigned(2109, 12), 1850 => to_unsigned(701, 12), 1851 => to_unsigned(1391, 12), 1852 => to_unsigned(706, 12), 1853 => to_unsigned(3001, 12), 1854 => to_unsigned(1177, 12), 1855 => to_unsigned(1932, 12), 1856 => to_unsigned(1780, 12), 1857 => to_unsigned(4029, 12), 1858 => to_unsigned(1913, 12), 1859 => to_unsigned(381, 12), 1860 => to_unsigned(1925, 12), 1861 => to_unsigned(2723, 12), 1862 => to_unsigned(3294, 12), 1863 => to_unsigned(1268, 12), 1864 => to_unsigned(1716, 12), 1865 => to_unsigned(2697, 12), 1866 => to_unsigned(3121, 12), 1867 => to_unsigned(4083, 12), 1868 => to_unsigned(1489, 12), 1869 => to_unsigned(1208, 12), 1870 => to_unsigned(2205, 12), 1871 => to_unsigned(2251, 12), 1872 => to_unsigned(3261, 12), 1873 => to_unsigned(3490, 12), 1874 => to_unsigned(2027, 12), 1875 => to_unsigned(1272, 12), 1876 => to_unsigned(2938, 12), 1877 => to_unsigned(939, 12), 1878 => to_unsigned(801, 12), 1879 => to_unsigned(2938, 12), 1880 => to_unsigned(1534, 12), 1881 => to_unsigned(2204, 12), 1882 => to_unsigned(2582, 12), 1883 => to_unsigned(2137, 12), 1884 => to_unsigned(2011, 12), 1885 => to_unsigned(1041, 12), 1886 => to_unsigned(1791, 12), 1887 => to_unsigned(1057, 12), 1888 => to_unsigned(609, 12), 1889 => to_unsigned(1012, 12), 1890 => to_unsigned(2649, 12), 1891 => to_unsigned(3540, 12), 1892 => to_unsigned(3451, 12), 1893 => to_unsigned(1031, 12), 1894 => to_unsigned(2240, 12), 1895 => to_unsigned(268, 12), 1896 => to_unsigned(241, 12), 1897 => to_unsigned(1351, 12), 1898 => to_unsigned(4012, 12), 1899 => to_unsigned(3671, 12), 1900 => to_unsigned(1574, 12), 1901 => to_unsigned(2050, 12), 1902 => to_unsigned(1979, 12), 1903 => to_unsigned(1609, 12), 1904 => to_unsigned(2974, 12), 1905 => to_unsigned(1214, 12), 1906 => to_unsigned(1330, 12), 1907 => to_unsigned(3738, 12), 1908 => to_unsigned(3596, 12), 1909 => to_unsigned(2962, 12), 1910 => to_unsigned(3559, 12), 1911 => to_unsigned(3825, 12), 1912 => to_unsigned(413, 12), 1913 => to_unsigned(2234, 12), 1914 => to_unsigned(1006, 12), 1915 => to_unsigned(2982, 12), 1916 => to_unsigned(2807, 12), 1917 => to_unsigned(3398, 12), 1918 => to_unsigned(66, 12), 1919 => to_unsigned(3708, 12), 1920 => to_unsigned(2353, 12), 1921 => to_unsigned(3533, 12), 1922 => to_unsigned(2296, 12), 1923 => to_unsigned(3763, 12), 1924 => to_unsigned(4095, 12), 1925 => to_unsigned(1872, 12), 1926 => to_unsigned(1823, 12), 1927 => to_unsigned(3720, 12), 1928 => to_unsigned(873, 12), 1929 => to_unsigned(871, 12), 1930 => to_unsigned(1695, 12), 1931 => to_unsigned(3993, 12), 1932 => to_unsigned(1042, 12), 1933 => to_unsigned(2003, 12), 1934 => to_unsigned(860, 12), 1935 => to_unsigned(2881, 12), 1936 => to_unsigned(441, 12), 1937 => to_unsigned(2394, 12), 1938 => to_unsigned(3187, 12), 1939 => to_unsigned(414, 12), 1940 => to_unsigned(405, 12), 1941 => to_unsigned(884, 12), 1942 => to_unsigned(2891, 12), 1943 => to_unsigned(3363, 12), 1944 => to_unsigned(2018, 12), 1945 => to_unsigned(1661, 12), 1946 => to_unsigned(3254, 12), 1947 => to_unsigned(832, 12), 1948 => to_unsigned(761, 12), 1949 => to_unsigned(2623, 12), 1950 => to_unsigned(2776, 12), 1951 => to_unsigned(174, 12), 1952 => to_unsigned(608, 12), 1953 => to_unsigned(2216, 12), 1954 => to_unsigned(3642, 12), 1955 => to_unsigned(324, 12), 1956 => to_unsigned(3485, 12), 1957 => to_unsigned(3123, 12), 1958 => to_unsigned(1078, 12), 1959 => to_unsigned(56, 12), 1960 => to_unsigned(4084, 12), 1961 => to_unsigned(3922, 12), 1962 => to_unsigned(3636, 12), 1963 => to_unsigned(1125, 12), 1964 => to_unsigned(3559, 12), 1965 => to_unsigned(2114, 12), 1966 => to_unsigned(883, 12), 1967 => to_unsigned(545, 12), 1968 => to_unsigned(985, 12), 1969 => to_unsigned(2971, 12), 1970 => to_unsigned(2925, 12), 1971 => to_unsigned(3542, 12), 1972 => to_unsigned(1834, 12), 1973 => to_unsigned(1905, 12), 1974 => to_unsigned(1030, 12), 1975 => to_unsigned(2997, 12), 1976 => to_unsigned(1629, 12), 1977 => to_unsigned(2080, 12), 1978 => to_unsigned(3943, 12), 1979 => to_unsigned(3479, 12), 1980 => to_unsigned(2213, 12), 1981 => to_unsigned(1674, 12), 1982 => to_unsigned(1929, 12), 1983 => to_unsigned(2369, 12), 1984 => to_unsigned(832, 12), 1985 => to_unsigned(515, 12), 1986 => to_unsigned(2713, 12), 1987 => to_unsigned(2237, 12), 1988 => to_unsigned(1640, 12), 1989 => to_unsigned(716, 12), 1990 => to_unsigned(195, 12), 1991 => to_unsigned(1762, 12), 1992 => to_unsigned(219, 12), 1993 => to_unsigned(3121, 12), 1994 => to_unsigned(513, 12), 1995 => to_unsigned(2824, 12), 1996 => to_unsigned(102, 12), 1997 => to_unsigned(97, 12), 1998 => to_unsigned(2411, 12), 1999 => to_unsigned(95, 12), 2000 => to_unsigned(669, 12), 2001 => to_unsigned(3632, 12), 2002 => to_unsigned(1212, 12), 2003 => to_unsigned(3836, 12), 2004 => to_unsigned(2413, 12), 2005 => to_unsigned(2253, 12), 2006 => to_unsigned(4046, 12), 2007 => to_unsigned(3740, 12), 2008 => to_unsigned(3152, 12), 2009 => to_unsigned(1763, 12), 2010 => to_unsigned(88, 12), 2011 => to_unsigned(2349, 12), 2012 => to_unsigned(3462, 12), 2013 => to_unsigned(2322, 12), 2014 => to_unsigned(1336, 12), 2015 => to_unsigned(673, 12), 2016 => to_unsigned(4092, 12), 2017 => to_unsigned(2568, 12), 2018 => to_unsigned(846, 12), 2019 => to_unsigned(1170, 12), 2020 => to_unsigned(2537, 12), 2021 => to_unsigned(699, 12), 2022 => to_unsigned(3623, 12), 2023 => to_unsigned(1688, 12), 2024 => to_unsigned(1932, 12), 2025 => to_unsigned(1545, 12), 2026 => to_unsigned(3568, 12), 2027 => to_unsigned(3425, 12), 2028 => to_unsigned(255, 12), 2029 => to_unsigned(2481, 12), 2030 => to_unsigned(1377, 12), 2031 => to_unsigned(2610, 12), 2032 => to_unsigned(728, 12), 2033 => to_unsigned(1423, 12), 2034 => to_unsigned(1262, 12), 2035 => to_unsigned(3239, 12), 2036 => to_unsigned(2374, 12), 2037 => to_unsigned(2877, 12), 2038 => to_unsigned(401, 12), 2039 => to_unsigned(3976, 12), 2040 => to_unsigned(111, 12), 2041 => to_unsigned(1473, 12), 2042 => to_unsigned(2695, 12), 2043 => to_unsigned(2324, 12), 2044 => to_unsigned(2728, 12), 2045 => to_unsigned(1096, 12), 2046 => to_unsigned(1396, 12), 2047 => to_unsigned(3200, 12)),
            4 => (0 => to_unsigned(2935, 12), 1 => to_unsigned(1577, 12), 2 => to_unsigned(898, 12), 3 => to_unsigned(3104, 12), 4 => to_unsigned(2518, 12), 5 => to_unsigned(2428, 12), 6 => to_unsigned(522, 12), 7 => to_unsigned(2014, 12), 8 => to_unsigned(904, 12), 9 => to_unsigned(3093, 12), 10 => to_unsigned(3703, 12), 11 => to_unsigned(2617, 12), 12 => to_unsigned(2605, 12), 13 => to_unsigned(2371, 12), 14 => to_unsigned(2245, 12), 15 => to_unsigned(2331, 12), 16 => to_unsigned(2266, 12), 17 => to_unsigned(1420, 12), 18 => to_unsigned(3392, 12), 19 => to_unsigned(2051, 12), 20 => to_unsigned(3005, 12), 21 => to_unsigned(1451, 12), 22 => to_unsigned(1632, 12), 23 => to_unsigned(2600, 12), 24 => to_unsigned(3092, 12), 25 => to_unsigned(1806, 12), 26 => to_unsigned(3608, 12), 27 => to_unsigned(2883, 12), 28 => to_unsigned(1312, 12), 29 => to_unsigned(3401, 12), 30 => to_unsigned(1350, 12), 31 => to_unsigned(67, 12), 32 => to_unsigned(3898, 12), 33 => to_unsigned(3484, 12), 34 => to_unsigned(1539, 12), 35 => to_unsigned(2511, 12), 36 => to_unsigned(3296, 12), 37 => to_unsigned(1446, 12), 38 => to_unsigned(620, 12), 39 => to_unsigned(1884, 12), 40 => to_unsigned(1013, 12), 41 => to_unsigned(2802, 12), 42 => to_unsigned(3781, 12), 43 => to_unsigned(1, 12), 44 => to_unsigned(1169, 12), 45 => to_unsigned(2238, 12), 46 => to_unsigned(431, 12), 47 => to_unsigned(2312, 12), 48 => to_unsigned(3401, 12), 49 => to_unsigned(436, 12), 50 => to_unsigned(1933, 12), 51 => to_unsigned(2928, 12), 52 => to_unsigned(553, 12), 53 => to_unsigned(2072, 12), 54 => to_unsigned(2623, 12), 55 => to_unsigned(1988, 12), 56 => to_unsigned(1095, 12), 57 => to_unsigned(1093, 12), 58 => to_unsigned(3687, 12), 59 => to_unsigned(2708, 12), 60 => to_unsigned(3907, 12), 61 => to_unsigned(3521, 12), 62 => to_unsigned(3273, 12), 63 => to_unsigned(346, 12), 64 => to_unsigned(1857, 12), 65 => to_unsigned(2216, 12), 66 => to_unsigned(368, 12), 67 => to_unsigned(358, 12), 68 => to_unsigned(2990, 12), 69 => to_unsigned(405, 12), 70 => to_unsigned(3404, 12), 71 => to_unsigned(2118, 12), 72 => to_unsigned(2464, 12), 73 => to_unsigned(426, 12), 74 => to_unsigned(1876, 12), 75 => to_unsigned(3788, 12), 76 => to_unsigned(3414, 12), 77 => to_unsigned(3092, 12), 78 => to_unsigned(109, 12), 79 => to_unsigned(1953, 12), 80 => to_unsigned(4000, 12), 81 => to_unsigned(777, 12), 82 => to_unsigned(3259, 12), 83 => to_unsigned(612, 12), 84 => to_unsigned(4095, 12), 85 => to_unsigned(3203, 12), 86 => to_unsigned(745, 12), 87 => to_unsigned(3647, 12), 88 => to_unsigned(2110, 12), 89 => to_unsigned(2440, 12), 90 => to_unsigned(2332, 12), 91 => to_unsigned(1267, 12), 92 => to_unsigned(3085, 12), 93 => to_unsigned(1495, 12), 94 => to_unsigned(1863, 12), 95 => to_unsigned(382, 12), 96 => to_unsigned(1535, 12), 97 => to_unsigned(2675, 12), 98 => to_unsigned(2444, 12), 99 => to_unsigned(1922, 12), 100 => to_unsigned(1764, 12), 101 => to_unsigned(109, 12), 102 => to_unsigned(2637, 12), 103 => to_unsigned(3351, 12), 104 => to_unsigned(2942, 12), 105 => to_unsigned(2279, 12), 106 => to_unsigned(1211, 12), 107 => to_unsigned(1273, 12), 108 => to_unsigned(2166, 12), 109 => to_unsigned(2249, 12), 110 => to_unsigned(231, 12), 111 => to_unsigned(1918, 12), 112 => to_unsigned(1871, 12), 113 => to_unsigned(11, 12), 114 => to_unsigned(2057, 12), 115 => to_unsigned(3902, 12), 116 => to_unsigned(2625, 12), 117 => to_unsigned(218, 12), 118 => to_unsigned(1419, 12), 119 => to_unsigned(2911, 12), 120 => to_unsigned(3888, 12), 121 => to_unsigned(3386, 12), 122 => to_unsigned(2123, 12), 123 => to_unsigned(129, 12), 124 => to_unsigned(1145, 12), 125 => to_unsigned(1992, 12), 126 => to_unsigned(2969, 12), 127 => to_unsigned(2040, 12), 128 => to_unsigned(2334, 12), 129 => to_unsigned(3489, 12), 130 => to_unsigned(3308, 12), 131 => to_unsigned(1111, 12), 132 => to_unsigned(788, 12), 133 => to_unsigned(817, 12), 134 => to_unsigned(904, 12), 135 => to_unsigned(320, 12), 136 => to_unsigned(1954, 12), 137 => to_unsigned(1694, 12), 138 => to_unsigned(1894, 12), 139 => to_unsigned(3540, 12), 140 => to_unsigned(165, 12), 141 => to_unsigned(1814, 12), 142 => to_unsigned(2621, 12), 143 => to_unsigned(2346, 12), 144 => to_unsigned(1328, 12), 145 => to_unsigned(4054, 12), 146 => to_unsigned(105, 12), 147 => to_unsigned(2068, 12), 148 => to_unsigned(1963, 12), 149 => to_unsigned(3463, 12), 150 => to_unsigned(2753, 12), 151 => to_unsigned(1144, 12), 152 => to_unsigned(429, 12), 153 => to_unsigned(542, 12), 154 => to_unsigned(3724, 12), 155 => to_unsigned(1477, 12), 156 => to_unsigned(1848, 12), 157 => to_unsigned(2197, 12), 158 => to_unsigned(2245, 12), 159 => to_unsigned(3088, 12), 160 => to_unsigned(1579, 12), 161 => to_unsigned(1406, 12), 162 => to_unsigned(535, 12), 163 => to_unsigned(1192, 12), 164 => to_unsigned(4094, 12), 165 => to_unsigned(3493, 12), 166 => to_unsigned(1391, 12), 167 => to_unsigned(1968, 12), 168 => to_unsigned(2855, 12), 169 => to_unsigned(1640, 12), 170 => to_unsigned(2854, 12), 171 => to_unsigned(3499, 12), 172 => to_unsigned(3066, 12), 173 => to_unsigned(3760, 12), 174 => to_unsigned(2944, 12), 175 => to_unsigned(2185, 12), 176 => to_unsigned(764, 12), 177 => to_unsigned(1935, 12), 178 => to_unsigned(3508, 12), 179 => to_unsigned(1772, 12), 180 => to_unsigned(1077, 12), 181 => to_unsigned(766, 12), 182 => to_unsigned(2436, 12), 183 => to_unsigned(1692, 12), 184 => to_unsigned(3569, 12), 185 => to_unsigned(3107, 12), 186 => to_unsigned(3604, 12), 187 => to_unsigned(3334, 12), 188 => to_unsigned(1577, 12), 189 => to_unsigned(927, 12), 190 => to_unsigned(1241, 12), 191 => to_unsigned(2896, 12), 192 => to_unsigned(964, 12), 193 => to_unsigned(2286, 12), 194 => to_unsigned(3469, 12), 195 => to_unsigned(1953, 12), 196 => to_unsigned(1169, 12), 197 => to_unsigned(111, 12), 198 => to_unsigned(1601, 12), 199 => to_unsigned(601, 12), 200 => to_unsigned(1583, 12), 201 => to_unsigned(2390, 12), 202 => to_unsigned(554, 12), 203 => to_unsigned(2198, 12), 204 => to_unsigned(2001, 12), 205 => to_unsigned(1859, 12), 206 => to_unsigned(1171, 12), 207 => to_unsigned(2862, 12), 208 => to_unsigned(3357, 12), 209 => to_unsigned(758, 12), 210 => to_unsigned(1348, 12), 211 => to_unsigned(1492, 12), 212 => to_unsigned(365, 12), 213 => to_unsigned(2974, 12), 214 => to_unsigned(1708, 12), 215 => to_unsigned(1487, 12), 216 => to_unsigned(2977, 12), 217 => to_unsigned(4092, 12), 218 => to_unsigned(3844, 12), 219 => to_unsigned(2003, 12), 220 => to_unsigned(2981, 12), 221 => to_unsigned(2100, 12), 222 => to_unsigned(1344, 12), 223 => to_unsigned(1553, 12), 224 => to_unsigned(657, 12), 225 => to_unsigned(2033, 12), 226 => to_unsigned(1447, 12), 227 => to_unsigned(616, 12), 228 => to_unsigned(1298, 12), 229 => to_unsigned(3461, 12), 230 => to_unsigned(3938, 12), 231 => to_unsigned(3971, 12), 232 => to_unsigned(1338, 12), 233 => to_unsigned(3584, 12), 234 => to_unsigned(2679, 12), 235 => to_unsigned(2595, 12), 236 => to_unsigned(2329, 12), 237 => to_unsigned(2388, 12), 238 => to_unsigned(3677, 12), 239 => to_unsigned(449, 12), 240 => to_unsigned(3982, 12), 241 => to_unsigned(3628, 12), 242 => to_unsigned(742, 12), 243 => to_unsigned(260, 12), 244 => to_unsigned(3782, 12), 245 => to_unsigned(1681, 12), 246 => to_unsigned(2269, 12), 247 => to_unsigned(2493, 12), 248 => to_unsigned(1848, 12), 249 => to_unsigned(3969, 12), 250 => to_unsigned(2320, 12), 251 => to_unsigned(3266, 12), 252 => to_unsigned(2638, 12), 253 => to_unsigned(3434, 12), 254 => to_unsigned(689, 12), 255 => to_unsigned(24, 12), 256 => to_unsigned(2885, 12), 257 => to_unsigned(1913, 12), 258 => to_unsigned(405, 12), 259 => to_unsigned(1544, 12), 260 => to_unsigned(712, 12), 261 => to_unsigned(1313, 12), 262 => to_unsigned(69, 12), 263 => to_unsigned(1632, 12), 264 => to_unsigned(2037, 12), 265 => to_unsigned(256, 12), 266 => to_unsigned(811, 12), 267 => to_unsigned(2419, 12), 268 => to_unsigned(262, 12), 269 => to_unsigned(398, 12), 270 => to_unsigned(1189, 12), 271 => to_unsigned(1372, 12), 272 => to_unsigned(3536, 12), 273 => to_unsigned(309, 12), 274 => to_unsigned(1053, 12), 275 => to_unsigned(4084, 12), 276 => to_unsigned(4050, 12), 277 => to_unsigned(861, 12), 278 => to_unsigned(3704, 12), 279 => to_unsigned(2170, 12), 280 => to_unsigned(741, 12), 281 => to_unsigned(131, 12), 282 => to_unsigned(3050, 12), 283 => to_unsigned(3146, 12), 284 => to_unsigned(1321, 12), 285 => to_unsigned(3495, 12), 286 => to_unsigned(96, 12), 287 => to_unsigned(416, 12), 288 => to_unsigned(3228, 12), 289 => to_unsigned(2318, 12), 290 => to_unsigned(3551, 12), 291 => to_unsigned(2914, 12), 292 => to_unsigned(3902, 12), 293 => to_unsigned(1853, 12), 294 => to_unsigned(3429, 12), 295 => to_unsigned(1251, 12), 296 => to_unsigned(1859, 12), 297 => to_unsigned(2957, 12), 298 => to_unsigned(3986, 12), 299 => to_unsigned(2385, 12), 300 => to_unsigned(3389, 12), 301 => to_unsigned(3362, 12), 302 => to_unsigned(1634, 12), 303 => to_unsigned(2387, 12), 304 => to_unsigned(1522, 12), 305 => to_unsigned(452, 12), 306 => to_unsigned(2635, 12), 307 => to_unsigned(2965, 12), 308 => to_unsigned(2179, 12), 309 => to_unsigned(2161, 12), 310 => to_unsigned(34, 12), 311 => to_unsigned(2259, 12), 312 => to_unsigned(858, 12), 313 => to_unsigned(1736, 12), 314 => to_unsigned(2537, 12), 315 => to_unsigned(3534, 12), 316 => to_unsigned(2979, 12), 317 => to_unsigned(2764, 12), 318 => to_unsigned(3537, 12), 319 => to_unsigned(106, 12), 320 => to_unsigned(2007, 12), 321 => to_unsigned(465, 12), 322 => to_unsigned(1248, 12), 323 => to_unsigned(177, 12), 324 => to_unsigned(523, 12), 325 => to_unsigned(1640, 12), 326 => to_unsigned(322, 12), 327 => to_unsigned(3824, 12), 328 => to_unsigned(790, 12), 329 => to_unsigned(2244, 12), 330 => to_unsigned(3369, 12), 331 => to_unsigned(1834, 12), 332 => to_unsigned(911, 12), 333 => to_unsigned(2235, 12), 334 => to_unsigned(1340, 12), 335 => to_unsigned(3409, 12), 336 => to_unsigned(2919, 12), 337 => to_unsigned(205, 12), 338 => to_unsigned(3679, 12), 339 => to_unsigned(3939, 12), 340 => to_unsigned(2940, 12), 341 => to_unsigned(3953, 12), 342 => to_unsigned(1539, 12), 343 => to_unsigned(1530, 12), 344 => to_unsigned(941, 12), 345 => to_unsigned(3737, 12), 346 => to_unsigned(307, 12), 347 => to_unsigned(1948, 12), 348 => to_unsigned(2386, 12), 349 => to_unsigned(2156, 12), 350 => to_unsigned(2783, 12), 351 => to_unsigned(919, 12), 352 => to_unsigned(1646, 12), 353 => to_unsigned(3338, 12), 354 => to_unsigned(1933, 12), 355 => to_unsigned(3917, 12), 356 => to_unsigned(1549, 12), 357 => to_unsigned(2003, 12), 358 => to_unsigned(3905, 12), 359 => to_unsigned(3075, 12), 360 => to_unsigned(1164, 12), 361 => to_unsigned(3080, 12), 362 => to_unsigned(2035, 12), 363 => to_unsigned(3850, 12), 364 => to_unsigned(2941, 12), 365 => to_unsigned(774, 12), 366 => to_unsigned(2868, 12), 367 => to_unsigned(1439, 12), 368 => to_unsigned(887, 12), 369 => to_unsigned(3371, 12), 370 => to_unsigned(2015, 12), 371 => to_unsigned(661, 12), 372 => to_unsigned(269, 12), 373 => to_unsigned(3399, 12), 374 => to_unsigned(1325, 12), 375 => to_unsigned(540, 12), 376 => to_unsigned(1362, 12), 377 => to_unsigned(3997, 12), 378 => to_unsigned(1341, 12), 379 => to_unsigned(410, 12), 380 => to_unsigned(306, 12), 381 => to_unsigned(1551, 12), 382 => to_unsigned(4014, 12), 383 => to_unsigned(2881, 12), 384 => to_unsigned(1133, 12), 385 => to_unsigned(1715, 12), 386 => to_unsigned(2841, 12), 387 => to_unsigned(1554, 12), 388 => to_unsigned(3061, 12), 389 => to_unsigned(2599, 12), 390 => to_unsigned(3760, 12), 391 => to_unsigned(3885, 12), 392 => to_unsigned(918, 12), 393 => to_unsigned(539, 12), 394 => to_unsigned(3531, 12), 395 => to_unsigned(3116, 12), 396 => to_unsigned(2726, 12), 397 => to_unsigned(3313, 12), 398 => to_unsigned(2048, 12), 399 => to_unsigned(1673, 12), 400 => to_unsigned(534, 12), 401 => to_unsigned(3909, 12), 402 => to_unsigned(1661, 12), 403 => to_unsigned(1943, 12), 404 => to_unsigned(2886, 12), 405 => to_unsigned(3926, 12), 406 => to_unsigned(3031, 12), 407 => to_unsigned(3905, 12), 408 => to_unsigned(1975, 12), 409 => to_unsigned(2231, 12), 410 => to_unsigned(2970, 12), 411 => to_unsigned(671, 12), 412 => to_unsigned(1939, 12), 413 => to_unsigned(957, 12), 414 => to_unsigned(281, 12), 415 => to_unsigned(2024, 12), 416 => to_unsigned(2887, 12), 417 => to_unsigned(3595, 12), 418 => to_unsigned(2427, 12), 419 => to_unsigned(1209, 12), 420 => to_unsigned(567, 12), 421 => to_unsigned(2833, 12), 422 => to_unsigned(1974, 12), 423 => to_unsigned(1128, 12), 424 => to_unsigned(3328, 12), 425 => to_unsigned(1803, 12), 426 => to_unsigned(3620, 12), 427 => to_unsigned(2787, 12), 428 => to_unsigned(1229, 12), 429 => to_unsigned(2812, 12), 430 => to_unsigned(264, 12), 431 => to_unsigned(319, 12), 432 => to_unsigned(2022, 12), 433 => to_unsigned(3466, 12), 434 => to_unsigned(729, 12), 435 => to_unsigned(1769, 12), 436 => to_unsigned(1033, 12), 437 => to_unsigned(2678, 12), 438 => to_unsigned(84, 12), 439 => to_unsigned(260, 12), 440 => to_unsigned(443, 12), 441 => to_unsigned(3111, 12), 442 => to_unsigned(2768, 12), 443 => to_unsigned(2514, 12), 444 => to_unsigned(3822, 12), 445 => to_unsigned(2766, 12), 446 => to_unsigned(3287, 12), 447 => to_unsigned(2798, 12), 448 => to_unsigned(2356, 12), 449 => to_unsigned(2403, 12), 450 => to_unsigned(2171, 12), 451 => to_unsigned(560, 12), 452 => to_unsigned(1310, 12), 453 => to_unsigned(1027, 12), 454 => to_unsigned(2058, 12), 455 => to_unsigned(2336, 12), 456 => to_unsigned(1173, 12), 457 => to_unsigned(4009, 12), 458 => to_unsigned(2938, 12), 459 => to_unsigned(3182, 12), 460 => to_unsigned(1377, 12), 461 => to_unsigned(2706, 12), 462 => to_unsigned(225, 12), 463 => to_unsigned(3251, 12), 464 => to_unsigned(3276, 12), 465 => to_unsigned(1215, 12), 466 => to_unsigned(564, 12), 467 => to_unsigned(3522, 12), 468 => to_unsigned(1881, 12), 469 => to_unsigned(2538, 12), 470 => to_unsigned(2526, 12), 471 => to_unsigned(1715, 12), 472 => to_unsigned(2396, 12), 473 => to_unsigned(3241, 12), 474 => to_unsigned(2833, 12), 475 => to_unsigned(910, 12), 476 => to_unsigned(1851, 12), 477 => to_unsigned(3900, 12), 478 => to_unsigned(13, 12), 479 => to_unsigned(2657, 12), 480 => to_unsigned(3862, 12), 481 => to_unsigned(3316, 12), 482 => to_unsigned(3005, 12), 483 => to_unsigned(3416, 12), 484 => to_unsigned(2462, 12), 485 => to_unsigned(906, 12), 486 => to_unsigned(643, 12), 487 => to_unsigned(3231, 12), 488 => to_unsigned(1009, 12), 489 => to_unsigned(3104, 12), 490 => to_unsigned(3981, 12), 491 => to_unsigned(1201, 12), 492 => to_unsigned(3623, 12), 493 => to_unsigned(1408, 12), 494 => to_unsigned(1774, 12), 495 => to_unsigned(1560, 12), 496 => to_unsigned(340, 12), 497 => to_unsigned(555, 12), 498 => to_unsigned(2409, 12), 499 => to_unsigned(730, 12), 500 => to_unsigned(1243, 12), 501 => to_unsigned(3031, 12), 502 => to_unsigned(3162, 12), 503 => to_unsigned(1481, 12), 504 => to_unsigned(3937, 12), 505 => to_unsigned(1370, 12), 506 => to_unsigned(1449, 12), 507 => to_unsigned(3055, 12), 508 => to_unsigned(3231, 12), 509 => to_unsigned(3624, 12), 510 => to_unsigned(223, 12), 511 => to_unsigned(1288, 12), 512 => to_unsigned(433, 12), 513 => to_unsigned(3748, 12), 514 => to_unsigned(1361, 12), 515 => to_unsigned(862, 12), 516 => to_unsigned(3457, 12), 517 => to_unsigned(186, 12), 518 => to_unsigned(2333, 12), 519 => to_unsigned(245, 12), 520 => to_unsigned(1232, 12), 521 => to_unsigned(1108, 12), 522 => to_unsigned(1672, 12), 523 => to_unsigned(3703, 12), 524 => to_unsigned(2340, 12), 525 => to_unsigned(2909, 12), 526 => to_unsigned(1723, 12), 527 => to_unsigned(235, 12), 528 => to_unsigned(108, 12), 529 => to_unsigned(1295, 12), 530 => to_unsigned(2061, 12), 531 => to_unsigned(3737, 12), 532 => to_unsigned(1790, 12), 533 => to_unsigned(1253, 12), 534 => to_unsigned(1744, 12), 535 => to_unsigned(2866, 12), 536 => to_unsigned(3979, 12), 537 => to_unsigned(302, 12), 538 => to_unsigned(130, 12), 539 => to_unsigned(3233, 12), 540 => to_unsigned(476, 12), 541 => to_unsigned(602, 12), 542 => to_unsigned(3753, 12), 543 => to_unsigned(1281, 12), 544 => to_unsigned(1434, 12), 545 => to_unsigned(3528, 12), 546 => to_unsigned(339, 12), 547 => to_unsigned(411, 12), 548 => to_unsigned(3833, 12), 549 => to_unsigned(1635, 12), 550 => to_unsigned(3222, 12), 551 => to_unsigned(2777, 12), 552 => to_unsigned(3288, 12), 553 => to_unsigned(364, 12), 554 => to_unsigned(1876, 12), 555 => to_unsigned(1956, 12), 556 => to_unsigned(3317, 12), 557 => to_unsigned(2968, 12), 558 => to_unsigned(2590, 12), 559 => to_unsigned(1676, 12), 560 => to_unsigned(1844, 12), 561 => to_unsigned(3319, 12), 562 => to_unsigned(2794, 12), 563 => to_unsigned(1592, 12), 564 => to_unsigned(220, 12), 565 => to_unsigned(3826, 12), 566 => to_unsigned(68, 12), 567 => to_unsigned(4033, 12), 568 => to_unsigned(69, 12), 569 => to_unsigned(1196, 12), 570 => to_unsigned(1365, 12), 571 => to_unsigned(2810, 12), 572 => to_unsigned(1649, 12), 573 => to_unsigned(920, 12), 574 => to_unsigned(1160, 12), 575 => to_unsigned(1784, 12), 576 => to_unsigned(492, 12), 577 => to_unsigned(2170, 12), 578 => to_unsigned(3440, 12), 579 => to_unsigned(1402, 12), 580 => to_unsigned(414, 12), 581 => to_unsigned(288, 12), 582 => to_unsigned(1365, 12), 583 => to_unsigned(4035, 12), 584 => to_unsigned(2233, 12), 585 => to_unsigned(3957, 12), 586 => to_unsigned(3924, 12), 587 => to_unsigned(1361, 12), 588 => to_unsigned(3198, 12), 589 => to_unsigned(3217, 12), 590 => to_unsigned(3403, 12), 591 => to_unsigned(402, 12), 592 => to_unsigned(1913, 12), 593 => to_unsigned(2723, 12), 594 => to_unsigned(826, 12), 595 => to_unsigned(2645, 12), 596 => to_unsigned(2541, 12), 597 => to_unsigned(299, 12), 598 => to_unsigned(2495, 12), 599 => to_unsigned(3426, 12), 600 => to_unsigned(371, 12), 601 => to_unsigned(2145, 12), 602 => to_unsigned(969, 12), 603 => to_unsigned(2203, 12), 604 => to_unsigned(4055, 12), 605 => to_unsigned(4031, 12), 606 => to_unsigned(1001, 12), 607 => to_unsigned(1587, 12), 608 => to_unsigned(3643, 12), 609 => to_unsigned(1700, 12), 610 => to_unsigned(688, 12), 611 => to_unsigned(225, 12), 612 => to_unsigned(395, 12), 613 => to_unsigned(237, 12), 614 => to_unsigned(3656, 12), 615 => to_unsigned(1771, 12), 616 => to_unsigned(1518, 12), 617 => to_unsigned(3933, 12), 618 => to_unsigned(417, 12), 619 => to_unsigned(3759, 12), 620 => to_unsigned(2190, 12), 621 => to_unsigned(4062, 12), 622 => to_unsigned(1390, 12), 623 => to_unsigned(2719, 12), 624 => to_unsigned(1239, 12), 625 => to_unsigned(3903, 12), 626 => to_unsigned(1707, 12), 627 => to_unsigned(3605, 12), 628 => to_unsigned(1410, 12), 629 => to_unsigned(666, 12), 630 => to_unsigned(3300, 12), 631 => to_unsigned(2542, 12), 632 => to_unsigned(2057, 12), 633 => to_unsigned(2433, 12), 634 => to_unsigned(1976, 12), 635 => to_unsigned(835, 12), 636 => to_unsigned(849, 12), 637 => to_unsigned(3329, 12), 638 => to_unsigned(1136, 12), 639 => to_unsigned(2334, 12), 640 => to_unsigned(3618, 12), 641 => to_unsigned(993, 12), 642 => to_unsigned(2991, 12), 643 => to_unsigned(4016, 12), 644 => to_unsigned(2058, 12), 645 => to_unsigned(1273, 12), 646 => to_unsigned(3718, 12), 647 => to_unsigned(517, 12), 648 => to_unsigned(2346, 12), 649 => to_unsigned(198, 12), 650 => to_unsigned(3177, 12), 651 => to_unsigned(1702, 12), 652 => to_unsigned(2565, 12), 653 => to_unsigned(1340, 12), 654 => to_unsigned(2718, 12), 655 => to_unsigned(571, 12), 656 => to_unsigned(8, 12), 657 => to_unsigned(1215, 12), 658 => to_unsigned(3281, 12), 659 => to_unsigned(375, 12), 660 => to_unsigned(1622, 12), 661 => to_unsigned(2179, 12), 662 => to_unsigned(783, 12), 663 => to_unsigned(614, 12), 664 => to_unsigned(2414, 12), 665 => to_unsigned(2548, 12), 666 => to_unsigned(3934, 12), 667 => to_unsigned(6, 12), 668 => to_unsigned(1629, 12), 669 => to_unsigned(3094, 12), 670 => to_unsigned(2058, 12), 671 => to_unsigned(668, 12), 672 => to_unsigned(1927, 12), 673 => to_unsigned(1371, 12), 674 => to_unsigned(1520, 12), 675 => to_unsigned(1107, 12), 676 => to_unsigned(3586, 12), 677 => to_unsigned(2419, 12), 678 => to_unsigned(3399, 12), 679 => to_unsigned(1484, 12), 680 => to_unsigned(179, 12), 681 => to_unsigned(2323, 12), 682 => to_unsigned(2291, 12), 683 => to_unsigned(3678, 12), 684 => to_unsigned(1822, 12), 685 => to_unsigned(126, 12), 686 => to_unsigned(1307, 12), 687 => to_unsigned(1807, 12), 688 => to_unsigned(47, 12), 689 => to_unsigned(2583, 12), 690 => to_unsigned(954, 12), 691 => to_unsigned(862, 12), 692 => to_unsigned(2003, 12), 693 => to_unsigned(1160, 12), 694 => to_unsigned(1677, 12), 695 => to_unsigned(1318, 12), 696 => to_unsigned(678, 12), 697 => to_unsigned(2306, 12), 698 => to_unsigned(810, 12), 699 => to_unsigned(3123, 12), 700 => to_unsigned(2116, 12), 701 => to_unsigned(806, 12), 702 => to_unsigned(2757, 12), 703 => to_unsigned(3643, 12), 704 => to_unsigned(1983, 12), 705 => to_unsigned(437, 12), 706 => to_unsigned(1086, 12), 707 => to_unsigned(1390, 12), 708 => to_unsigned(1650, 12), 709 => to_unsigned(1441, 12), 710 => to_unsigned(88, 12), 711 => to_unsigned(2668, 12), 712 => to_unsigned(3292, 12), 713 => to_unsigned(3797, 12), 714 => to_unsigned(2301, 12), 715 => to_unsigned(2220, 12), 716 => to_unsigned(1678, 12), 717 => to_unsigned(3314, 12), 718 => to_unsigned(2420, 12), 719 => to_unsigned(2756, 12), 720 => to_unsigned(1385, 12), 721 => to_unsigned(2129, 12), 722 => to_unsigned(1743, 12), 723 => to_unsigned(3737, 12), 724 => to_unsigned(959, 12), 725 => to_unsigned(164, 12), 726 => to_unsigned(1420, 12), 727 => to_unsigned(550, 12), 728 => to_unsigned(3259, 12), 729 => to_unsigned(2525, 12), 730 => to_unsigned(3614, 12), 731 => to_unsigned(354, 12), 732 => to_unsigned(3539, 12), 733 => to_unsigned(3050, 12), 734 => to_unsigned(3923, 12), 735 => to_unsigned(1567, 12), 736 => to_unsigned(1001, 12), 737 => to_unsigned(868, 12), 738 => to_unsigned(3305, 12), 739 => to_unsigned(1867, 12), 740 => to_unsigned(2055, 12), 741 => to_unsigned(1093, 12), 742 => to_unsigned(333, 12), 743 => to_unsigned(1982, 12), 744 => to_unsigned(3554, 12), 745 => to_unsigned(430, 12), 746 => to_unsigned(1568, 12), 747 => to_unsigned(1056, 12), 748 => to_unsigned(1564, 12), 749 => to_unsigned(12, 12), 750 => to_unsigned(1117, 12), 751 => to_unsigned(3059, 12), 752 => to_unsigned(3146, 12), 753 => to_unsigned(3050, 12), 754 => to_unsigned(3127, 12), 755 => to_unsigned(2889, 12), 756 => to_unsigned(3059, 12), 757 => to_unsigned(2353, 12), 758 => to_unsigned(1531, 12), 759 => to_unsigned(1043, 12), 760 => to_unsigned(3286, 12), 761 => to_unsigned(2455, 12), 762 => to_unsigned(2590, 12), 763 => to_unsigned(956, 12), 764 => to_unsigned(436, 12), 765 => to_unsigned(3853, 12), 766 => to_unsigned(1522, 12), 767 => to_unsigned(1823, 12), 768 => to_unsigned(186, 12), 769 => to_unsigned(3324, 12), 770 => to_unsigned(1680, 12), 771 => to_unsigned(2834, 12), 772 => to_unsigned(3969, 12), 773 => to_unsigned(2063, 12), 774 => to_unsigned(1696, 12), 775 => to_unsigned(78, 12), 776 => to_unsigned(3913, 12), 777 => to_unsigned(774, 12), 778 => to_unsigned(3827, 12), 779 => to_unsigned(2927, 12), 780 => to_unsigned(2243, 12), 781 => to_unsigned(3142, 12), 782 => to_unsigned(3958, 12), 783 => to_unsigned(3279, 12), 784 => to_unsigned(3805, 12), 785 => to_unsigned(1877, 12), 786 => to_unsigned(3251, 12), 787 => to_unsigned(3914, 12), 788 => to_unsigned(2234, 12), 789 => to_unsigned(973, 12), 790 => to_unsigned(859, 12), 791 => to_unsigned(2970, 12), 792 => to_unsigned(1562, 12), 793 => to_unsigned(3817, 12), 794 => to_unsigned(2628, 12), 795 => to_unsigned(3899, 12), 796 => to_unsigned(925, 12), 797 => to_unsigned(3760, 12), 798 => to_unsigned(2396, 12), 799 => to_unsigned(3389, 12), 800 => to_unsigned(3772, 12), 801 => to_unsigned(3983, 12), 802 => to_unsigned(3950, 12), 803 => to_unsigned(505, 12), 804 => to_unsigned(91, 12), 805 => to_unsigned(3496, 12), 806 => to_unsigned(2208, 12), 807 => to_unsigned(2733, 12), 808 => to_unsigned(113, 12), 809 => to_unsigned(398, 12), 810 => to_unsigned(2884, 12), 811 => to_unsigned(2393, 12), 812 => to_unsigned(1504, 12), 813 => to_unsigned(3340, 12), 814 => to_unsigned(3756, 12), 815 => to_unsigned(3945, 12), 816 => to_unsigned(1339, 12), 817 => to_unsigned(1450, 12), 818 => to_unsigned(3007, 12), 819 => to_unsigned(820, 12), 820 => to_unsigned(3469, 12), 821 => to_unsigned(2484, 12), 822 => to_unsigned(1202, 12), 823 => to_unsigned(120, 12), 824 => to_unsigned(946, 12), 825 => to_unsigned(1905, 12), 826 => to_unsigned(4037, 12), 827 => to_unsigned(2519, 12), 828 => to_unsigned(2789, 12), 829 => to_unsigned(3700, 12), 830 => to_unsigned(3038, 12), 831 => to_unsigned(3548, 12), 832 => to_unsigned(1206, 12), 833 => to_unsigned(3029, 12), 834 => to_unsigned(1875, 12), 835 => to_unsigned(2904, 12), 836 => to_unsigned(2425, 12), 837 => to_unsigned(1711, 12), 838 => to_unsigned(599, 12), 839 => to_unsigned(2989, 12), 840 => to_unsigned(3134, 12), 841 => to_unsigned(2314, 12), 842 => to_unsigned(2654, 12), 843 => to_unsigned(1120, 12), 844 => to_unsigned(2005, 12), 845 => to_unsigned(2920, 12), 846 => to_unsigned(1078, 12), 847 => to_unsigned(862, 12), 848 => to_unsigned(1670, 12), 849 => to_unsigned(1945, 12), 850 => to_unsigned(2565, 12), 851 => to_unsigned(695, 12), 852 => to_unsigned(3807, 12), 853 => to_unsigned(3119, 12), 854 => to_unsigned(1518, 12), 855 => to_unsigned(411, 12), 856 => to_unsigned(3417, 12), 857 => to_unsigned(2465, 12), 858 => to_unsigned(731, 12), 859 => to_unsigned(3984, 12), 860 => to_unsigned(1680, 12), 861 => to_unsigned(2383, 12), 862 => to_unsigned(3806, 12), 863 => to_unsigned(3490, 12), 864 => to_unsigned(2491, 12), 865 => to_unsigned(3141, 12), 866 => to_unsigned(3144, 12), 867 => to_unsigned(1680, 12), 868 => to_unsigned(2278, 12), 869 => to_unsigned(1843, 12), 870 => to_unsigned(3559, 12), 871 => to_unsigned(1628, 12), 872 => to_unsigned(3717, 12), 873 => to_unsigned(0, 12), 874 => to_unsigned(723, 12), 875 => to_unsigned(535, 12), 876 => to_unsigned(1532, 12), 877 => to_unsigned(3230, 12), 878 => to_unsigned(756, 12), 879 => to_unsigned(622, 12), 880 => to_unsigned(806, 12), 881 => to_unsigned(2728, 12), 882 => to_unsigned(738, 12), 883 => to_unsigned(1617, 12), 884 => to_unsigned(2687, 12), 885 => to_unsigned(911, 12), 886 => to_unsigned(2122, 12), 887 => to_unsigned(3346, 12), 888 => to_unsigned(1512, 12), 889 => to_unsigned(1307, 12), 890 => to_unsigned(2355, 12), 891 => to_unsigned(892, 12), 892 => to_unsigned(426, 12), 893 => to_unsigned(1510, 12), 894 => to_unsigned(718, 12), 895 => to_unsigned(1839, 12), 896 => to_unsigned(3409, 12), 897 => to_unsigned(252, 12), 898 => to_unsigned(3447, 12), 899 => to_unsigned(3241, 12), 900 => to_unsigned(236, 12), 901 => to_unsigned(899, 12), 902 => to_unsigned(3568, 12), 903 => to_unsigned(3189, 12), 904 => to_unsigned(1945, 12), 905 => to_unsigned(216, 12), 906 => to_unsigned(2924, 12), 907 => to_unsigned(991, 12), 908 => to_unsigned(3287, 12), 909 => to_unsigned(2045, 12), 910 => to_unsigned(2383, 12), 911 => to_unsigned(2069, 12), 912 => to_unsigned(3132, 12), 913 => to_unsigned(3101, 12), 914 => to_unsigned(2582, 12), 915 => to_unsigned(24, 12), 916 => to_unsigned(2115, 12), 917 => to_unsigned(1673, 12), 918 => to_unsigned(550, 12), 919 => to_unsigned(1856, 12), 920 => to_unsigned(2383, 12), 921 => to_unsigned(492, 12), 922 => to_unsigned(3049, 12), 923 => to_unsigned(142, 12), 924 => to_unsigned(2629, 12), 925 => to_unsigned(3153, 12), 926 => to_unsigned(698, 12), 927 => to_unsigned(361, 12), 928 => to_unsigned(579, 12), 929 => to_unsigned(240, 12), 930 => to_unsigned(2259, 12), 931 => to_unsigned(2130, 12), 932 => to_unsigned(363, 12), 933 => to_unsigned(689, 12), 934 => to_unsigned(1649, 12), 935 => to_unsigned(385, 12), 936 => to_unsigned(1671, 12), 937 => to_unsigned(520, 12), 938 => to_unsigned(3615, 12), 939 => to_unsigned(636, 12), 940 => to_unsigned(3342, 12), 941 => to_unsigned(206, 12), 942 => to_unsigned(3476, 12), 943 => to_unsigned(2194, 12), 944 => to_unsigned(1775, 12), 945 => to_unsigned(1187, 12), 946 => to_unsigned(812, 12), 947 => to_unsigned(1000, 12), 948 => to_unsigned(2407, 12), 949 => to_unsigned(1695, 12), 950 => to_unsigned(3265, 12), 951 => to_unsigned(2778, 12), 952 => to_unsigned(3321, 12), 953 => to_unsigned(2456, 12), 954 => to_unsigned(1318, 12), 955 => to_unsigned(41, 12), 956 => to_unsigned(2783, 12), 957 => to_unsigned(1208, 12), 958 => to_unsigned(2635, 12), 959 => to_unsigned(2544, 12), 960 => to_unsigned(2619, 12), 961 => to_unsigned(3875, 12), 962 => to_unsigned(331, 12), 963 => to_unsigned(2801, 12), 964 => to_unsigned(3631, 12), 965 => to_unsigned(1457, 12), 966 => to_unsigned(2801, 12), 967 => to_unsigned(3442, 12), 968 => to_unsigned(2287, 12), 969 => to_unsigned(1906, 12), 970 => to_unsigned(1389, 12), 971 => to_unsigned(2333, 12), 972 => to_unsigned(996, 12), 973 => to_unsigned(818, 12), 974 => to_unsigned(2169, 12), 975 => to_unsigned(2954, 12), 976 => to_unsigned(554, 12), 977 => to_unsigned(3610, 12), 978 => to_unsigned(1020, 12), 979 => to_unsigned(1227, 12), 980 => to_unsigned(697, 12), 981 => to_unsigned(1129, 12), 982 => to_unsigned(3527, 12), 983 => to_unsigned(2941, 12), 984 => to_unsigned(372, 12), 985 => to_unsigned(1760, 12), 986 => to_unsigned(3291, 12), 987 => to_unsigned(2311, 12), 988 => to_unsigned(439, 12), 989 => to_unsigned(3284, 12), 990 => to_unsigned(401, 12), 991 => to_unsigned(74, 12), 992 => to_unsigned(988, 12), 993 => to_unsigned(710, 12), 994 => to_unsigned(1592, 12), 995 => to_unsigned(2460, 12), 996 => to_unsigned(2303, 12), 997 => to_unsigned(1680, 12), 998 => to_unsigned(61, 12), 999 => to_unsigned(1860, 12), 1000 => to_unsigned(2245, 12), 1001 => to_unsigned(472, 12), 1002 => to_unsigned(3756, 12), 1003 => to_unsigned(2358, 12), 1004 => to_unsigned(1008, 12), 1005 => to_unsigned(1952, 12), 1006 => to_unsigned(3694, 12), 1007 => to_unsigned(3788, 12), 1008 => to_unsigned(2487, 12), 1009 => to_unsigned(1473, 12), 1010 => to_unsigned(751, 12), 1011 => to_unsigned(2316, 12), 1012 => to_unsigned(1433, 12), 1013 => to_unsigned(1600, 12), 1014 => to_unsigned(2373, 12), 1015 => to_unsigned(76, 12), 1016 => to_unsigned(926, 12), 1017 => to_unsigned(680, 12), 1018 => to_unsigned(3985, 12), 1019 => to_unsigned(3484, 12), 1020 => to_unsigned(500, 12), 1021 => to_unsigned(2332, 12), 1022 => to_unsigned(11, 12), 1023 => to_unsigned(2653, 12), 1024 => to_unsigned(1601, 12), 1025 => to_unsigned(3176, 12), 1026 => to_unsigned(1408, 12), 1027 => to_unsigned(108, 12), 1028 => to_unsigned(690, 12), 1029 => to_unsigned(762, 12), 1030 => to_unsigned(2459, 12), 1031 => to_unsigned(2232, 12), 1032 => to_unsigned(3068, 12), 1033 => to_unsigned(2127, 12), 1034 => to_unsigned(875, 12), 1035 => to_unsigned(3764, 12), 1036 => to_unsigned(2320, 12), 1037 => to_unsigned(346, 12), 1038 => to_unsigned(589, 12), 1039 => to_unsigned(3609, 12), 1040 => to_unsigned(3049, 12), 1041 => to_unsigned(919, 12), 1042 => to_unsigned(2364, 12), 1043 => to_unsigned(3015, 12), 1044 => to_unsigned(3475, 12), 1045 => to_unsigned(2534, 12), 1046 => to_unsigned(1601, 12), 1047 => to_unsigned(2155, 12), 1048 => to_unsigned(2494, 12), 1049 => to_unsigned(2216, 12), 1050 => to_unsigned(324, 12), 1051 => to_unsigned(2191, 12), 1052 => to_unsigned(21, 12), 1053 => to_unsigned(275, 12), 1054 => to_unsigned(3740, 12), 1055 => to_unsigned(3809, 12), 1056 => to_unsigned(650, 12), 1057 => to_unsigned(1048, 12), 1058 => to_unsigned(153, 12), 1059 => to_unsigned(1205, 12), 1060 => to_unsigned(3591, 12), 1061 => to_unsigned(1428, 12), 1062 => to_unsigned(1891, 12), 1063 => to_unsigned(1239, 12), 1064 => to_unsigned(2750, 12), 1065 => to_unsigned(2494, 12), 1066 => to_unsigned(3022, 12), 1067 => to_unsigned(3215, 12), 1068 => to_unsigned(1668, 12), 1069 => to_unsigned(1387, 12), 1070 => to_unsigned(1636, 12), 1071 => to_unsigned(3294, 12), 1072 => to_unsigned(1120, 12), 1073 => to_unsigned(871, 12), 1074 => to_unsigned(490, 12), 1075 => to_unsigned(2645, 12), 1076 => to_unsigned(2675, 12), 1077 => to_unsigned(2945, 12), 1078 => to_unsigned(690, 12), 1079 => to_unsigned(3095, 12), 1080 => to_unsigned(3136, 12), 1081 => to_unsigned(270, 12), 1082 => to_unsigned(475, 12), 1083 => to_unsigned(3572, 12), 1084 => to_unsigned(1229, 12), 1085 => to_unsigned(3365, 12), 1086 => to_unsigned(2612, 12), 1087 => to_unsigned(3426, 12), 1088 => to_unsigned(716, 12), 1089 => to_unsigned(1410, 12), 1090 => to_unsigned(114, 12), 1091 => to_unsigned(2401, 12), 1092 => to_unsigned(1527, 12), 1093 => to_unsigned(1230, 12), 1094 => to_unsigned(2961, 12), 1095 => to_unsigned(2025, 12), 1096 => to_unsigned(3372, 12), 1097 => to_unsigned(1735, 12), 1098 => to_unsigned(3099, 12), 1099 => to_unsigned(1431, 12), 1100 => to_unsigned(3171, 12), 1101 => to_unsigned(751, 12), 1102 => to_unsigned(577, 12), 1103 => to_unsigned(3143, 12), 1104 => to_unsigned(2105, 12), 1105 => to_unsigned(1527, 12), 1106 => to_unsigned(2891, 12), 1107 => to_unsigned(2233, 12), 1108 => to_unsigned(231, 12), 1109 => to_unsigned(266, 12), 1110 => to_unsigned(2056, 12), 1111 => to_unsigned(2830, 12), 1112 => to_unsigned(2013, 12), 1113 => to_unsigned(607, 12), 1114 => to_unsigned(1818, 12), 1115 => to_unsigned(1843, 12), 1116 => to_unsigned(425, 12), 1117 => to_unsigned(976, 12), 1118 => to_unsigned(3113, 12), 1119 => to_unsigned(2807, 12), 1120 => to_unsigned(2301, 12), 1121 => to_unsigned(813, 12), 1122 => to_unsigned(2399, 12), 1123 => to_unsigned(666, 12), 1124 => to_unsigned(3829, 12), 1125 => to_unsigned(3173, 12), 1126 => to_unsigned(2815, 12), 1127 => to_unsigned(3013, 12), 1128 => to_unsigned(589, 12), 1129 => to_unsigned(2825, 12), 1130 => to_unsigned(3349, 12), 1131 => to_unsigned(2, 12), 1132 => to_unsigned(2287, 12), 1133 => to_unsigned(416, 12), 1134 => to_unsigned(1604, 12), 1135 => to_unsigned(124, 12), 1136 => to_unsigned(1960, 12), 1137 => to_unsigned(2822, 12), 1138 => to_unsigned(193, 12), 1139 => to_unsigned(309, 12), 1140 => to_unsigned(3446, 12), 1141 => to_unsigned(2407, 12), 1142 => to_unsigned(3124, 12), 1143 => to_unsigned(1598, 12), 1144 => to_unsigned(3306, 12), 1145 => to_unsigned(1855, 12), 1146 => to_unsigned(3447, 12), 1147 => to_unsigned(3276, 12), 1148 => to_unsigned(826, 12), 1149 => to_unsigned(3501, 12), 1150 => to_unsigned(3926, 12), 1151 => to_unsigned(1000, 12), 1152 => to_unsigned(1612, 12), 1153 => to_unsigned(1296, 12), 1154 => to_unsigned(3395, 12), 1155 => to_unsigned(3286, 12), 1156 => to_unsigned(767, 12), 1157 => to_unsigned(1816, 12), 1158 => to_unsigned(2181, 12), 1159 => to_unsigned(3796, 12), 1160 => to_unsigned(765, 12), 1161 => to_unsigned(1802, 12), 1162 => to_unsigned(1128, 12), 1163 => to_unsigned(1212, 12), 1164 => to_unsigned(345, 12), 1165 => to_unsigned(3098, 12), 1166 => to_unsigned(1689, 12), 1167 => to_unsigned(1246, 12), 1168 => to_unsigned(2329, 12), 1169 => to_unsigned(2629, 12), 1170 => to_unsigned(3355, 12), 1171 => to_unsigned(1216, 12), 1172 => to_unsigned(3873, 12), 1173 => to_unsigned(1794, 12), 1174 => to_unsigned(1481, 12), 1175 => to_unsigned(2254, 12), 1176 => to_unsigned(3517, 12), 1177 => to_unsigned(3879, 12), 1178 => to_unsigned(1431, 12), 1179 => to_unsigned(2027, 12), 1180 => to_unsigned(2484, 12), 1181 => to_unsigned(1221, 12), 1182 => to_unsigned(34, 12), 1183 => to_unsigned(1503, 12), 1184 => to_unsigned(1922, 12), 1185 => to_unsigned(1380, 12), 1186 => to_unsigned(3790, 12), 1187 => to_unsigned(2843, 12), 1188 => to_unsigned(667, 12), 1189 => to_unsigned(2240, 12), 1190 => to_unsigned(3413, 12), 1191 => to_unsigned(2026, 12), 1192 => to_unsigned(1272, 12), 1193 => to_unsigned(2789, 12), 1194 => to_unsigned(3857, 12), 1195 => to_unsigned(840, 12), 1196 => to_unsigned(3208, 12), 1197 => to_unsigned(813, 12), 1198 => to_unsigned(2829, 12), 1199 => to_unsigned(1556, 12), 1200 => to_unsigned(3696, 12), 1201 => to_unsigned(3477, 12), 1202 => to_unsigned(3415, 12), 1203 => to_unsigned(129, 12), 1204 => to_unsigned(1958, 12), 1205 => to_unsigned(750, 12), 1206 => to_unsigned(824, 12), 1207 => to_unsigned(2635, 12), 1208 => to_unsigned(664, 12), 1209 => to_unsigned(2039, 12), 1210 => to_unsigned(2909, 12), 1211 => to_unsigned(1439, 12), 1212 => to_unsigned(1685, 12), 1213 => to_unsigned(1756, 12), 1214 => to_unsigned(2764, 12), 1215 => to_unsigned(3804, 12), 1216 => to_unsigned(3560, 12), 1217 => to_unsigned(2369, 12), 1218 => to_unsigned(2655, 12), 1219 => to_unsigned(1974, 12), 1220 => to_unsigned(650, 12), 1221 => to_unsigned(2780, 12), 1222 => to_unsigned(2096, 12), 1223 => to_unsigned(3946, 12), 1224 => to_unsigned(3045, 12), 1225 => to_unsigned(2837, 12), 1226 => to_unsigned(1739, 12), 1227 => to_unsigned(3571, 12), 1228 => to_unsigned(132, 12), 1229 => to_unsigned(2044, 12), 1230 => to_unsigned(486, 12), 1231 => to_unsigned(3195, 12), 1232 => to_unsigned(2156, 12), 1233 => to_unsigned(1230, 12), 1234 => to_unsigned(2485, 12), 1235 => to_unsigned(2531, 12), 1236 => to_unsigned(3576, 12), 1237 => to_unsigned(3767, 12), 1238 => to_unsigned(999, 12), 1239 => to_unsigned(426, 12), 1240 => to_unsigned(1784, 12), 1241 => to_unsigned(2655, 12), 1242 => to_unsigned(3627, 12), 1243 => to_unsigned(1352, 12), 1244 => to_unsigned(1787, 12), 1245 => to_unsigned(918, 12), 1246 => to_unsigned(2599, 12), 1247 => to_unsigned(4008, 12), 1248 => to_unsigned(34, 12), 1249 => to_unsigned(291, 12), 1250 => to_unsigned(2548, 12), 1251 => to_unsigned(996, 12), 1252 => to_unsigned(1460, 12), 1253 => to_unsigned(223, 12), 1254 => to_unsigned(2814, 12), 1255 => to_unsigned(1723, 12), 1256 => to_unsigned(3492, 12), 1257 => to_unsigned(2609, 12), 1258 => to_unsigned(530, 12), 1259 => to_unsigned(3509, 12), 1260 => to_unsigned(3469, 12), 1261 => to_unsigned(2358, 12), 1262 => to_unsigned(246, 12), 1263 => to_unsigned(191, 12), 1264 => to_unsigned(1721, 12), 1265 => to_unsigned(1071, 12), 1266 => to_unsigned(3979, 12), 1267 => to_unsigned(2795, 12), 1268 => to_unsigned(2290, 12), 1269 => to_unsigned(2005, 12), 1270 => to_unsigned(1728, 12), 1271 => to_unsigned(2942, 12), 1272 => to_unsigned(2682, 12), 1273 => to_unsigned(1705, 12), 1274 => to_unsigned(2705, 12), 1275 => to_unsigned(3217, 12), 1276 => to_unsigned(3837, 12), 1277 => to_unsigned(2465, 12), 1278 => to_unsigned(3112, 12), 1279 => to_unsigned(227, 12), 1280 => to_unsigned(419, 12), 1281 => to_unsigned(3362, 12), 1282 => to_unsigned(2907, 12), 1283 => to_unsigned(2531, 12), 1284 => to_unsigned(3187, 12), 1285 => to_unsigned(3616, 12), 1286 => to_unsigned(3736, 12), 1287 => to_unsigned(3707, 12), 1288 => to_unsigned(2057, 12), 1289 => to_unsigned(2651, 12), 1290 => to_unsigned(4013, 12), 1291 => to_unsigned(2970, 12), 1292 => to_unsigned(1549, 12), 1293 => to_unsigned(1188, 12), 1294 => to_unsigned(3370, 12), 1295 => to_unsigned(3836, 12), 1296 => to_unsigned(1304, 12), 1297 => to_unsigned(816, 12), 1298 => to_unsigned(1331, 12), 1299 => to_unsigned(988, 12), 1300 => to_unsigned(3568, 12), 1301 => to_unsigned(504, 12), 1302 => to_unsigned(3555, 12), 1303 => to_unsigned(2207, 12), 1304 => to_unsigned(672, 12), 1305 => to_unsigned(1196, 12), 1306 => to_unsigned(2650, 12), 1307 => to_unsigned(3208, 12), 1308 => to_unsigned(1041, 12), 1309 => to_unsigned(1647, 12), 1310 => to_unsigned(2710, 12), 1311 => to_unsigned(413, 12), 1312 => to_unsigned(1792, 12), 1313 => to_unsigned(3566, 12), 1314 => to_unsigned(2566, 12), 1315 => to_unsigned(207, 12), 1316 => to_unsigned(149, 12), 1317 => to_unsigned(594, 12), 1318 => to_unsigned(3011, 12), 1319 => to_unsigned(3189, 12), 1320 => to_unsigned(3187, 12), 1321 => to_unsigned(2583, 12), 1322 => to_unsigned(2362, 12), 1323 => to_unsigned(2187, 12), 1324 => to_unsigned(3126, 12), 1325 => to_unsigned(3392, 12), 1326 => to_unsigned(228, 12), 1327 => to_unsigned(1048, 12), 1328 => to_unsigned(4036, 12), 1329 => to_unsigned(3113, 12), 1330 => to_unsigned(290, 12), 1331 => to_unsigned(2242, 12), 1332 => to_unsigned(2184, 12), 1333 => to_unsigned(2979, 12), 1334 => to_unsigned(4074, 12), 1335 => to_unsigned(644, 12), 1336 => to_unsigned(195, 12), 1337 => to_unsigned(2468, 12), 1338 => to_unsigned(1602, 12), 1339 => to_unsigned(2956, 12), 1340 => to_unsigned(2879, 12), 1341 => to_unsigned(2393, 12), 1342 => to_unsigned(1660, 12), 1343 => to_unsigned(1816, 12), 1344 => to_unsigned(3617, 12), 1345 => to_unsigned(1967, 12), 1346 => to_unsigned(2480, 12), 1347 => to_unsigned(300, 12), 1348 => to_unsigned(2019, 12), 1349 => to_unsigned(824, 12), 1350 => to_unsigned(739, 12), 1351 => to_unsigned(2441, 12), 1352 => to_unsigned(175, 12), 1353 => to_unsigned(900, 12), 1354 => to_unsigned(3403, 12), 1355 => to_unsigned(1384, 12), 1356 => to_unsigned(1050, 12), 1357 => to_unsigned(777, 12), 1358 => to_unsigned(1881, 12), 1359 => to_unsigned(123, 12), 1360 => to_unsigned(1865, 12), 1361 => to_unsigned(3484, 12), 1362 => to_unsigned(89, 12), 1363 => to_unsigned(3821, 12), 1364 => to_unsigned(2372, 12), 1365 => to_unsigned(542, 12), 1366 => to_unsigned(3631, 12), 1367 => to_unsigned(1441, 12), 1368 => to_unsigned(117, 12), 1369 => to_unsigned(3677, 12), 1370 => to_unsigned(1757, 12), 1371 => to_unsigned(3540, 12), 1372 => to_unsigned(2357, 12), 1373 => to_unsigned(2808, 12), 1374 => to_unsigned(3831, 12), 1375 => to_unsigned(336, 12), 1376 => to_unsigned(2911, 12), 1377 => to_unsigned(3494, 12), 1378 => to_unsigned(193, 12), 1379 => to_unsigned(1345, 12), 1380 => to_unsigned(1517, 12), 1381 => to_unsigned(1694, 12), 1382 => to_unsigned(2857, 12), 1383 => to_unsigned(2047, 12), 1384 => to_unsigned(4084, 12), 1385 => to_unsigned(2213, 12), 1386 => to_unsigned(2346, 12), 1387 => to_unsigned(3585, 12), 1388 => to_unsigned(702, 12), 1389 => to_unsigned(5, 12), 1390 => to_unsigned(654, 12), 1391 => to_unsigned(2185, 12), 1392 => to_unsigned(2005, 12), 1393 => to_unsigned(3651, 12), 1394 => to_unsigned(2078, 12), 1395 => to_unsigned(1687, 12), 1396 => to_unsigned(337, 12), 1397 => to_unsigned(138, 12), 1398 => to_unsigned(559, 12), 1399 => to_unsigned(1021, 12), 1400 => to_unsigned(1463, 12), 1401 => to_unsigned(688, 12), 1402 => to_unsigned(2438, 12), 1403 => to_unsigned(3398, 12), 1404 => to_unsigned(2069, 12), 1405 => to_unsigned(2467, 12), 1406 => to_unsigned(2283, 12), 1407 => to_unsigned(1307, 12), 1408 => to_unsigned(912, 12), 1409 => to_unsigned(1830, 12), 1410 => to_unsigned(1188, 12), 1411 => to_unsigned(3335, 12), 1412 => to_unsigned(1038, 12), 1413 => to_unsigned(549, 12), 1414 => to_unsigned(1988, 12), 1415 => to_unsigned(287, 12), 1416 => to_unsigned(584, 12), 1417 => to_unsigned(419, 12), 1418 => to_unsigned(327, 12), 1419 => to_unsigned(87, 12), 1420 => to_unsigned(314, 12), 1421 => to_unsigned(1976, 12), 1422 => to_unsigned(3651, 12), 1423 => to_unsigned(875, 12), 1424 => to_unsigned(1489, 12), 1425 => to_unsigned(872, 12), 1426 => to_unsigned(892, 12), 1427 => to_unsigned(309, 12), 1428 => to_unsigned(3995, 12), 1429 => to_unsigned(2340, 12), 1430 => to_unsigned(4068, 12), 1431 => to_unsigned(3281, 12), 1432 => to_unsigned(1697, 12), 1433 => to_unsigned(936, 12), 1434 => to_unsigned(2413, 12), 1435 => to_unsigned(1448, 12), 1436 => to_unsigned(723, 12), 1437 => to_unsigned(287, 12), 1438 => to_unsigned(1906, 12), 1439 => to_unsigned(3670, 12), 1440 => to_unsigned(515, 12), 1441 => to_unsigned(3436, 12), 1442 => to_unsigned(512, 12), 1443 => to_unsigned(2848, 12), 1444 => to_unsigned(1925, 12), 1445 => to_unsigned(232, 12), 1446 => to_unsigned(2823, 12), 1447 => to_unsigned(2245, 12), 1448 => to_unsigned(2191, 12), 1449 => to_unsigned(621, 12), 1450 => to_unsigned(984, 12), 1451 => to_unsigned(3818, 12), 1452 => to_unsigned(3659, 12), 1453 => to_unsigned(960, 12), 1454 => to_unsigned(2298, 12), 1455 => to_unsigned(1313, 12), 1456 => to_unsigned(418, 12), 1457 => to_unsigned(2592, 12), 1458 => to_unsigned(3390, 12), 1459 => to_unsigned(1838, 12), 1460 => to_unsigned(184, 12), 1461 => to_unsigned(3394, 12), 1462 => to_unsigned(312, 12), 1463 => to_unsigned(2079, 12), 1464 => to_unsigned(1616, 12), 1465 => to_unsigned(198, 12), 1466 => to_unsigned(1546, 12), 1467 => to_unsigned(1814, 12), 1468 => to_unsigned(2230, 12), 1469 => to_unsigned(2190, 12), 1470 => to_unsigned(163, 12), 1471 => to_unsigned(180, 12), 1472 => to_unsigned(2627, 12), 1473 => to_unsigned(1642, 12), 1474 => to_unsigned(3888, 12), 1475 => to_unsigned(435, 12), 1476 => to_unsigned(3302, 12), 1477 => to_unsigned(2922, 12), 1478 => to_unsigned(2618, 12), 1479 => to_unsigned(470, 12), 1480 => to_unsigned(3245, 12), 1481 => to_unsigned(557, 12), 1482 => to_unsigned(758, 12), 1483 => to_unsigned(741, 12), 1484 => to_unsigned(1913, 12), 1485 => to_unsigned(464, 12), 1486 => to_unsigned(1889, 12), 1487 => to_unsigned(1684, 12), 1488 => to_unsigned(510, 12), 1489 => to_unsigned(1959, 12), 1490 => to_unsigned(3682, 12), 1491 => to_unsigned(2218, 12), 1492 => to_unsigned(1469, 12), 1493 => to_unsigned(2870, 12), 1494 => to_unsigned(2912, 12), 1495 => to_unsigned(1633, 12), 1496 => to_unsigned(1521, 12), 1497 => to_unsigned(1840, 12), 1498 => to_unsigned(689, 12), 1499 => to_unsigned(991, 12), 1500 => to_unsigned(2389, 12), 1501 => to_unsigned(3200, 12), 1502 => to_unsigned(2582, 12), 1503 => to_unsigned(2623, 12), 1504 => to_unsigned(2897, 12), 1505 => to_unsigned(4032, 12), 1506 => to_unsigned(1317, 12), 1507 => to_unsigned(3708, 12), 1508 => to_unsigned(557, 12), 1509 => to_unsigned(502, 12), 1510 => to_unsigned(2095, 12), 1511 => to_unsigned(1032, 12), 1512 => to_unsigned(2038, 12), 1513 => to_unsigned(432, 12), 1514 => to_unsigned(2089, 12), 1515 => to_unsigned(2977, 12), 1516 => to_unsigned(3319, 12), 1517 => to_unsigned(85, 12), 1518 => to_unsigned(3173, 12), 1519 => to_unsigned(1632, 12), 1520 => to_unsigned(3536, 12), 1521 => to_unsigned(17, 12), 1522 => to_unsigned(2586, 12), 1523 => to_unsigned(3845, 12), 1524 => to_unsigned(939, 12), 1525 => to_unsigned(2966, 12), 1526 => to_unsigned(1732, 12), 1527 => to_unsigned(1336, 12), 1528 => to_unsigned(1609, 12), 1529 => to_unsigned(3285, 12), 1530 => to_unsigned(2859, 12), 1531 => to_unsigned(917, 12), 1532 => to_unsigned(1343, 12), 1533 => to_unsigned(3000, 12), 1534 => to_unsigned(2713, 12), 1535 => to_unsigned(1935, 12), 1536 => to_unsigned(1953, 12), 1537 => to_unsigned(3186, 12), 1538 => to_unsigned(1496, 12), 1539 => to_unsigned(1221, 12), 1540 => to_unsigned(3390, 12), 1541 => to_unsigned(710, 12), 1542 => to_unsigned(695, 12), 1543 => to_unsigned(1165, 12), 1544 => to_unsigned(2011, 12), 1545 => to_unsigned(1292, 12), 1546 => to_unsigned(1154, 12), 1547 => to_unsigned(2644, 12), 1548 => to_unsigned(3134, 12), 1549 => to_unsigned(3830, 12), 1550 => to_unsigned(768, 12), 1551 => to_unsigned(2067, 12), 1552 => to_unsigned(2723, 12), 1553 => to_unsigned(2902, 12), 1554 => to_unsigned(1555, 12), 1555 => to_unsigned(761, 12), 1556 => to_unsigned(1659, 12), 1557 => to_unsigned(385, 12), 1558 => to_unsigned(3614, 12), 1559 => to_unsigned(1527, 12), 1560 => to_unsigned(1773, 12), 1561 => to_unsigned(2019, 12), 1562 => to_unsigned(1980, 12), 1563 => to_unsigned(3276, 12), 1564 => to_unsigned(3955, 12), 1565 => to_unsigned(2291, 12), 1566 => to_unsigned(1727, 12), 1567 => to_unsigned(1049, 12), 1568 => to_unsigned(1841, 12), 1569 => to_unsigned(3601, 12), 1570 => to_unsigned(1360, 12), 1571 => to_unsigned(2319, 12), 1572 => to_unsigned(1014, 12), 1573 => to_unsigned(3865, 12), 1574 => to_unsigned(79, 12), 1575 => to_unsigned(3897, 12), 1576 => to_unsigned(2047, 12), 1577 => to_unsigned(1960, 12), 1578 => to_unsigned(2331, 12), 1579 => to_unsigned(3338, 12), 1580 => to_unsigned(3336, 12), 1581 => to_unsigned(1777, 12), 1582 => to_unsigned(1752, 12), 1583 => to_unsigned(510, 12), 1584 => to_unsigned(3732, 12), 1585 => to_unsigned(236, 12), 1586 => to_unsigned(3791, 12), 1587 => to_unsigned(222, 12), 1588 => to_unsigned(3251, 12), 1589 => to_unsigned(1881, 12), 1590 => to_unsigned(2532, 12), 1591 => to_unsigned(568, 12), 1592 => to_unsigned(3838, 12), 1593 => to_unsigned(3721, 12), 1594 => to_unsigned(2926, 12), 1595 => to_unsigned(2911, 12), 1596 => to_unsigned(163, 12), 1597 => to_unsigned(2505, 12), 1598 => to_unsigned(3465, 12), 1599 => to_unsigned(3856, 12), 1600 => to_unsigned(3175, 12), 1601 => to_unsigned(2829, 12), 1602 => to_unsigned(4065, 12), 1603 => to_unsigned(880, 12), 1604 => to_unsigned(552, 12), 1605 => to_unsigned(2401, 12), 1606 => to_unsigned(1647, 12), 1607 => to_unsigned(437, 12), 1608 => to_unsigned(2155, 12), 1609 => to_unsigned(4013, 12), 1610 => to_unsigned(2963, 12), 1611 => to_unsigned(3962, 12), 1612 => to_unsigned(2700, 12), 1613 => to_unsigned(3081, 12), 1614 => to_unsigned(2089, 12), 1615 => to_unsigned(2320, 12), 1616 => to_unsigned(35, 12), 1617 => to_unsigned(2373, 12), 1618 => to_unsigned(3045, 12), 1619 => to_unsigned(2977, 12), 1620 => to_unsigned(3619, 12), 1621 => to_unsigned(1477, 12), 1622 => to_unsigned(474, 12), 1623 => to_unsigned(93, 12), 1624 => to_unsigned(1329, 12), 1625 => to_unsigned(2336, 12), 1626 => to_unsigned(2811, 12), 1627 => to_unsigned(2478, 12), 1628 => to_unsigned(1356, 12), 1629 => to_unsigned(2467, 12), 1630 => to_unsigned(3691, 12), 1631 => to_unsigned(813, 12), 1632 => to_unsigned(2820, 12), 1633 => to_unsigned(2939, 12), 1634 => to_unsigned(3562, 12), 1635 => to_unsigned(773, 12), 1636 => to_unsigned(1961, 12), 1637 => to_unsigned(1369, 12), 1638 => to_unsigned(1881, 12), 1639 => to_unsigned(2230, 12), 1640 => to_unsigned(2101, 12), 1641 => to_unsigned(2051, 12), 1642 => to_unsigned(3628, 12), 1643 => to_unsigned(3611, 12), 1644 => to_unsigned(3417, 12), 1645 => to_unsigned(2348, 12), 1646 => to_unsigned(433, 12), 1647 => to_unsigned(1705, 12), 1648 => to_unsigned(978, 12), 1649 => to_unsigned(970, 12), 1650 => to_unsigned(4027, 12), 1651 => to_unsigned(1626, 12), 1652 => to_unsigned(84, 12), 1653 => to_unsigned(3808, 12), 1654 => to_unsigned(12, 12), 1655 => to_unsigned(1361, 12), 1656 => to_unsigned(2653, 12), 1657 => to_unsigned(2377, 12), 1658 => to_unsigned(4037, 12), 1659 => to_unsigned(194, 12), 1660 => to_unsigned(2753, 12), 1661 => to_unsigned(3768, 12), 1662 => to_unsigned(3171, 12), 1663 => to_unsigned(1811, 12), 1664 => to_unsigned(231, 12), 1665 => to_unsigned(148, 12), 1666 => to_unsigned(639, 12), 1667 => to_unsigned(3365, 12), 1668 => to_unsigned(2038, 12), 1669 => to_unsigned(267, 12), 1670 => to_unsigned(3730, 12), 1671 => to_unsigned(2679, 12), 1672 => to_unsigned(3874, 12), 1673 => to_unsigned(2102, 12), 1674 => to_unsigned(1689, 12), 1675 => to_unsigned(2642, 12), 1676 => to_unsigned(362, 12), 1677 => to_unsigned(1707, 12), 1678 => to_unsigned(4013, 12), 1679 => to_unsigned(4016, 12), 1680 => to_unsigned(1673, 12), 1681 => to_unsigned(3828, 12), 1682 => to_unsigned(3611, 12), 1683 => to_unsigned(1303, 12), 1684 => to_unsigned(1793, 12), 1685 => to_unsigned(1974, 12), 1686 => to_unsigned(3987, 12), 1687 => to_unsigned(3450, 12), 1688 => to_unsigned(774, 12), 1689 => to_unsigned(28, 12), 1690 => to_unsigned(3164, 12), 1691 => to_unsigned(3549, 12), 1692 => to_unsigned(1119, 12), 1693 => to_unsigned(3920, 12), 1694 => to_unsigned(2353, 12), 1695 => to_unsigned(357, 12), 1696 => to_unsigned(3695, 12), 1697 => to_unsigned(1639, 12), 1698 => to_unsigned(2148, 12), 1699 => to_unsigned(3243, 12), 1700 => to_unsigned(1055, 12), 1701 => to_unsigned(1089, 12), 1702 => to_unsigned(2298, 12), 1703 => to_unsigned(2968, 12), 1704 => to_unsigned(2082, 12), 1705 => to_unsigned(2429, 12), 1706 => to_unsigned(100, 12), 1707 => to_unsigned(1322, 12), 1708 => to_unsigned(203, 12), 1709 => to_unsigned(1243, 12), 1710 => to_unsigned(2289, 12), 1711 => to_unsigned(1503, 12), 1712 => to_unsigned(3752, 12), 1713 => to_unsigned(3328, 12), 1714 => to_unsigned(2755, 12), 1715 => to_unsigned(3394, 12), 1716 => to_unsigned(1090, 12), 1717 => to_unsigned(1325, 12), 1718 => to_unsigned(209, 12), 1719 => to_unsigned(780, 12), 1720 => to_unsigned(1012, 12), 1721 => to_unsigned(1383, 12), 1722 => to_unsigned(2537, 12), 1723 => to_unsigned(3415, 12), 1724 => to_unsigned(2310, 12), 1725 => to_unsigned(86, 12), 1726 => to_unsigned(828, 12), 1727 => to_unsigned(1663, 12), 1728 => to_unsigned(2099, 12), 1729 => to_unsigned(2616, 12), 1730 => to_unsigned(1230, 12), 1731 => to_unsigned(2989, 12), 1732 => to_unsigned(2368, 12), 1733 => to_unsigned(2172, 12), 1734 => to_unsigned(3988, 12), 1735 => to_unsigned(3364, 12), 1736 => to_unsigned(96, 12), 1737 => to_unsigned(740, 12), 1738 => to_unsigned(3602, 12), 1739 => to_unsigned(946, 12), 1740 => to_unsigned(1955, 12), 1741 => to_unsigned(3865, 12), 1742 => to_unsigned(1886, 12), 1743 => to_unsigned(2527, 12), 1744 => to_unsigned(510, 12), 1745 => to_unsigned(3771, 12), 1746 => to_unsigned(2045, 12), 1747 => to_unsigned(527, 12), 1748 => to_unsigned(1752, 12), 1749 => to_unsigned(790, 12), 1750 => to_unsigned(3906, 12), 1751 => to_unsigned(2071, 12), 1752 => to_unsigned(161, 12), 1753 => to_unsigned(3445, 12), 1754 => to_unsigned(3946, 12), 1755 => to_unsigned(2420, 12), 1756 => to_unsigned(456, 12), 1757 => to_unsigned(2665, 12), 1758 => to_unsigned(3503, 12), 1759 => to_unsigned(3387, 12), 1760 => to_unsigned(3437, 12), 1761 => to_unsigned(1464, 12), 1762 => to_unsigned(2511, 12), 1763 => to_unsigned(2067, 12), 1764 => to_unsigned(2126, 12), 1765 => to_unsigned(3366, 12), 1766 => to_unsigned(1061, 12), 1767 => to_unsigned(2851, 12), 1768 => to_unsigned(3339, 12), 1769 => to_unsigned(870, 12), 1770 => to_unsigned(2716, 12), 1771 => to_unsigned(227, 12), 1772 => to_unsigned(3882, 12), 1773 => to_unsigned(1247, 12), 1774 => to_unsigned(3757, 12), 1775 => to_unsigned(3281, 12), 1776 => to_unsigned(2601, 12), 1777 => to_unsigned(2382, 12), 1778 => to_unsigned(3624, 12), 1779 => to_unsigned(1138, 12), 1780 => to_unsigned(2979, 12), 1781 => to_unsigned(3262, 12), 1782 => to_unsigned(1445, 12), 1783 => to_unsigned(3807, 12), 1784 => to_unsigned(2615, 12), 1785 => to_unsigned(2850, 12), 1786 => to_unsigned(2798, 12), 1787 => to_unsigned(2335, 12), 1788 => to_unsigned(2515, 12), 1789 => to_unsigned(3475, 12), 1790 => to_unsigned(3385, 12), 1791 => to_unsigned(613, 12), 1792 => to_unsigned(3095, 12), 1793 => to_unsigned(588, 12), 1794 => to_unsigned(238, 12), 1795 => to_unsigned(1104, 12), 1796 => to_unsigned(2913, 12), 1797 => to_unsigned(1975, 12), 1798 => to_unsigned(3614, 12), 1799 => to_unsigned(2139, 12), 1800 => to_unsigned(3576, 12), 1801 => to_unsigned(2278, 12), 1802 => to_unsigned(2435, 12), 1803 => to_unsigned(854, 12), 1804 => to_unsigned(3457, 12), 1805 => to_unsigned(1550, 12), 1806 => to_unsigned(2971, 12), 1807 => to_unsigned(3712, 12), 1808 => to_unsigned(3819, 12), 1809 => to_unsigned(3081, 12), 1810 => to_unsigned(2339, 12), 1811 => to_unsigned(2894, 12), 1812 => to_unsigned(3616, 12), 1813 => to_unsigned(1722, 12), 1814 => to_unsigned(3738, 12), 1815 => to_unsigned(268, 12), 1816 => to_unsigned(820, 12), 1817 => to_unsigned(953, 12), 1818 => to_unsigned(1197, 12), 1819 => to_unsigned(3918, 12), 1820 => to_unsigned(3091, 12), 1821 => to_unsigned(2653, 12), 1822 => to_unsigned(2035, 12), 1823 => to_unsigned(1398, 12), 1824 => to_unsigned(891, 12), 1825 => to_unsigned(1873, 12), 1826 => to_unsigned(70, 12), 1827 => to_unsigned(2287, 12), 1828 => to_unsigned(161, 12), 1829 => to_unsigned(3277, 12), 1830 => to_unsigned(214, 12), 1831 => to_unsigned(3371, 12), 1832 => to_unsigned(1792, 12), 1833 => to_unsigned(1081, 12), 1834 => to_unsigned(662, 12), 1835 => to_unsigned(1262, 12), 1836 => to_unsigned(782, 12), 1837 => to_unsigned(868, 12), 1838 => to_unsigned(3576, 12), 1839 => to_unsigned(1605, 12), 1840 => to_unsigned(1290, 12), 1841 => to_unsigned(67, 12), 1842 => to_unsigned(4, 12), 1843 => to_unsigned(2228, 12), 1844 => to_unsigned(2108, 12), 1845 => to_unsigned(308, 12), 1846 => to_unsigned(959, 12), 1847 => to_unsigned(1758, 12), 1848 => to_unsigned(389, 12), 1849 => to_unsigned(1547, 12), 1850 => to_unsigned(60, 12), 1851 => to_unsigned(1165, 12), 1852 => to_unsigned(652, 12), 1853 => to_unsigned(2951, 12), 1854 => to_unsigned(1336, 12), 1855 => to_unsigned(1413, 12), 1856 => to_unsigned(3897, 12), 1857 => to_unsigned(906, 12), 1858 => to_unsigned(1438, 12), 1859 => to_unsigned(1411, 12), 1860 => to_unsigned(1762, 12), 1861 => to_unsigned(2426, 12), 1862 => to_unsigned(1341, 12), 1863 => to_unsigned(1665, 12), 1864 => to_unsigned(3883, 12), 1865 => to_unsigned(1424, 12), 1866 => to_unsigned(1959, 12), 1867 => to_unsigned(3985, 12), 1868 => to_unsigned(2612, 12), 1869 => to_unsigned(3054, 12), 1870 => to_unsigned(436, 12), 1871 => to_unsigned(2682, 12), 1872 => to_unsigned(880, 12), 1873 => to_unsigned(1543, 12), 1874 => to_unsigned(2194, 12), 1875 => to_unsigned(3477, 12), 1876 => to_unsigned(3734, 12), 1877 => to_unsigned(3870, 12), 1878 => to_unsigned(1348, 12), 1879 => to_unsigned(863, 12), 1880 => to_unsigned(3459, 12), 1881 => to_unsigned(689, 12), 1882 => to_unsigned(1776, 12), 1883 => to_unsigned(137, 12), 1884 => to_unsigned(1161, 12), 1885 => to_unsigned(2722, 12), 1886 => to_unsigned(3814, 12), 1887 => to_unsigned(1271, 12), 1888 => to_unsigned(3934, 12), 1889 => to_unsigned(3148, 12), 1890 => to_unsigned(2480, 12), 1891 => to_unsigned(4017, 12), 1892 => to_unsigned(2184, 12), 1893 => to_unsigned(2943, 12), 1894 => to_unsigned(3063, 12), 1895 => to_unsigned(238, 12), 1896 => to_unsigned(24, 12), 1897 => to_unsigned(1188, 12), 1898 => to_unsigned(1143, 12), 1899 => to_unsigned(3337, 12), 1900 => to_unsigned(6, 12), 1901 => to_unsigned(1800, 12), 1902 => to_unsigned(1784, 12), 1903 => to_unsigned(1105, 12), 1904 => to_unsigned(2377, 12), 1905 => to_unsigned(953, 12), 1906 => to_unsigned(3962, 12), 1907 => to_unsigned(1153, 12), 1908 => to_unsigned(3748, 12), 1909 => to_unsigned(3072, 12), 1910 => to_unsigned(2618, 12), 1911 => to_unsigned(2345, 12), 1912 => to_unsigned(2766, 12), 1913 => to_unsigned(2614, 12), 1914 => to_unsigned(3547, 12), 1915 => to_unsigned(3610, 12), 1916 => to_unsigned(1698, 12), 1917 => to_unsigned(1221, 12), 1918 => to_unsigned(3198, 12), 1919 => to_unsigned(7, 12), 1920 => to_unsigned(754, 12), 1921 => to_unsigned(210, 12), 1922 => to_unsigned(2296, 12), 1923 => to_unsigned(2959, 12), 1924 => to_unsigned(1181, 12), 1925 => to_unsigned(511, 12), 1926 => to_unsigned(3302, 12), 1927 => to_unsigned(3280, 12), 1928 => to_unsigned(2877, 12), 1929 => to_unsigned(562, 12), 1930 => to_unsigned(2819, 12), 1931 => to_unsigned(1713, 12), 1932 => to_unsigned(453, 12), 1933 => to_unsigned(485, 12), 1934 => to_unsigned(602, 12), 1935 => to_unsigned(674, 12), 1936 => to_unsigned(2401, 12), 1937 => to_unsigned(3288, 12), 1938 => to_unsigned(437, 12), 1939 => to_unsigned(298, 12), 1940 => to_unsigned(1698, 12), 1941 => to_unsigned(202, 12), 1942 => to_unsigned(3906, 12), 1943 => to_unsigned(577, 12), 1944 => to_unsigned(960, 12), 1945 => to_unsigned(2987, 12), 1946 => to_unsigned(505, 12), 1947 => to_unsigned(1291, 12), 1948 => to_unsigned(3958, 12), 1949 => to_unsigned(1863, 12), 1950 => to_unsigned(2467, 12), 1951 => to_unsigned(3729, 12), 1952 => to_unsigned(3944, 12), 1953 => to_unsigned(456, 12), 1954 => to_unsigned(3109, 12), 1955 => to_unsigned(288, 12), 1956 => to_unsigned(1217, 12), 1957 => to_unsigned(1641, 12), 1958 => to_unsigned(516, 12), 1959 => to_unsigned(3822, 12), 1960 => to_unsigned(209, 12), 1961 => to_unsigned(2524, 12), 1962 => to_unsigned(443, 12), 1963 => to_unsigned(2911, 12), 1964 => to_unsigned(209, 12), 1965 => to_unsigned(164, 12), 1966 => to_unsigned(1472, 12), 1967 => to_unsigned(2285, 12), 1968 => to_unsigned(2131, 12), 1969 => to_unsigned(1305, 12), 1970 => to_unsigned(2077, 12), 1971 => to_unsigned(2303, 12), 1972 => to_unsigned(263, 12), 1973 => to_unsigned(1626, 12), 1974 => to_unsigned(2438, 12), 1975 => to_unsigned(1183, 12), 1976 => to_unsigned(443, 12), 1977 => to_unsigned(3053, 12), 1978 => to_unsigned(67, 12), 1979 => to_unsigned(3332, 12), 1980 => to_unsigned(769, 12), 1981 => to_unsigned(2636, 12), 1982 => to_unsigned(3059, 12), 1983 => to_unsigned(648, 12), 1984 => to_unsigned(3903, 12), 1985 => to_unsigned(1313, 12), 1986 => to_unsigned(161, 12), 1987 => to_unsigned(3447, 12), 1988 => to_unsigned(29, 12), 1989 => to_unsigned(1949, 12), 1990 => to_unsigned(3798, 12), 1991 => to_unsigned(1855, 12), 1992 => to_unsigned(1433, 12), 1993 => to_unsigned(1117, 12), 1994 => to_unsigned(2616, 12), 1995 => to_unsigned(2243, 12), 1996 => to_unsigned(3434, 12), 1997 => to_unsigned(347, 12), 1998 => to_unsigned(3368, 12), 1999 => to_unsigned(2804, 12), 2000 => to_unsigned(108, 12), 2001 => to_unsigned(269, 12), 2002 => to_unsigned(1114, 12), 2003 => to_unsigned(1196, 12), 2004 => to_unsigned(536, 12), 2005 => to_unsigned(3426, 12), 2006 => to_unsigned(2224, 12), 2007 => to_unsigned(2713, 12), 2008 => to_unsigned(2748, 12), 2009 => to_unsigned(1445, 12), 2010 => to_unsigned(503, 12), 2011 => to_unsigned(2079, 12), 2012 => to_unsigned(3599, 12), 2013 => to_unsigned(2262, 12), 2014 => to_unsigned(481, 12), 2015 => to_unsigned(3211, 12), 2016 => to_unsigned(2022, 12), 2017 => to_unsigned(2022, 12), 2018 => to_unsigned(3217, 12), 2019 => to_unsigned(284, 12), 2020 => to_unsigned(3371, 12), 2021 => to_unsigned(1663, 12), 2022 => to_unsigned(3860, 12), 2023 => to_unsigned(364, 12), 2024 => to_unsigned(3108, 12), 2025 => to_unsigned(1288, 12), 2026 => to_unsigned(2351, 12), 2027 => to_unsigned(3845, 12), 2028 => to_unsigned(2590, 12), 2029 => to_unsigned(3772, 12), 2030 => to_unsigned(4019, 12), 2031 => to_unsigned(175, 12), 2032 => to_unsigned(3891, 12), 2033 => to_unsigned(2562, 12), 2034 => to_unsigned(2260, 12), 2035 => to_unsigned(856, 12), 2036 => to_unsigned(3564, 12), 2037 => to_unsigned(909, 12), 2038 => to_unsigned(702, 12), 2039 => to_unsigned(3411, 12), 2040 => to_unsigned(3617, 12), 2041 => to_unsigned(2854, 12), 2042 => to_unsigned(988, 12), 2043 => to_unsigned(1104, 12), 2044 => to_unsigned(1299, 12), 2045 => to_unsigned(1700, 12), 2046 => to_unsigned(2319, 12), 2047 => to_unsigned(2725, 12)),
            5 => (0 => to_unsigned(2166, 12), 1 => to_unsigned(870, 12), 2 => to_unsigned(266, 12), 3 => to_unsigned(2793, 12), 4 => to_unsigned(1526, 12), 5 => to_unsigned(2355, 12), 6 => to_unsigned(4090, 12), 7 => to_unsigned(1171, 12), 8 => to_unsigned(3765, 12), 9 => to_unsigned(3497, 12), 10 => to_unsigned(1914, 12), 11 => to_unsigned(2026, 12), 12 => to_unsigned(2825, 12), 13 => to_unsigned(4045, 12), 14 => to_unsigned(73, 12), 15 => to_unsigned(669, 12), 16 => to_unsigned(65, 12), 17 => to_unsigned(891, 12), 18 => to_unsigned(373, 12), 19 => to_unsigned(311, 12), 20 => to_unsigned(83, 12), 21 => to_unsigned(2144, 12), 22 => to_unsigned(1442, 12), 23 => to_unsigned(570, 12), 24 => to_unsigned(3230, 12), 25 => to_unsigned(4021, 12), 26 => to_unsigned(804, 12), 27 => to_unsigned(3482, 12), 28 => to_unsigned(680, 12), 29 => to_unsigned(1152, 12), 30 => to_unsigned(3473, 12), 31 => to_unsigned(2874, 12), 32 => to_unsigned(1503, 12), 33 => to_unsigned(3031, 12), 34 => to_unsigned(2080, 12), 35 => to_unsigned(2065, 12), 36 => to_unsigned(455, 12), 37 => to_unsigned(3335, 12), 38 => to_unsigned(374, 12), 39 => to_unsigned(949, 12), 40 => to_unsigned(1680, 12), 41 => to_unsigned(3711, 12), 42 => to_unsigned(874, 12), 43 => to_unsigned(2078, 12), 44 => to_unsigned(3358, 12), 45 => to_unsigned(502, 12), 46 => to_unsigned(930, 12), 47 => to_unsigned(409, 12), 48 => to_unsigned(3922, 12), 49 => to_unsigned(1737, 12), 50 => to_unsigned(3026, 12), 51 => to_unsigned(3732, 12), 52 => to_unsigned(1209, 12), 53 => to_unsigned(204, 12), 54 => to_unsigned(783, 12), 55 => to_unsigned(1749, 12), 56 => to_unsigned(682, 12), 57 => to_unsigned(678, 12), 58 => to_unsigned(1429, 12), 59 => to_unsigned(2187, 12), 60 => to_unsigned(3314, 12), 61 => to_unsigned(3397, 12), 62 => to_unsigned(3157, 12), 63 => to_unsigned(1142, 12), 64 => to_unsigned(2518, 12), 65 => to_unsigned(107, 12), 66 => to_unsigned(2522, 12), 67 => to_unsigned(3985, 12), 68 => to_unsigned(968, 12), 69 => to_unsigned(785, 12), 70 => to_unsigned(661, 12), 71 => to_unsigned(3891, 12), 72 => to_unsigned(2306, 12), 73 => to_unsigned(3642, 12), 74 => to_unsigned(3055, 12), 75 => to_unsigned(3002, 12), 76 => to_unsigned(1584, 12), 77 => to_unsigned(3568, 12), 78 => to_unsigned(2601, 12), 79 => to_unsigned(1821, 12), 80 => to_unsigned(3801, 12), 81 => to_unsigned(3027, 12), 82 => to_unsigned(1888, 12), 83 => to_unsigned(1100, 12), 84 => to_unsigned(3633, 12), 85 => to_unsigned(687, 12), 86 => to_unsigned(2165, 12), 87 => to_unsigned(2598, 12), 88 => to_unsigned(1836, 12), 89 => to_unsigned(3665, 12), 90 => to_unsigned(383, 12), 91 => to_unsigned(1693, 12), 92 => to_unsigned(3396, 12), 93 => to_unsigned(918, 12), 94 => to_unsigned(1230, 12), 95 => to_unsigned(2212, 12), 96 => to_unsigned(2225, 12), 97 => to_unsigned(464, 12), 98 => to_unsigned(79, 12), 99 => to_unsigned(1439, 12), 100 => to_unsigned(2961, 12), 101 => to_unsigned(2112, 12), 102 => to_unsigned(2575, 12), 103 => to_unsigned(2498, 12), 104 => to_unsigned(3933, 12), 105 => to_unsigned(2919, 12), 106 => to_unsigned(4013, 12), 107 => to_unsigned(2234, 12), 108 => to_unsigned(2850, 12), 109 => to_unsigned(1918, 12), 110 => to_unsigned(2125, 12), 111 => to_unsigned(434, 12), 112 => to_unsigned(1147, 12), 113 => to_unsigned(734, 12), 114 => to_unsigned(963, 12), 115 => to_unsigned(2401, 12), 116 => to_unsigned(2870, 12), 117 => to_unsigned(1140, 12), 118 => to_unsigned(1251, 12), 119 => to_unsigned(1339, 12), 120 => to_unsigned(3708, 12), 121 => to_unsigned(2451, 12), 122 => to_unsigned(1028, 12), 123 => to_unsigned(3275, 12), 124 => to_unsigned(1202, 12), 125 => to_unsigned(2981, 12), 126 => to_unsigned(590, 12), 127 => to_unsigned(2223, 12), 128 => to_unsigned(1484, 12), 129 => to_unsigned(3942, 12), 130 => to_unsigned(682, 12), 131 => to_unsigned(2865, 12), 132 => to_unsigned(1564, 12), 133 => to_unsigned(2644, 12), 134 => to_unsigned(3296, 12), 135 => to_unsigned(875, 12), 136 => to_unsigned(1926, 12), 137 => to_unsigned(1660, 12), 138 => to_unsigned(1486, 12), 139 => to_unsigned(1776, 12), 140 => to_unsigned(3301, 12), 141 => to_unsigned(2488, 12), 142 => to_unsigned(2360, 12), 143 => to_unsigned(2733, 12), 144 => to_unsigned(770, 12), 145 => to_unsigned(2040, 12), 146 => to_unsigned(1972, 12), 147 => to_unsigned(3913, 12), 148 => to_unsigned(539, 12), 149 => to_unsigned(879, 12), 150 => to_unsigned(861, 12), 151 => to_unsigned(1314, 12), 152 => to_unsigned(1925, 12), 153 => to_unsigned(3384, 12), 154 => to_unsigned(2328, 12), 155 => to_unsigned(2218, 12), 156 => to_unsigned(2605, 12), 157 => to_unsigned(3274, 12), 158 => to_unsigned(493, 12), 159 => to_unsigned(2572, 12), 160 => to_unsigned(1028, 12), 161 => to_unsigned(3830, 12), 162 => to_unsigned(3809, 12), 163 => to_unsigned(100, 12), 164 => to_unsigned(1700, 12), 165 => to_unsigned(93, 12), 166 => to_unsigned(1702, 12), 167 => to_unsigned(1354, 12), 168 => to_unsigned(3626, 12), 169 => to_unsigned(803, 12), 170 => to_unsigned(1890, 12), 171 => to_unsigned(570, 12), 172 => to_unsigned(2764, 12), 173 => to_unsigned(533, 12), 174 => to_unsigned(3654, 12), 175 => to_unsigned(479, 12), 176 => to_unsigned(2700, 12), 177 => to_unsigned(1322, 12), 178 => to_unsigned(3778, 12), 179 => to_unsigned(1971, 12), 180 => to_unsigned(1175, 12), 181 => to_unsigned(2968, 12), 182 => to_unsigned(3455, 12), 183 => to_unsigned(3914, 12), 184 => to_unsigned(1265, 12), 185 => to_unsigned(3787, 12), 186 => to_unsigned(54, 12), 187 => to_unsigned(3176, 12), 188 => to_unsigned(3509, 12), 189 => to_unsigned(964, 12), 190 => to_unsigned(2274, 12), 191 => to_unsigned(593, 12), 192 => to_unsigned(1604, 12), 193 => to_unsigned(3226, 12), 194 => to_unsigned(2600, 12), 195 => to_unsigned(775, 12), 196 => to_unsigned(3202, 12), 197 => to_unsigned(2037, 12), 198 => to_unsigned(1122, 12), 199 => to_unsigned(3169, 12), 200 => to_unsigned(171, 12), 201 => to_unsigned(2516, 12), 202 => to_unsigned(285, 12), 203 => to_unsigned(2796, 12), 204 => to_unsigned(1858, 12), 205 => to_unsigned(3534, 12), 206 => to_unsigned(753, 12), 207 => to_unsigned(2931, 12), 208 => to_unsigned(1226, 12), 209 => to_unsigned(1228, 12), 210 => to_unsigned(2522, 12), 211 => to_unsigned(3886, 12), 212 => to_unsigned(1959, 12), 213 => to_unsigned(880, 12), 214 => to_unsigned(1333, 12), 215 => to_unsigned(4086, 12), 216 => to_unsigned(1038, 12), 217 => to_unsigned(1182, 12), 218 => to_unsigned(1987, 12), 219 => to_unsigned(1742, 12), 220 => to_unsigned(2026, 12), 221 => to_unsigned(241, 12), 222 => to_unsigned(917, 12), 223 => to_unsigned(1956, 12), 224 => to_unsigned(69, 12), 225 => to_unsigned(2472, 12), 226 => to_unsigned(1265, 12), 227 => to_unsigned(3692, 12), 228 => to_unsigned(3216, 12), 229 => to_unsigned(1790, 12), 230 => to_unsigned(3847, 12), 231 => to_unsigned(980, 12), 232 => to_unsigned(1683, 12), 233 => to_unsigned(3330, 12), 234 => to_unsigned(316, 12), 235 => to_unsigned(1696, 12), 236 => to_unsigned(3683, 12), 237 => to_unsigned(658, 12), 238 => to_unsigned(51, 12), 239 => to_unsigned(3631, 12), 240 => to_unsigned(1913, 12), 241 => to_unsigned(2621, 12), 242 => to_unsigned(1937, 12), 243 => to_unsigned(1858, 12), 244 => to_unsigned(694, 12), 245 => to_unsigned(777, 12), 246 => to_unsigned(682, 12), 247 => to_unsigned(2374, 12), 248 => to_unsigned(1045, 12), 249 => to_unsigned(2481, 12), 250 => to_unsigned(1325, 12), 251 => to_unsigned(3335, 12), 252 => to_unsigned(3541, 12), 253 => to_unsigned(585, 12), 254 => to_unsigned(2159, 12), 255 => to_unsigned(2777, 12), 256 => to_unsigned(1938, 12), 257 => to_unsigned(1526, 12), 258 => to_unsigned(444, 12), 259 => to_unsigned(3783, 12), 260 => to_unsigned(3022, 12), 261 => to_unsigned(260, 12), 262 => to_unsigned(1137, 12), 263 => to_unsigned(2012, 12), 264 => to_unsigned(3283, 12), 265 => to_unsigned(2761, 12), 266 => to_unsigned(731, 12), 267 => to_unsigned(2708, 12), 268 => to_unsigned(4034, 12), 269 => to_unsigned(781, 12), 270 => to_unsigned(445, 12), 271 => to_unsigned(1910, 12), 272 => to_unsigned(3296, 12), 273 => to_unsigned(2703, 12), 274 => to_unsigned(3706, 12), 275 => to_unsigned(2738, 12), 276 => to_unsigned(3125, 12), 277 => to_unsigned(3909, 12), 278 => to_unsigned(3788, 12), 279 => to_unsigned(3242, 12), 280 => to_unsigned(933, 12), 281 => to_unsigned(3717, 12), 282 => to_unsigned(820, 12), 283 => to_unsigned(1648, 12), 284 => to_unsigned(1596, 12), 285 => to_unsigned(3899, 12), 286 => to_unsigned(3870, 12), 287 => to_unsigned(1159, 12), 288 => to_unsigned(3284, 12), 289 => to_unsigned(851, 12), 290 => to_unsigned(3362, 12), 291 => to_unsigned(2586, 12), 292 => to_unsigned(1319, 12), 293 => to_unsigned(971, 12), 294 => to_unsigned(3666, 12), 295 => to_unsigned(3729, 12), 296 => to_unsigned(3455, 12), 297 => to_unsigned(3776, 12), 298 => to_unsigned(3182, 12), 299 => to_unsigned(2749, 12), 300 => to_unsigned(1590, 12), 301 => to_unsigned(644, 12), 302 => to_unsigned(2000, 12), 303 => to_unsigned(4074, 12), 304 => to_unsigned(1080, 12), 305 => to_unsigned(729, 12), 306 => to_unsigned(737, 12), 307 => to_unsigned(412, 12), 308 => to_unsigned(378, 12), 309 => to_unsigned(3438, 12), 310 => to_unsigned(1250, 12), 311 => to_unsigned(2961, 12), 312 => to_unsigned(1159, 12), 313 => to_unsigned(3243, 12), 314 => to_unsigned(3264, 12), 315 => to_unsigned(1329, 12), 316 => to_unsigned(2504, 12), 317 => to_unsigned(3540, 12), 318 => to_unsigned(513, 12), 319 => to_unsigned(3813, 12), 320 => to_unsigned(2556, 12), 321 => to_unsigned(2715, 12), 322 => to_unsigned(171, 12), 323 => to_unsigned(3386, 12), 324 => to_unsigned(1807, 12), 325 => to_unsigned(2996, 12), 326 => to_unsigned(1545, 12), 327 => to_unsigned(792, 12), 328 => to_unsigned(968, 12), 329 => to_unsigned(2924, 12), 330 => to_unsigned(89, 12), 331 => to_unsigned(2802, 12), 332 => to_unsigned(3043, 12), 333 => to_unsigned(2734, 12), 334 => to_unsigned(1499, 12), 335 => to_unsigned(1378, 12), 336 => to_unsigned(3117, 12), 337 => to_unsigned(577, 12), 338 => to_unsigned(4022, 12), 339 => to_unsigned(1224, 12), 340 => to_unsigned(719, 12), 341 => to_unsigned(3736, 12), 342 => to_unsigned(2173, 12), 343 => to_unsigned(629, 12), 344 => to_unsigned(3080, 12), 345 => to_unsigned(2961, 12), 346 => to_unsigned(1657, 12), 347 => to_unsigned(295, 12), 348 => to_unsigned(596, 12), 349 => to_unsigned(3078, 12), 350 => to_unsigned(1252, 12), 351 => to_unsigned(1326, 12), 352 => to_unsigned(3026, 12), 353 => to_unsigned(2714, 12), 354 => to_unsigned(1264, 12), 355 => to_unsigned(1615, 12), 356 => to_unsigned(7, 12), 357 => to_unsigned(1409, 12), 358 => to_unsigned(2332, 12), 359 => to_unsigned(1296, 12), 360 => to_unsigned(2205, 12), 361 => to_unsigned(3916, 12), 362 => to_unsigned(353, 12), 363 => to_unsigned(2177, 12), 364 => to_unsigned(3570, 12), 365 => to_unsigned(2717, 12), 366 => to_unsigned(1198, 12), 367 => to_unsigned(606, 12), 368 => to_unsigned(2001, 12), 369 => to_unsigned(2417, 12), 370 => to_unsigned(3461, 12), 371 => to_unsigned(1429, 12), 372 => to_unsigned(3973, 12), 373 => to_unsigned(1015, 12), 374 => to_unsigned(3672, 12), 375 => to_unsigned(2025, 12), 376 => to_unsigned(2447, 12), 377 => to_unsigned(3382, 12), 378 => to_unsigned(4071, 12), 379 => to_unsigned(2027, 12), 380 => to_unsigned(2920, 12), 381 => to_unsigned(301, 12), 382 => to_unsigned(599, 12), 383 => to_unsigned(3631, 12), 384 => to_unsigned(2517, 12), 385 => to_unsigned(1066, 12), 386 => to_unsigned(1174, 12), 387 => to_unsigned(2792, 12), 388 => to_unsigned(1056, 12), 389 => to_unsigned(1993, 12), 390 => to_unsigned(3432, 12), 391 => to_unsigned(1244, 12), 392 => to_unsigned(3643, 12), 393 => to_unsigned(3375, 12), 394 => to_unsigned(877, 12), 395 => to_unsigned(3740, 12), 396 => to_unsigned(2698, 12), 397 => to_unsigned(789, 12), 398 => to_unsigned(715, 12), 399 => to_unsigned(3449, 12), 400 => to_unsigned(2451, 12), 401 => to_unsigned(3919, 12), 402 => to_unsigned(137, 12), 403 => to_unsigned(2072, 12), 404 => to_unsigned(2353, 12), 405 => to_unsigned(2866, 12), 406 => to_unsigned(2484, 12), 407 => to_unsigned(3027, 12), 408 => to_unsigned(3342, 12), 409 => to_unsigned(2404, 12), 410 => to_unsigned(287, 12), 411 => to_unsigned(1990, 12), 412 => to_unsigned(1381, 12), 413 => to_unsigned(797, 12), 414 => to_unsigned(2276, 12), 415 => to_unsigned(933, 12), 416 => to_unsigned(2684, 12), 417 => to_unsigned(2221, 12), 418 => to_unsigned(4060, 12), 419 => to_unsigned(80, 12), 420 => to_unsigned(2618, 12), 421 => to_unsigned(3333, 12), 422 => to_unsigned(594, 12), 423 => to_unsigned(3761, 12), 424 => to_unsigned(209, 12), 425 => to_unsigned(1185, 12), 426 => to_unsigned(474, 12), 427 => to_unsigned(983, 12), 428 => to_unsigned(3178, 12), 429 => to_unsigned(306, 12), 430 => to_unsigned(3577, 12), 431 => to_unsigned(16, 12), 432 => to_unsigned(3669, 12), 433 => to_unsigned(1325, 12), 434 => to_unsigned(428, 12), 435 => to_unsigned(2197, 12), 436 => to_unsigned(2479, 12), 437 => to_unsigned(2842, 12), 438 => to_unsigned(3118, 12), 439 => to_unsigned(1394, 12), 440 => to_unsigned(1515, 12), 441 => to_unsigned(730, 12), 442 => to_unsigned(1284, 12), 443 => to_unsigned(550, 12), 444 => to_unsigned(1357, 12), 445 => to_unsigned(1609, 12), 446 => to_unsigned(2374, 12), 447 => to_unsigned(291, 12), 448 => to_unsigned(3084, 12), 449 => to_unsigned(2693, 12), 450 => to_unsigned(991, 12), 451 => to_unsigned(3128, 12), 452 => to_unsigned(1820, 12), 453 => to_unsigned(1234, 12), 454 => to_unsigned(958, 12), 455 => to_unsigned(729, 12), 456 => to_unsigned(3036, 12), 457 => to_unsigned(1251, 12), 458 => to_unsigned(1900, 12), 459 => to_unsigned(1039, 12), 460 => to_unsigned(351, 12), 461 => to_unsigned(1967, 12), 462 => to_unsigned(291, 12), 463 => to_unsigned(1531, 12), 464 => to_unsigned(766, 12), 465 => to_unsigned(3804, 12), 466 => to_unsigned(607, 12), 467 => to_unsigned(2187, 12), 468 => to_unsigned(153, 12), 469 => to_unsigned(3602, 12), 470 => to_unsigned(3680, 12), 471 => to_unsigned(1084, 12), 472 => to_unsigned(483, 12), 473 => to_unsigned(90, 12), 474 => to_unsigned(1843, 12), 475 => to_unsigned(2938, 12), 476 => to_unsigned(478, 12), 477 => to_unsigned(68, 12), 478 => to_unsigned(939, 12), 479 => to_unsigned(2318, 12), 480 => to_unsigned(261, 12), 481 => to_unsigned(3040, 12), 482 => to_unsigned(2176, 12), 483 => to_unsigned(2222, 12), 484 => to_unsigned(260, 12), 485 => to_unsigned(829, 12), 486 => to_unsigned(3861, 12), 487 => to_unsigned(1787, 12), 488 => to_unsigned(1236, 12), 489 => to_unsigned(2610, 12), 490 => to_unsigned(383, 12), 491 => to_unsigned(1135, 12), 492 => to_unsigned(615, 12), 493 => to_unsigned(14, 12), 494 => to_unsigned(1207, 12), 495 => to_unsigned(3781, 12), 496 => to_unsigned(1420, 12), 497 => to_unsigned(3696, 12), 498 => to_unsigned(3513, 12), 499 => to_unsigned(515, 12), 500 => to_unsigned(2845, 12), 501 => to_unsigned(2849, 12), 502 => to_unsigned(1840, 12), 503 => to_unsigned(2937, 12), 504 => to_unsigned(1701, 12), 505 => to_unsigned(786, 12), 506 => to_unsigned(1225, 12), 507 => to_unsigned(2212, 12), 508 => to_unsigned(624, 12), 509 => to_unsigned(67, 12), 510 => to_unsigned(752, 12), 511 => to_unsigned(1157, 12), 512 => to_unsigned(4028, 12), 513 => to_unsigned(575, 12), 514 => to_unsigned(200, 12), 515 => to_unsigned(2761, 12), 516 => to_unsigned(2449, 12), 517 => to_unsigned(1386, 12), 518 => to_unsigned(3942, 12), 519 => to_unsigned(1135, 12), 520 => to_unsigned(3543, 12), 521 => to_unsigned(3948, 12), 522 => to_unsigned(3060, 12), 523 => to_unsigned(1475, 12), 524 => to_unsigned(1639, 12), 525 => to_unsigned(3587, 12), 526 => to_unsigned(1771, 12), 527 => to_unsigned(3653, 12), 528 => to_unsigned(684, 12), 529 => to_unsigned(2554, 12), 530 => to_unsigned(2507, 12), 531 => to_unsigned(553, 12), 532 => to_unsigned(3006, 12), 533 => to_unsigned(299, 12), 534 => to_unsigned(2939, 12), 535 => to_unsigned(2020, 12), 536 => to_unsigned(2127, 12), 537 => to_unsigned(862, 12), 538 => to_unsigned(3456, 12), 539 => to_unsigned(3728, 12), 540 => to_unsigned(502, 12), 541 => to_unsigned(2209, 12), 542 => to_unsigned(173, 12), 543 => to_unsigned(2603, 12), 544 => to_unsigned(583, 12), 545 => to_unsigned(1105, 12), 546 => to_unsigned(3493, 12), 547 => to_unsigned(3241, 12), 548 => to_unsigned(1318, 12), 549 => to_unsigned(35, 12), 550 => to_unsigned(1329, 12), 551 => to_unsigned(209, 12), 552 => to_unsigned(527, 12), 553 => to_unsigned(2102, 12), 554 => to_unsigned(2602, 12), 555 => to_unsigned(345, 12), 556 => to_unsigned(3400, 12), 557 => to_unsigned(685, 12), 558 => to_unsigned(2989, 12), 559 => to_unsigned(2191, 12), 560 => to_unsigned(3006, 12), 561 => to_unsigned(1263, 12), 562 => to_unsigned(3194, 12), 563 => to_unsigned(2612, 12), 564 => to_unsigned(3435, 12), 565 => to_unsigned(3812, 12), 566 => to_unsigned(291, 12), 567 => to_unsigned(2658, 12), 568 => to_unsigned(2156, 12), 569 => to_unsigned(1848, 12), 570 => to_unsigned(2945, 12), 571 => to_unsigned(3062, 12), 572 => to_unsigned(3811, 12), 573 => to_unsigned(4023, 12), 574 => to_unsigned(92, 12), 575 => to_unsigned(2587, 12), 576 => to_unsigned(1277, 12), 577 => to_unsigned(2943, 12), 578 => to_unsigned(1193, 12), 579 => to_unsigned(3314, 12), 580 => to_unsigned(514, 12), 581 => to_unsigned(2190, 12), 582 => to_unsigned(3352, 12), 583 => to_unsigned(984, 12), 584 => to_unsigned(3562, 12), 585 => to_unsigned(1023, 12), 586 => to_unsigned(3091, 12), 587 => to_unsigned(1925, 12), 588 => to_unsigned(2147, 12), 589 => to_unsigned(123, 12), 590 => to_unsigned(2339, 12), 591 => to_unsigned(1953, 12), 592 => to_unsigned(2266, 12), 593 => to_unsigned(1228, 12), 594 => to_unsigned(3738, 12), 595 => to_unsigned(3950, 12), 596 => to_unsigned(3855, 12), 597 => to_unsigned(1448, 12), 598 => to_unsigned(3173, 12), 599 => to_unsigned(1039, 12), 600 => to_unsigned(4003, 12), 601 => to_unsigned(3925, 12), 602 => to_unsigned(1949, 12), 603 => to_unsigned(3222, 12), 604 => to_unsigned(3770, 12), 605 => to_unsigned(123, 12), 606 => to_unsigned(4013, 12), 607 => to_unsigned(742, 12), 608 => to_unsigned(3, 12), 609 => to_unsigned(1625, 12), 610 => to_unsigned(3919, 12), 611 => to_unsigned(217, 12), 612 => to_unsigned(2755, 12), 613 => to_unsigned(3130, 12), 614 => to_unsigned(2285, 12), 615 => to_unsigned(916, 12), 616 => to_unsigned(1977, 12), 617 => to_unsigned(1212, 12), 618 => to_unsigned(3820, 12), 619 => to_unsigned(279, 12), 620 => to_unsigned(2691, 12), 621 => to_unsigned(1879, 12), 622 => to_unsigned(2913, 12), 623 => to_unsigned(1987, 12), 624 => to_unsigned(1673, 12), 625 => to_unsigned(2462, 12), 626 => to_unsigned(2447, 12), 627 => to_unsigned(640, 12), 628 => to_unsigned(1487, 12), 629 => to_unsigned(4007, 12), 630 => to_unsigned(2330, 12), 631 => to_unsigned(3645, 12), 632 => to_unsigned(3544, 12), 633 => to_unsigned(3503, 12), 634 => to_unsigned(1341, 12), 635 => to_unsigned(2650, 12), 636 => to_unsigned(2674, 12), 637 => to_unsigned(2, 12), 638 => to_unsigned(1225, 12), 639 => to_unsigned(2425, 12), 640 => to_unsigned(3746, 12), 641 => to_unsigned(800, 12), 642 => to_unsigned(2508, 12), 643 => to_unsigned(1621, 12), 644 => to_unsigned(1602, 12), 645 => to_unsigned(700, 12), 646 => to_unsigned(29, 12), 647 => to_unsigned(1032, 12), 648 => to_unsigned(1108, 12), 649 => to_unsigned(2041, 12), 650 => to_unsigned(2784, 12), 651 => to_unsigned(1081, 12), 652 => to_unsigned(3228, 12), 653 => to_unsigned(3491, 12), 654 => to_unsigned(2304, 12), 655 => to_unsigned(2997, 12), 656 => to_unsigned(3822, 12), 657 => to_unsigned(1267, 12), 658 => to_unsigned(3786, 12), 659 => to_unsigned(1411, 12), 660 => to_unsigned(2158, 12), 661 => to_unsigned(1345, 12), 662 => to_unsigned(1433, 12), 663 => to_unsigned(1420, 12), 664 => to_unsigned(2620, 12), 665 => to_unsigned(2122, 12), 666 => to_unsigned(697, 12), 667 => to_unsigned(2544, 12), 668 => to_unsigned(3478, 12), 669 => to_unsigned(1901, 12), 670 => to_unsigned(3805, 12), 671 => to_unsigned(2634, 12), 672 => to_unsigned(3387, 12), 673 => to_unsigned(1080, 12), 674 => to_unsigned(1074, 12), 675 => to_unsigned(1135, 12), 676 => to_unsigned(3651, 12), 677 => to_unsigned(3831, 12), 678 => to_unsigned(288, 12), 679 => to_unsigned(1828, 12), 680 => to_unsigned(2505, 12), 681 => to_unsigned(3187, 12), 682 => to_unsigned(1249, 12), 683 => to_unsigned(1315, 12), 684 => to_unsigned(1513, 12), 685 => to_unsigned(517, 12), 686 => to_unsigned(222, 12), 687 => to_unsigned(171, 12), 688 => to_unsigned(97, 12), 689 => to_unsigned(3013, 12), 690 => to_unsigned(2332, 12), 691 => to_unsigned(3465, 12), 692 => to_unsigned(2149, 12), 693 => to_unsigned(1790, 12), 694 => to_unsigned(3947, 12), 695 => to_unsigned(829, 12), 696 => to_unsigned(3181, 12), 697 => to_unsigned(94, 12), 698 => to_unsigned(1503, 12), 699 => to_unsigned(3129, 12), 700 => to_unsigned(3521, 12), 701 => to_unsigned(3218, 12), 702 => to_unsigned(766, 12), 703 => to_unsigned(3255, 12), 704 => to_unsigned(3011, 12), 705 => to_unsigned(2949, 12), 706 => to_unsigned(2769, 12), 707 => to_unsigned(166, 12), 708 => to_unsigned(155, 12), 709 => to_unsigned(1770, 12), 710 => to_unsigned(3335, 12), 711 => to_unsigned(3319, 12), 712 => to_unsigned(1515, 12), 713 => to_unsigned(1771, 12), 714 => to_unsigned(1142, 12), 715 => to_unsigned(1723, 12), 716 => to_unsigned(872, 12), 717 => to_unsigned(991, 12), 718 => to_unsigned(2809, 12), 719 => to_unsigned(2294, 12), 720 => to_unsigned(3296, 12), 721 => to_unsigned(865, 12), 722 => to_unsigned(3817, 12), 723 => to_unsigned(730, 12), 724 => to_unsigned(3760, 12), 725 => to_unsigned(1694, 12), 726 => to_unsigned(88, 12), 727 => to_unsigned(359, 12), 728 => to_unsigned(1580, 12), 729 => to_unsigned(698, 12), 730 => to_unsigned(437, 12), 731 => to_unsigned(2897, 12), 732 => to_unsigned(3793, 12), 733 => to_unsigned(556, 12), 734 => to_unsigned(2209, 12), 735 => to_unsigned(2872, 12), 736 => to_unsigned(2693, 12), 737 => to_unsigned(2478, 12), 738 => to_unsigned(2310, 12), 739 => to_unsigned(231, 12), 740 => to_unsigned(2012, 12), 741 => to_unsigned(2196, 12), 742 => to_unsigned(1921, 12), 743 => to_unsigned(721, 12), 744 => to_unsigned(2631, 12), 745 => to_unsigned(548, 12), 746 => to_unsigned(3989, 12), 747 => to_unsigned(360, 12), 748 => to_unsigned(3625, 12), 749 => to_unsigned(2217, 12), 750 => to_unsigned(3988, 12), 751 => to_unsigned(1854, 12), 752 => to_unsigned(2762, 12), 753 => to_unsigned(1543, 12), 754 => to_unsigned(4023, 12), 755 => to_unsigned(2877, 12), 756 => to_unsigned(72, 12), 757 => to_unsigned(2929, 12), 758 => to_unsigned(3029, 12), 759 => to_unsigned(3510, 12), 760 => to_unsigned(1463, 12), 761 => to_unsigned(3734, 12), 762 => to_unsigned(3343, 12), 763 => to_unsigned(1241, 12), 764 => to_unsigned(1450, 12), 765 => to_unsigned(1569, 12), 766 => to_unsigned(3811, 12), 767 => to_unsigned(2214, 12), 768 => to_unsigned(2933, 12), 769 => to_unsigned(1310, 12), 770 => to_unsigned(2924, 12), 771 => to_unsigned(1321, 12), 772 => to_unsigned(2381, 12), 773 => to_unsigned(2518, 12), 774 => to_unsigned(675, 12), 775 => to_unsigned(1609, 12), 776 => to_unsigned(2412, 12), 777 => to_unsigned(4059, 12), 778 => to_unsigned(1787, 12), 779 => to_unsigned(2974, 12), 780 => to_unsigned(3340, 12), 781 => to_unsigned(2110, 12), 782 => to_unsigned(3726, 12), 783 => to_unsigned(482, 12), 784 => to_unsigned(2559, 12), 785 => to_unsigned(2018, 12), 786 => to_unsigned(2764, 12), 787 => to_unsigned(3433, 12), 788 => to_unsigned(624, 12), 789 => to_unsigned(2401, 12), 790 => to_unsigned(1355, 12), 791 => to_unsigned(3320, 12), 792 => to_unsigned(3771, 12), 793 => to_unsigned(2011, 12), 794 => to_unsigned(566, 12), 795 => to_unsigned(1750, 12), 796 => to_unsigned(2916, 12), 797 => to_unsigned(2229, 12), 798 => to_unsigned(3050, 12), 799 => to_unsigned(3895, 12), 800 => to_unsigned(2498, 12), 801 => to_unsigned(3034, 12), 802 => to_unsigned(1090, 12), 803 => to_unsigned(2112, 12), 804 => to_unsigned(2383, 12), 805 => to_unsigned(2618, 12), 806 => to_unsigned(1940, 12), 807 => to_unsigned(2545, 12), 808 => to_unsigned(811, 12), 809 => to_unsigned(3801, 12), 810 => to_unsigned(3983, 12), 811 => to_unsigned(1688, 12), 812 => to_unsigned(3772, 12), 813 => to_unsigned(2563, 12), 814 => to_unsigned(3976, 12), 815 => to_unsigned(3437, 12), 816 => to_unsigned(2324, 12), 817 => to_unsigned(2883, 12), 818 => to_unsigned(1071, 12), 819 => to_unsigned(1582, 12), 820 => to_unsigned(3834, 12), 821 => to_unsigned(3902, 12), 822 => to_unsigned(3987, 12), 823 => to_unsigned(3808, 12), 824 => to_unsigned(2160, 12), 825 => to_unsigned(3757, 12), 826 => to_unsigned(3515, 12), 827 => to_unsigned(444, 12), 828 => to_unsigned(1652, 12), 829 => to_unsigned(3770, 12), 830 => to_unsigned(1542, 12), 831 => to_unsigned(80, 12), 832 => to_unsigned(2674, 12), 833 => to_unsigned(2111, 12), 834 => to_unsigned(882, 12), 835 => to_unsigned(1479, 12), 836 => to_unsigned(1623, 12), 837 => to_unsigned(1428, 12), 838 => to_unsigned(2941, 12), 839 => to_unsigned(962, 12), 840 => to_unsigned(3385, 12), 841 => to_unsigned(3935, 12), 842 => to_unsigned(3610, 12), 843 => to_unsigned(942, 12), 844 => to_unsigned(710, 12), 845 => to_unsigned(2026, 12), 846 => to_unsigned(2253, 12), 847 => to_unsigned(1840, 12), 848 => to_unsigned(2747, 12), 849 => to_unsigned(186, 12), 850 => to_unsigned(2610, 12), 851 => to_unsigned(2398, 12), 852 => to_unsigned(2150, 12), 853 => to_unsigned(1259, 12), 854 => to_unsigned(2616, 12), 855 => to_unsigned(3581, 12), 856 => to_unsigned(357, 12), 857 => to_unsigned(557, 12), 858 => to_unsigned(2864, 12), 859 => to_unsigned(637, 12), 860 => to_unsigned(3297, 12), 861 => to_unsigned(1431, 12), 862 => to_unsigned(68, 12), 863 => to_unsigned(840, 12), 864 => to_unsigned(2832, 12), 865 => to_unsigned(2166, 12), 866 => to_unsigned(3841, 12), 867 => to_unsigned(1203, 12), 868 => to_unsigned(3757, 12), 869 => to_unsigned(1616, 12), 870 => to_unsigned(294, 12), 871 => to_unsigned(2544, 12), 872 => to_unsigned(506, 12), 873 => to_unsigned(1284, 12), 874 => to_unsigned(2675, 12), 875 => to_unsigned(794, 12), 876 => to_unsigned(2796, 12), 877 => to_unsigned(75, 12), 878 => to_unsigned(2821, 12), 879 => to_unsigned(1396, 12), 880 => to_unsigned(3238, 12), 881 => to_unsigned(2539, 12), 882 => to_unsigned(3742, 12), 883 => to_unsigned(24, 12), 884 => to_unsigned(1995, 12), 885 => to_unsigned(3117, 12), 886 => to_unsigned(145, 12), 887 => to_unsigned(3557, 12), 888 => to_unsigned(709, 12), 889 => to_unsigned(1719, 12), 890 => to_unsigned(318, 12), 891 => to_unsigned(3162, 12), 892 => to_unsigned(409, 12), 893 => to_unsigned(3853, 12), 894 => to_unsigned(276, 12), 895 => to_unsigned(2173, 12), 896 => to_unsigned(516, 12), 897 => to_unsigned(2255, 12), 898 => to_unsigned(3065, 12), 899 => to_unsigned(4003, 12), 900 => to_unsigned(1338, 12), 901 => to_unsigned(3261, 12), 902 => to_unsigned(2088, 12), 903 => to_unsigned(3970, 12), 904 => to_unsigned(1991, 12), 905 => to_unsigned(330, 12), 906 => to_unsigned(1371, 12), 907 => to_unsigned(653, 12), 908 => to_unsigned(1420, 12), 909 => to_unsigned(1891, 12), 910 => to_unsigned(3659, 12), 911 => to_unsigned(1728, 12), 912 => to_unsigned(2468, 12), 913 => to_unsigned(670, 12), 914 => to_unsigned(3206, 12), 915 => to_unsigned(1789, 12), 916 => to_unsigned(991, 12), 917 => to_unsigned(1916, 12), 918 => to_unsigned(3184, 12), 919 => to_unsigned(2538, 12), 920 => to_unsigned(383, 12), 921 => to_unsigned(2550, 12), 922 => to_unsigned(2548, 12), 923 => to_unsigned(1511, 12), 924 => to_unsigned(897, 12), 925 => to_unsigned(3729, 12), 926 => to_unsigned(2601, 12), 927 => to_unsigned(3682, 12), 928 => to_unsigned(641, 12), 929 => to_unsigned(2982, 12), 930 => to_unsigned(3408, 12), 931 => to_unsigned(908, 12), 932 => to_unsigned(3136, 12), 933 => to_unsigned(2996, 12), 934 => to_unsigned(214, 12), 935 => to_unsigned(4000, 12), 936 => to_unsigned(4048, 12), 937 => to_unsigned(795, 12), 938 => to_unsigned(2165, 12), 939 => to_unsigned(1954, 12), 940 => to_unsigned(152, 12), 941 => to_unsigned(2274, 12), 942 => to_unsigned(642, 12), 943 => to_unsigned(798, 12), 944 => to_unsigned(1535, 12), 945 => to_unsigned(286, 12), 946 => to_unsigned(837, 12), 947 => to_unsigned(319, 12), 948 => to_unsigned(2555, 12), 949 => to_unsigned(1904, 12), 950 => to_unsigned(2776, 12), 951 => to_unsigned(2950, 12), 952 => to_unsigned(461, 12), 953 => to_unsigned(401, 12), 954 => to_unsigned(1573, 12), 955 => to_unsigned(466, 12), 956 => to_unsigned(3347, 12), 957 => to_unsigned(322, 12), 958 => to_unsigned(2744, 12), 959 => to_unsigned(2455, 12), 960 => to_unsigned(529, 12), 961 => to_unsigned(3424, 12), 962 => to_unsigned(3900, 12), 963 => to_unsigned(545, 12), 964 => to_unsigned(2027, 12), 965 => to_unsigned(2483, 12), 966 => to_unsigned(786, 12), 967 => to_unsigned(3498, 12), 968 => to_unsigned(1633, 12), 969 => to_unsigned(1992, 12), 970 => to_unsigned(809, 12), 971 => to_unsigned(4044, 12), 972 => to_unsigned(2541, 12), 973 => to_unsigned(129, 12), 974 => to_unsigned(989, 12), 975 => to_unsigned(3001, 12), 976 => to_unsigned(1134, 12), 977 => to_unsigned(3069, 12), 978 => to_unsigned(1100, 12), 979 => to_unsigned(3136, 12), 980 => to_unsigned(2364, 12), 981 => to_unsigned(4001, 12), 982 => to_unsigned(1882, 12), 983 => to_unsigned(1579, 12), 984 => to_unsigned(2215, 12), 985 => to_unsigned(3384, 12), 986 => to_unsigned(1246, 12), 987 => to_unsigned(3479, 12), 988 => to_unsigned(1128, 12), 989 => to_unsigned(3862, 12), 990 => to_unsigned(1996, 12), 991 => to_unsigned(3138, 12), 992 => to_unsigned(3545, 12), 993 => to_unsigned(3770, 12), 994 => to_unsigned(1660, 12), 995 => to_unsigned(1168, 12), 996 => to_unsigned(353, 12), 997 => to_unsigned(4052, 12), 998 => to_unsigned(3763, 12), 999 => to_unsigned(955, 12), 1000 => to_unsigned(3187, 12), 1001 => to_unsigned(2638, 12), 1002 => to_unsigned(2949, 12), 1003 => to_unsigned(3807, 12), 1004 => to_unsigned(47, 12), 1005 => to_unsigned(912, 12), 1006 => to_unsigned(896, 12), 1007 => to_unsigned(559, 12), 1008 => to_unsigned(1530, 12), 1009 => to_unsigned(110, 12), 1010 => to_unsigned(22, 12), 1011 => to_unsigned(1490, 12), 1012 => to_unsigned(2019, 12), 1013 => to_unsigned(3100, 12), 1014 => to_unsigned(331, 12), 1015 => to_unsigned(3494, 12), 1016 => to_unsigned(2121, 12), 1017 => to_unsigned(2945, 12), 1018 => to_unsigned(2447, 12), 1019 => to_unsigned(2659, 12), 1020 => to_unsigned(1812, 12), 1021 => to_unsigned(858, 12), 1022 => to_unsigned(3707, 12), 1023 => to_unsigned(172, 12), 1024 => to_unsigned(1420, 12), 1025 => to_unsigned(1263, 12), 1026 => to_unsigned(1641, 12), 1027 => to_unsigned(682, 12), 1028 => to_unsigned(3151, 12), 1029 => to_unsigned(1844, 12), 1030 => to_unsigned(1019, 12), 1031 => to_unsigned(3781, 12), 1032 => to_unsigned(725, 12), 1033 => to_unsigned(796, 12), 1034 => to_unsigned(2342, 12), 1035 => to_unsigned(2439, 12), 1036 => to_unsigned(531, 12), 1037 => to_unsigned(1414, 12), 1038 => to_unsigned(2636, 12), 1039 => to_unsigned(3209, 12), 1040 => to_unsigned(1050, 12), 1041 => to_unsigned(2196, 12), 1042 => to_unsigned(3430, 12), 1043 => to_unsigned(3620, 12), 1044 => to_unsigned(3958, 12), 1045 => to_unsigned(1183, 12), 1046 => to_unsigned(297, 12), 1047 => to_unsigned(212, 12), 1048 => to_unsigned(1680, 12), 1049 => to_unsigned(1440, 12), 1050 => to_unsigned(475, 12), 1051 => to_unsigned(2508, 12), 1052 => to_unsigned(2207, 12), 1053 => to_unsigned(2095, 12), 1054 => to_unsigned(2291, 12), 1055 => to_unsigned(614, 12), 1056 => to_unsigned(3620, 12), 1057 => to_unsigned(2801, 12), 1058 => to_unsigned(151, 12), 1059 => to_unsigned(914, 12), 1060 => to_unsigned(282, 12), 1061 => to_unsigned(307, 12), 1062 => to_unsigned(3632, 12), 1063 => to_unsigned(511, 12), 1064 => to_unsigned(845, 12), 1065 => to_unsigned(1141, 12), 1066 => to_unsigned(1694, 12), 1067 => to_unsigned(3191, 12), 1068 => to_unsigned(3444, 12), 1069 => to_unsigned(2127, 12), 1070 => to_unsigned(3778, 12), 1071 => to_unsigned(3915, 12), 1072 => to_unsigned(2436, 12), 1073 => to_unsigned(1991, 12), 1074 => to_unsigned(465, 12), 1075 => to_unsigned(4051, 12), 1076 => to_unsigned(576, 12), 1077 => to_unsigned(2204, 12), 1078 => to_unsigned(740, 12), 1079 => to_unsigned(2487, 12), 1080 => to_unsigned(3175, 12), 1081 => to_unsigned(1342, 12), 1082 => to_unsigned(2286, 12), 1083 => to_unsigned(1722, 12), 1084 => to_unsigned(463, 12), 1085 => to_unsigned(2274, 12), 1086 => to_unsigned(326, 12), 1087 => to_unsigned(3629, 12), 1088 => to_unsigned(2211, 12), 1089 => to_unsigned(1589, 12), 1090 => to_unsigned(392, 12), 1091 => to_unsigned(3277, 12), 1092 => to_unsigned(2447, 12), 1093 => to_unsigned(3791, 12), 1094 => to_unsigned(3826, 12), 1095 => to_unsigned(2284, 12), 1096 => to_unsigned(2557, 12), 1097 => to_unsigned(3803, 12), 1098 => to_unsigned(1939, 12), 1099 => to_unsigned(448, 12), 1100 => to_unsigned(842, 12), 1101 => to_unsigned(2314, 12), 1102 => to_unsigned(4021, 12), 1103 => to_unsigned(2542, 12), 1104 => to_unsigned(1504, 12), 1105 => to_unsigned(3972, 12), 1106 => to_unsigned(3267, 12), 1107 => to_unsigned(680, 12), 1108 => to_unsigned(3977, 12), 1109 => to_unsigned(311, 12), 1110 => to_unsigned(896, 12), 1111 => to_unsigned(803, 12), 1112 => to_unsigned(2716, 12), 1113 => to_unsigned(2398, 12), 1114 => to_unsigned(2745, 12), 1115 => to_unsigned(81, 12), 1116 => to_unsigned(2117, 12), 1117 => to_unsigned(3809, 12), 1118 => to_unsigned(886, 12), 1119 => to_unsigned(1259, 12), 1120 => to_unsigned(813, 12), 1121 => to_unsigned(3333, 12), 1122 => to_unsigned(792, 12), 1123 => to_unsigned(751, 12), 1124 => to_unsigned(469, 12), 1125 => to_unsigned(525, 12), 1126 => to_unsigned(1535, 12), 1127 => to_unsigned(3735, 12), 1128 => to_unsigned(2978, 12), 1129 => to_unsigned(349, 12), 1130 => to_unsigned(971, 12), 1131 => to_unsigned(1227, 12), 1132 => to_unsigned(4053, 12), 1133 => to_unsigned(475, 12), 1134 => to_unsigned(954, 12), 1135 => to_unsigned(3582, 12), 1136 => to_unsigned(685, 12), 1137 => to_unsigned(2283, 12), 1138 => to_unsigned(2242, 12), 1139 => to_unsigned(1449, 12), 1140 => to_unsigned(3591, 12), 1141 => to_unsigned(2703, 12), 1142 => to_unsigned(3456, 12), 1143 => to_unsigned(1502, 12), 1144 => to_unsigned(3503, 12), 1145 => to_unsigned(123, 12), 1146 => to_unsigned(1066, 12), 1147 => to_unsigned(2790, 12), 1148 => to_unsigned(241, 12), 1149 => to_unsigned(1356, 12), 1150 => to_unsigned(464, 12), 1151 => to_unsigned(3229, 12), 1152 => to_unsigned(3927, 12), 1153 => to_unsigned(1863, 12), 1154 => to_unsigned(1646, 12), 1155 => to_unsigned(2884, 12), 1156 => to_unsigned(543, 12), 1157 => to_unsigned(2208, 12), 1158 => to_unsigned(3971, 12), 1159 => to_unsigned(1125, 12), 1160 => to_unsigned(3470, 12), 1161 => to_unsigned(2370, 12), 1162 => to_unsigned(2064, 12), 1163 => to_unsigned(3231, 12), 1164 => to_unsigned(1150, 12), 1165 => to_unsigned(2163, 12), 1166 => to_unsigned(3095, 12), 1167 => to_unsigned(3801, 12), 1168 => to_unsigned(1307, 12), 1169 => to_unsigned(733, 12), 1170 => to_unsigned(1303, 12), 1171 => to_unsigned(844, 12), 1172 => to_unsigned(2789, 12), 1173 => to_unsigned(808, 12), 1174 => to_unsigned(999, 12), 1175 => to_unsigned(2482, 12), 1176 => to_unsigned(2316, 12), 1177 => to_unsigned(2361, 12), 1178 => to_unsigned(3747, 12), 1179 => to_unsigned(2752, 12), 1180 => to_unsigned(2398, 12), 1181 => to_unsigned(2577, 12), 1182 => to_unsigned(2034, 12), 1183 => to_unsigned(1079, 12), 1184 => to_unsigned(3356, 12), 1185 => to_unsigned(3248, 12), 1186 => to_unsigned(3913, 12), 1187 => to_unsigned(1154, 12), 1188 => to_unsigned(3875, 12), 1189 => to_unsigned(778, 12), 1190 => to_unsigned(924, 12), 1191 => to_unsigned(553, 12), 1192 => to_unsigned(1410, 12), 1193 => to_unsigned(2120, 12), 1194 => to_unsigned(2156, 12), 1195 => to_unsigned(3024, 12), 1196 => to_unsigned(26, 12), 1197 => to_unsigned(1234, 12), 1198 => to_unsigned(2020, 12), 1199 => to_unsigned(2708, 12), 1200 => to_unsigned(443, 12), 1201 => to_unsigned(3562, 12), 1202 => to_unsigned(3533, 12), 1203 => to_unsigned(3085, 12), 1204 => to_unsigned(1038, 12), 1205 => to_unsigned(4090, 12), 1206 => to_unsigned(480, 12), 1207 => to_unsigned(2997, 12), 1208 => to_unsigned(3211, 12), 1209 => to_unsigned(1391, 12), 1210 => to_unsigned(3888, 12), 1211 => to_unsigned(2234, 12), 1212 => to_unsigned(1288, 12), 1213 => to_unsigned(1521, 12), 1214 => to_unsigned(2540, 12), 1215 => to_unsigned(3112, 12), 1216 => to_unsigned(2096, 12), 1217 => to_unsigned(2210, 12), 1218 => to_unsigned(165, 12), 1219 => to_unsigned(2915, 12), 1220 => to_unsigned(621, 12), 1221 => to_unsigned(2856, 12), 1222 => to_unsigned(3705, 12), 1223 => to_unsigned(522, 12), 1224 => to_unsigned(3119, 12), 1225 => to_unsigned(3963, 12), 1226 => to_unsigned(535, 12), 1227 => to_unsigned(2104, 12), 1228 => to_unsigned(1702, 12), 1229 => to_unsigned(132, 12), 1230 => to_unsigned(948, 12), 1231 => to_unsigned(2878, 12), 1232 => to_unsigned(1020, 12), 1233 => to_unsigned(3063, 12), 1234 => to_unsigned(2735, 12), 1235 => to_unsigned(2842, 12), 1236 => to_unsigned(3783, 12), 1237 => to_unsigned(2292, 12), 1238 => to_unsigned(2291, 12), 1239 => to_unsigned(3162, 12), 1240 => to_unsigned(2073, 12), 1241 => to_unsigned(1321, 12), 1242 => to_unsigned(20, 12), 1243 => to_unsigned(3069, 12), 1244 => to_unsigned(1183, 12), 1245 => to_unsigned(3438, 12), 1246 => to_unsigned(2807, 12), 1247 => to_unsigned(182, 12), 1248 => to_unsigned(2178, 12), 1249 => to_unsigned(446, 12), 1250 => to_unsigned(2871, 12), 1251 => to_unsigned(3716, 12), 1252 => to_unsigned(4062, 12), 1253 => to_unsigned(3612, 12), 1254 => to_unsigned(2317, 12), 1255 => to_unsigned(25, 12), 1256 => to_unsigned(2909, 12), 1257 => to_unsigned(2161, 12), 1258 => to_unsigned(3154, 12), 1259 => to_unsigned(3606, 12), 1260 => to_unsigned(3972, 12), 1261 => to_unsigned(1458, 12), 1262 => to_unsigned(2423, 12), 1263 => to_unsigned(3963, 12), 1264 => to_unsigned(2547, 12), 1265 => to_unsigned(1133, 12), 1266 => to_unsigned(3424, 12), 1267 => to_unsigned(3623, 12), 1268 => to_unsigned(1681, 12), 1269 => to_unsigned(3650, 12), 1270 => to_unsigned(3036, 12), 1271 => to_unsigned(1336, 12), 1272 => to_unsigned(1691, 12), 1273 => to_unsigned(3150, 12), 1274 => to_unsigned(1364, 12), 1275 => to_unsigned(3232, 12), 1276 => to_unsigned(631, 12), 1277 => to_unsigned(3224, 12), 1278 => to_unsigned(3403, 12), 1279 => to_unsigned(2126, 12), 1280 => to_unsigned(3086, 12), 1281 => to_unsigned(4077, 12), 1282 => to_unsigned(1772, 12), 1283 => to_unsigned(1956, 12), 1284 => to_unsigned(1416, 12), 1285 => to_unsigned(1837, 12), 1286 => to_unsigned(1525, 12), 1287 => to_unsigned(2265, 12), 1288 => to_unsigned(3953, 12), 1289 => to_unsigned(1457, 12), 1290 => to_unsigned(2135, 12), 1291 => to_unsigned(1960, 12), 1292 => to_unsigned(2313, 12), 1293 => to_unsigned(3891, 12), 1294 => to_unsigned(2664, 12), 1295 => to_unsigned(2989, 12), 1296 => to_unsigned(473, 12), 1297 => to_unsigned(62, 12), 1298 => to_unsigned(1034, 12), 1299 => to_unsigned(2548, 12), 1300 => to_unsigned(2127, 12), 1301 => to_unsigned(4072, 12), 1302 => to_unsigned(423, 12), 1303 => to_unsigned(1958, 12), 1304 => to_unsigned(2428, 12), 1305 => to_unsigned(1796, 12), 1306 => to_unsigned(767, 12), 1307 => to_unsigned(1697, 12), 1308 => to_unsigned(1226, 12), 1309 => to_unsigned(3961, 12), 1310 => to_unsigned(1589, 12), 1311 => to_unsigned(162, 12), 1312 => to_unsigned(1346, 12), 1313 => to_unsigned(3247, 12), 1314 => to_unsigned(1853, 12), 1315 => to_unsigned(3524, 12), 1316 => to_unsigned(484, 12), 1317 => to_unsigned(418, 12), 1318 => to_unsigned(2037, 12), 1319 => to_unsigned(34, 12), 1320 => to_unsigned(274, 12), 1321 => to_unsigned(1388, 12), 1322 => to_unsigned(2565, 12), 1323 => to_unsigned(1013, 12), 1324 => to_unsigned(283, 12), 1325 => to_unsigned(1171, 12), 1326 => to_unsigned(2165, 12), 1327 => to_unsigned(3152, 12), 1328 => to_unsigned(611, 12), 1329 => to_unsigned(1833, 12), 1330 => to_unsigned(1446, 12), 1331 => to_unsigned(4060, 12), 1332 => to_unsigned(1675, 12), 1333 => to_unsigned(3450, 12), 1334 => to_unsigned(2287, 12), 1335 => to_unsigned(3066, 12), 1336 => to_unsigned(2361, 12), 1337 => to_unsigned(1472, 12), 1338 => to_unsigned(3474, 12), 1339 => to_unsigned(1317, 12), 1340 => to_unsigned(1574, 12), 1341 => to_unsigned(3854, 12), 1342 => to_unsigned(3787, 12), 1343 => to_unsigned(4005, 12), 1344 => to_unsigned(1802, 12), 1345 => to_unsigned(2775, 12), 1346 => to_unsigned(1159, 12), 1347 => to_unsigned(1239, 12), 1348 => to_unsigned(3160, 12), 1349 => to_unsigned(3217, 12), 1350 => to_unsigned(1808, 12), 1351 => to_unsigned(120, 12), 1352 => to_unsigned(2844, 12), 1353 => to_unsigned(2418, 12), 1354 => to_unsigned(3511, 12), 1355 => to_unsigned(21, 12), 1356 => to_unsigned(2770, 12), 1357 => to_unsigned(1547, 12), 1358 => to_unsigned(2264, 12), 1359 => to_unsigned(2137, 12), 1360 => to_unsigned(346, 12), 1361 => to_unsigned(2278, 12), 1362 => to_unsigned(1006, 12), 1363 => to_unsigned(1039, 12), 1364 => to_unsigned(1914, 12), 1365 => to_unsigned(2551, 12), 1366 => to_unsigned(3877, 12), 1367 => to_unsigned(609, 12), 1368 => to_unsigned(3093, 12), 1369 => to_unsigned(2125, 12), 1370 => to_unsigned(1630, 12), 1371 => to_unsigned(2132, 12), 1372 => to_unsigned(990, 12), 1373 => to_unsigned(2715, 12), 1374 => to_unsigned(1762, 12), 1375 => to_unsigned(1629, 12), 1376 => to_unsigned(1538, 12), 1377 => to_unsigned(1419, 12), 1378 => to_unsigned(3035, 12), 1379 => to_unsigned(1314, 12), 1380 => to_unsigned(1910, 12), 1381 => to_unsigned(3963, 12), 1382 => to_unsigned(1019, 12), 1383 => to_unsigned(321, 12), 1384 => to_unsigned(3315, 12), 1385 => to_unsigned(3145, 12), 1386 => to_unsigned(86, 12), 1387 => to_unsigned(407, 12), 1388 => to_unsigned(3416, 12), 1389 => to_unsigned(323, 12), 1390 => to_unsigned(2237, 12), 1391 => to_unsigned(1633, 12), 1392 => to_unsigned(3928, 12), 1393 => to_unsigned(1919, 12), 1394 => to_unsigned(3227, 12), 1395 => to_unsigned(1395, 12), 1396 => to_unsigned(2508, 12), 1397 => to_unsigned(3070, 12), 1398 => to_unsigned(1127, 12), 1399 => to_unsigned(2138, 12), 1400 => to_unsigned(1125, 12), 1401 => to_unsigned(3700, 12), 1402 => to_unsigned(1183, 12), 1403 => to_unsigned(3878, 12), 1404 => to_unsigned(3643, 12), 1405 => to_unsigned(156, 12), 1406 => to_unsigned(420, 12), 1407 => to_unsigned(979, 12), 1408 => to_unsigned(2501, 12), 1409 => to_unsigned(2991, 12), 1410 => to_unsigned(1671, 12), 1411 => to_unsigned(3855, 12), 1412 => to_unsigned(546, 12), 1413 => to_unsigned(141, 12), 1414 => to_unsigned(2136, 12), 1415 => to_unsigned(1717, 12), 1416 => to_unsigned(759, 12), 1417 => to_unsigned(367, 12), 1418 => to_unsigned(171, 12), 1419 => to_unsigned(2515, 12), 1420 => to_unsigned(3129, 12), 1421 => to_unsigned(2480, 12), 1422 => to_unsigned(2443, 12), 1423 => to_unsigned(3810, 12), 1424 => to_unsigned(1112, 12), 1425 => to_unsigned(661, 12), 1426 => to_unsigned(3953, 12), 1427 => to_unsigned(470, 12), 1428 => to_unsigned(3000, 12), 1429 => to_unsigned(481, 12), 1430 => to_unsigned(1779, 12), 1431 => to_unsigned(1063, 12), 1432 => to_unsigned(1707, 12), 1433 => to_unsigned(1888, 12), 1434 => to_unsigned(2450, 12), 1435 => to_unsigned(1148, 12), 1436 => to_unsigned(1168, 12), 1437 => to_unsigned(3077, 12), 1438 => to_unsigned(2463, 12), 1439 => to_unsigned(1044, 12), 1440 => to_unsigned(283, 12), 1441 => to_unsigned(3050, 12), 1442 => to_unsigned(2261, 12), 1443 => to_unsigned(2758, 12), 1444 => to_unsigned(1815, 12), 1445 => to_unsigned(2800, 12), 1446 => to_unsigned(743, 12), 1447 => to_unsigned(1719, 12), 1448 => to_unsigned(3615, 12), 1449 => to_unsigned(2100, 12), 1450 => to_unsigned(1661, 12), 1451 => to_unsigned(2952, 12), 1452 => to_unsigned(824, 12), 1453 => to_unsigned(2218, 12), 1454 => to_unsigned(756, 12), 1455 => to_unsigned(4095, 12), 1456 => to_unsigned(3811, 12), 1457 => to_unsigned(1755, 12), 1458 => to_unsigned(1763, 12), 1459 => to_unsigned(1793, 12), 1460 => to_unsigned(633, 12), 1461 => to_unsigned(1318, 12), 1462 => to_unsigned(2530, 12), 1463 => to_unsigned(3548, 12), 1464 => to_unsigned(2532, 12), 1465 => to_unsigned(2710, 12), 1466 => to_unsigned(3977, 12), 1467 => to_unsigned(3231, 12), 1468 => to_unsigned(2926, 12), 1469 => to_unsigned(3961, 12), 1470 => to_unsigned(89, 12), 1471 => to_unsigned(3330, 12), 1472 => to_unsigned(3205, 12), 1473 => to_unsigned(2783, 12), 1474 => to_unsigned(3229, 12), 1475 => to_unsigned(2920, 12), 1476 => to_unsigned(472, 12), 1477 => to_unsigned(2549, 12), 1478 => to_unsigned(944, 12), 1479 => to_unsigned(2014, 12), 1480 => to_unsigned(1364, 12), 1481 => to_unsigned(205, 12), 1482 => to_unsigned(440, 12), 1483 => to_unsigned(2530, 12), 1484 => to_unsigned(1689, 12), 1485 => to_unsigned(3116, 12), 1486 => to_unsigned(2949, 12), 1487 => to_unsigned(3808, 12), 1488 => to_unsigned(3689, 12), 1489 => to_unsigned(3460, 12), 1490 => to_unsigned(3875, 12), 1491 => to_unsigned(2135, 12), 1492 => to_unsigned(2538, 12), 1493 => to_unsigned(3962, 12), 1494 => to_unsigned(1026, 12), 1495 => to_unsigned(1362, 12), 1496 => to_unsigned(1802, 12), 1497 => to_unsigned(2736, 12), 1498 => to_unsigned(816, 12), 1499 => to_unsigned(3611, 12), 1500 => to_unsigned(3100, 12), 1501 => to_unsigned(120, 12), 1502 => to_unsigned(470, 12), 1503 => to_unsigned(2546, 12), 1504 => to_unsigned(3685, 12), 1505 => to_unsigned(3297, 12), 1506 => to_unsigned(1655, 12), 1507 => to_unsigned(3721, 12), 1508 => to_unsigned(3950, 12), 1509 => to_unsigned(1812, 12), 1510 => to_unsigned(1003, 12), 1511 => to_unsigned(1435, 12), 1512 => to_unsigned(3056, 12), 1513 => to_unsigned(483, 12), 1514 => to_unsigned(5, 12), 1515 => to_unsigned(219, 12), 1516 => to_unsigned(1462, 12), 1517 => to_unsigned(3786, 12), 1518 => to_unsigned(229, 12), 1519 => to_unsigned(1957, 12), 1520 => to_unsigned(1953, 12), 1521 => to_unsigned(496, 12), 1522 => to_unsigned(791, 12), 1523 => to_unsigned(3571, 12), 1524 => to_unsigned(2403, 12), 1525 => to_unsigned(2097, 12), 1526 => to_unsigned(2404, 12), 1527 => to_unsigned(1086, 12), 1528 => to_unsigned(2504, 12), 1529 => to_unsigned(3445, 12), 1530 => to_unsigned(2571, 12), 1531 => to_unsigned(2296, 12), 1532 => to_unsigned(3574, 12), 1533 => to_unsigned(2381, 12), 1534 => to_unsigned(2807, 12), 1535 => to_unsigned(3085, 12), 1536 => to_unsigned(1774, 12), 1537 => to_unsigned(2965, 12), 1538 => to_unsigned(223, 12), 1539 => to_unsigned(2448, 12), 1540 => to_unsigned(2868, 12), 1541 => to_unsigned(1406, 12), 1542 => to_unsigned(835, 12), 1543 => to_unsigned(1325, 12), 1544 => to_unsigned(3672, 12), 1545 => to_unsigned(1515, 12), 1546 => to_unsigned(2341, 12), 1547 => to_unsigned(2678, 12), 1548 => to_unsigned(2389, 12), 1549 => to_unsigned(3797, 12), 1550 => to_unsigned(1803, 12), 1551 => to_unsigned(3626, 12), 1552 => to_unsigned(2300, 12), 1553 => to_unsigned(2863, 12), 1554 => to_unsigned(3760, 12), 1555 => to_unsigned(1037, 12), 1556 => to_unsigned(1184, 12), 1557 => to_unsigned(711, 12), 1558 => to_unsigned(3275, 12), 1559 => to_unsigned(3303, 12), 1560 => to_unsigned(872, 12), 1561 => to_unsigned(1986, 12), 1562 => to_unsigned(1710, 12), 1563 => to_unsigned(74, 12), 1564 => to_unsigned(1969, 12), 1565 => to_unsigned(1623, 12), 1566 => to_unsigned(2399, 12), 1567 => to_unsigned(3622, 12), 1568 => to_unsigned(672, 12), 1569 => to_unsigned(3119, 12), 1570 => to_unsigned(3166, 12), 1571 => to_unsigned(2496, 12), 1572 => to_unsigned(3958, 12), 1573 => to_unsigned(821, 12), 1574 => to_unsigned(3788, 12), 1575 => to_unsigned(2965, 12), 1576 => to_unsigned(3723, 12), 1577 => to_unsigned(2332, 12), 1578 => to_unsigned(3402, 12), 1579 => to_unsigned(3351, 12), 1580 => to_unsigned(2061, 12), 1581 => to_unsigned(3328, 12), 1582 => to_unsigned(525, 12), 1583 => to_unsigned(1680, 12), 1584 => to_unsigned(2588, 12), 1585 => to_unsigned(2581, 12), 1586 => to_unsigned(3916, 12), 1587 => to_unsigned(421, 12), 1588 => to_unsigned(2129, 12), 1589 => to_unsigned(2277, 12), 1590 => to_unsigned(2593, 12), 1591 => to_unsigned(1326, 12), 1592 => to_unsigned(709, 12), 1593 => to_unsigned(73, 12), 1594 => to_unsigned(3927, 12), 1595 => to_unsigned(468, 12), 1596 => to_unsigned(347, 12), 1597 => to_unsigned(1117, 12), 1598 => to_unsigned(599, 12), 1599 => to_unsigned(412, 12), 1600 => to_unsigned(4093, 12), 1601 => to_unsigned(1314, 12), 1602 => to_unsigned(2048, 12), 1603 => to_unsigned(787, 12), 1604 => to_unsigned(1576, 12), 1605 => to_unsigned(923, 12), 1606 => to_unsigned(1579, 12), 1607 => to_unsigned(866, 12), 1608 => to_unsigned(1965, 12), 1609 => to_unsigned(2254, 12), 1610 => to_unsigned(1690, 12), 1611 => to_unsigned(3698, 12), 1612 => to_unsigned(1936, 12), 1613 => to_unsigned(1562, 12), 1614 => to_unsigned(643, 12), 1615 => to_unsigned(544, 12), 1616 => to_unsigned(1223, 12), 1617 => to_unsigned(1571, 12), 1618 => to_unsigned(2743, 12), 1619 => to_unsigned(1249, 12), 1620 => to_unsigned(629, 12), 1621 => to_unsigned(1397, 12), 1622 => to_unsigned(2519, 12), 1623 => to_unsigned(688, 12), 1624 => to_unsigned(3171, 12), 1625 => to_unsigned(2499, 12), 1626 => to_unsigned(3494, 12), 1627 => to_unsigned(1728, 12), 1628 => to_unsigned(433, 12), 1629 => to_unsigned(2487, 12), 1630 => to_unsigned(3686, 12), 1631 => to_unsigned(3112, 12), 1632 => to_unsigned(2682, 12), 1633 => to_unsigned(711, 12), 1634 => to_unsigned(2970, 12), 1635 => to_unsigned(2962, 12), 1636 => to_unsigned(652, 12), 1637 => to_unsigned(1030, 12), 1638 => to_unsigned(1249, 12), 1639 => to_unsigned(648, 12), 1640 => to_unsigned(3108, 12), 1641 => to_unsigned(4057, 12), 1642 => to_unsigned(517, 12), 1643 => to_unsigned(4059, 12), 1644 => to_unsigned(1304, 12), 1645 => to_unsigned(1362, 12), 1646 => to_unsigned(3897, 12), 1647 => to_unsigned(3835, 12), 1648 => to_unsigned(287, 12), 1649 => to_unsigned(97, 12), 1650 => to_unsigned(1715, 12), 1651 => to_unsigned(2785, 12), 1652 => to_unsigned(666, 12), 1653 => to_unsigned(3423, 12), 1654 => to_unsigned(3086, 12), 1655 => to_unsigned(12, 12), 1656 => to_unsigned(1406, 12), 1657 => to_unsigned(803, 12), 1658 => to_unsigned(2840, 12), 1659 => to_unsigned(3656, 12), 1660 => to_unsigned(3191, 12), 1661 => to_unsigned(2441, 12), 1662 => to_unsigned(1204, 12), 1663 => to_unsigned(3687, 12), 1664 => to_unsigned(1355, 12), 1665 => to_unsigned(4044, 12), 1666 => to_unsigned(913, 12), 1667 => to_unsigned(1891, 12), 1668 => to_unsigned(864, 12), 1669 => to_unsigned(896, 12), 1670 => to_unsigned(2798, 12), 1671 => to_unsigned(1291, 12), 1672 => to_unsigned(2771, 12), 1673 => to_unsigned(1723, 12), 1674 => to_unsigned(3672, 12), 1675 => to_unsigned(1931, 12), 1676 => to_unsigned(766, 12), 1677 => to_unsigned(1907, 12), 1678 => to_unsigned(860, 12), 1679 => to_unsigned(849, 12), 1680 => to_unsigned(2692, 12), 1681 => to_unsigned(697, 12), 1682 => to_unsigned(3350, 12), 1683 => to_unsigned(3670, 12), 1684 => to_unsigned(2230, 12), 1685 => to_unsigned(1025, 12), 1686 => to_unsigned(2797, 12), 1687 => to_unsigned(129, 12), 1688 => to_unsigned(136, 12), 1689 => to_unsigned(1303, 12), 1690 => to_unsigned(2927, 12), 1691 => to_unsigned(3920, 12), 1692 => to_unsigned(2406, 12), 1693 => to_unsigned(3798, 12), 1694 => to_unsigned(4043, 12), 1695 => to_unsigned(3519, 12), 1696 => to_unsigned(236, 12), 1697 => to_unsigned(1116, 12), 1698 => to_unsigned(1955, 12), 1699 => to_unsigned(2508, 12), 1700 => to_unsigned(2371, 12), 1701 => to_unsigned(3050, 12), 1702 => to_unsigned(3532, 12), 1703 => to_unsigned(3000, 12), 1704 => to_unsigned(2306, 12), 1705 => to_unsigned(2059, 12), 1706 => to_unsigned(1224, 12), 1707 => to_unsigned(3708, 12), 1708 => to_unsigned(4033, 12), 1709 => to_unsigned(2195, 12), 1710 => to_unsigned(3044, 12), 1711 => to_unsigned(3188, 12), 1712 => to_unsigned(926, 12), 1713 => to_unsigned(2899, 12), 1714 => to_unsigned(147, 12), 1715 => to_unsigned(867, 12), 1716 => to_unsigned(3956, 12), 1717 => to_unsigned(1479, 12), 1718 => to_unsigned(2442, 12), 1719 => to_unsigned(1517, 12), 1720 => to_unsigned(3449, 12), 1721 => to_unsigned(2076, 12), 1722 => to_unsigned(2851, 12), 1723 => to_unsigned(1714, 12), 1724 => to_unsigned(2927, 12), 1725 => to_unsigned(689, 12), 1726 => to_unsigned(2994, 12), 1727 => to_unsigned(1155, 12), 1728 => to_unsigned(3401, 12), 1729 => to_unsigned(2666, 12), 1730 => to_unsigned(82, 12), 1731 => to_unsigned(3711, 12), 1732 => to_unsigned(1462, 12), 1733 => to_unsigned(1093, 12), 1734 => to_unsigned(3994, 12), 1735 => to_unsigned(3261, 12), 1736 => to_unsigned(2999, 12), 1737 => to_unsigned(1871, 12), 1738 => to_unsigned(1917, 12), 1739 => to_unsigned(2710, 12), 1740 => to_unsigned(375, 12), 1741 => to_unsigned(269, 12), 1742 => to_unsigned(3326, 12), 1743 => to_unsigned(1745, 12), 1744 => to_unsigned(43, 12), 1745 => to_unsigned(825, 12), 1746 => to_unsigned(4002, 12), 1747 => to_unsigned(3854, 12), 1748 => to_unsigned(2570, 12), 1749 => to_unsigned(835, 12), 1750 => to_unsigned(328, 12), 1751 => to_unsigned(987, 12), 1752 => to_unsigned(3137, 12), 1753 => to_unsigned(2919, 12), 1754 => to_unsigned(690, 12), 1755 => to_unsigned(492, 12), 1756 => to_unsigned(2706, 12), 1757 => to_unsigned(695, 12), 1758 => to_unsigned(3070, 12), 1759 => to_unsigned(328, 12), 1760 => to_unsigned(2048, 12), 1761 => to_unsigned(2291, 12), 1762 => to_unsigned(3404, 12), 1763 => to_unsigned(3453, 12), 1764 => to_unsigned(3199, 12), 1765 => to_unsigned(3497, 12), 1766 => to_unsigned(1739, 12), 1767 => to_unsigned(2186, 12), 1768 => to_unsigned(3116, 12), 1769 => to_unsigned(618, 12), 1770 => to_unsigned(2054, 12), 1771 => to_unsigned(2262, 12), 1772 => to_unsigned(4076, 12), 1773 => to_unsigned(3527, 12), 1774 => to_unsigned(1548, 12), 1775 => to_unsigned(1876, 12), 1776 => to_unsigned(553, 12), 1777 => to_unsigned(1629, 12), 1778 => to_unsigned(356, 12), 1779 => to_unsigned(387, 12), 1780 => to_unsigned(376, 12), 1781 => to_unsigned(2924, 12), 1782 => to_unsigned(775, 12), 1783 => to_unsigned(1485, 12), 1784 => to_unsigned(3385, 12), 1785 => to_unsigned(2706, 12), 1786 => to_unsigned(444, 12), 1787 => to_unsigned(1624, 12), 1788 => to_unsigned(3065, 12), 1789 => to_unsigned(3297, 12), 1790 => to_unsigned(2146, 12), 1791 => to_unsigned(2924, 12), 1792 => to_unsigned(3541, 12), 1793 => to_unsigned(2083, 12), 1794 => to_unsigned(1628, 12), 1795 => to_unsigned(241, 12), 1796 => to_unsigned(3455, 12), 1797 => to_unsigned(1638, 12), 1798 => to_unsigned(236, 12), 1799 => to_unsigned(3867, 12), 1800 => to_unsigned(2654, 12), 1801 => to_unsigned(1755, 12), 1802 => to_unsigned(2881, 12), 1803 => to_unsigned(2056, 12), 1804 => to_unsigned(3957, 12), 1805 => to_unsigned(2905, 12), 1806 => to_unsigned(1309, 12), 1807 => to_unsigned(3727, 12), 1808 => to_unsigned(2307, 12), 1809 => to_unsigned(435, 12), 1810 => to_unsigned(2711, 12), 1811 => to_unsigned(863, 12), 1812 => to_unsigned(1910, 12), 1813 => to_unsigned(1252, 12), 1814 => to_unsigned(1045, 12), 1815 => to_unsigned(341, 12), 1816 => to_unsigned(3010, 12), 1817 => to_unsigned(371, 12), 1818 => to_unsigned(4063, 12), 1819 => to_unsigned(3272, 12), 1820 => to_unsigned(1733, 12), 1821 => to_unsigned(2489, 12), 1822 => to_unsigned(2611, 12), 1823 => to_unsigned(3596, 12), 1824 => to_unsigned(1636, 12), 1825 => to_unsigned(1162, 12), 1826 => to_unsigned(185, 12), 1827 => to_unsigned(870, 12), 1828 => to_unsigned(2235, 12), 1829 => to_unsigned(3378, 12), 1830 => to_unsigned(232, 12), 1831 => to_unsigned(203, 12), 1832 => to_unsigned(3114, 12), 1833 => to_unsigned(2815, 12), 1834 => to_unsigned(413, 12), 1835 => to_unsigned(357, 12), 1836 => to_unsigned(3637, 12), 1837 => to_unsigned(1448, 12), 1838 => to_unsigned(428, 12), 1839 => to_unsigned(3401, 12), 1840 => to_unsigned(3497, 12), 1841 => to_unsigned(1112, 12), 1842 => to_unsigned(2859, 12), 1843 => to_unsigned(2983, 12), 1844 => to_unsigned(3553, 12), 1845 => to_unsigned(3017, 12), 1846 => to_unsigned(3590, 12), 1847 => to_unsigned(600, 12), 1848 => to_unsigned(1687, 12), 1849 => to_unsigned(1832, 12), 1850 => to_unsigned(2565, 12), 1851 => to_unsigned(3726, 12), 1852 => to_unsigned(2044, 12), 1853 => to_unsigned(983, 12), 1854 => to_unsigned(3728, 12), 1855 => to_unsigned(3240, 12), 1856 => to_unsigned(3354, 12), 1857 => to_unsigned(526, 12), 1858 => to_unsigned(2507, 12), 1859 => to_unsigned(2362, 12), 1860 => to_unsigned(719, 12), 1861 => to_unsigned(1768, 12), 1862 => to_unsigned(271, 12), 1863 => to_unsigned(3772, 12), 1864 => to_unsigned(1683, 12), 1865 => to_unsigned(2170, 12), 1866 => to_unsigned(3410, 12), 1867 => to_unsigned(1214, 12), 1868 => to_unsigned(2367, 12), 1869 => to_unsigned(2427, 12), 1870 => to_unsigned(2639, 12), 1871 => to_unsigned(2693, 12), 1872 => to_unsigned(2375, 12), 1873 => to_unsigned(583, 12), 1874 => to_unsigned(918, 12), 1875 => to_unsigned(2608, 12), 1876 => to_unsigned(2899, 12), 1877 => to_unsigned(2830, 12), 1878 => to_unsigned(3842, 12), 1879 => to_unsigned(1017, 12), 1880 => to_unsigned(875, 12), 1881 => to_unsigned(975, 12), 1882 => to_unsigned(916, 12), 1883 => to_unsigned(394, 12), 1884 => to_unsigned(2389, 12), 1885 => to_unsigned(2410, 12), 1886 => to_unsigned(3369, 12), 1887 => to_unsigned(2609, 12), 1888 => to_unsigned(1977, 12), 1889 => to_unsigned(4017, 12), 1890 => to_unsigned(3568, 12), 1891 => to_unsigned(3485, 12), 1892 => to_unsigned(3691, 12), 1893 => to_unsigned(2372, 12), 1894 => to_unsigned(676, 12), 1895 => to_unsigned(2762, 12), 1896 => to_unsigned(3392, 12), 1897 => to_unsigned(3218, 12), 1898 => to_unsigned(1068, 12), 1899 => to_unsigned(387, 12), 1900 => to_unsigned(2608, 12), 1901 => to_unsigned(856, 12), 1902 => to_unsigned(3228, 12), 1903 => to_unsigned(2850, 12), 1904 => to_unsigned(747, 12), 1905 => to_unsigned(2888, 12), 1906 => to_unsigned(3194, 12), 1907 => to_unsigned(1336, 12), 1908 => to_unsigned(805, 12), 1909 => to_unsigned(3306, 12), 1910 => to_unsigned(1759, 12), 1911 => to_unsigned(2409, 12), 1912 => to_unsigned(2930, 12), 1913 => to_unsigned(3980, 12), 1914 => to_unsigned(3371, 12), 1915 => to_unsigned(3366, 12), 1916 => to_unsigned(2736, 12), 1917 => to_unsigned(2522, 12), 1918 => to_unsigned(3844, 12), 1919 => to_unsigned(1958, 12), 1920 => to_unsigned(207, 12), 1921 => to_unsigned(1691, 12), 1922 => to_unsigned(2293, 12), 1923 => to_unsigned(1034, 12), 1924 => to_unsigned(1130, 12), 1925 => to_unsigned(1799, 12), 1926 => to_unsigned(3766, 12), 1927 => to_unsigned(3800, 12), 1928 => to_unsigned(1953, 12), 1929 => to_unsigned(2784, 12), 1930 => to_unsigned(3385, 12), 1931 => to_unsigned(1470, 12), 1932 => to_unsigned(1787, 12), 1933 => to_unsigned(216, 12), 1934 => to_unsigned(3284, 12), 1935 => to_unsigned(3806, 12), 1936 => to_unsigned(3332, 12), 1937 => to_unsigned(2101, 12), 1938 => to_unsigned(908, 12), 1939 => to_unsigned(158, 12), 1940 => to_unsigned(1326, 12), 1941 => to_unsigned(20, 12), 1942 => to_unsigned(1505, 12), 1943 => to_unsigned(1594, 12), 1944 => to_unsigned(1587, 12), 1945 => to_unsigned(3973, 12), 1946 => to_unsigned(1084, 12), 1947 => to_unsigned(2387, 12), 1948 => to_unsigned(2951, 12), 1949 => to_unsigned(430, 12), 1950 => to_unsigned(472, 12), 1951 => to_unsigned(393, 12), 1952 => to_unsigned(1073, 12), 1953 => to_unsigned(1809, 12), 1954 => to_unsigned(866, 12), 1955 => to_unsigned(1934, 12), 1956 => to_unsigned(3266, 12), 1957 => to_unsigned(103, 12), 1958 => to_unsigned(1417, 12), 1959 => to_unsigned(2490, 12), 1960 => to_unsigned(1435, 12), 1961 => to_unsigned(4043, 12), 1962 => to_unsigned(2107, 12), 1963 => to_unsigned(2155, 12), 1964 => to_unsigned(3631, 12), 1965 => to_unsigned(2549, 12), 1966 => to_unsigned(1839, 12), 1967 => to_unsigned(1750, 12), 1968 => to_unsigned(416, 12), 1969 => to_unsigned(1384, 12), 1970 => to_unsigned(3561, 12), 1971 => to_unsigned(1333, 12), 1972 => to_unsigned(388, 12), 1973 => to_unsigned(1565, 12), 1974 => to_unsigned(1189, 12), 1975 => to_unsigned(3114, 12), 1976 => to_unsigned(1250, 12), 1977 => to_unsigned(3311, 12), 1978 => to_unsigned(102, 12), 1979 => to_unsigned(2837, 12), 1980 => to_unsigned(3734, 12), 1981 => to_unsigned(2870, 12), 1982 => to_unsigned(2366, 12), 1983 => to_unsigned(1425, 12), 1984 => to_unsigned(2418, 12), 1985 => to_unsigned(1027, 12), 1986 => to_unsigned(786, 12), 1987 => to_unsigned(4037, 12), 1988 => to_unsigned(1065, 12), 1989 => to_unsigned(3618, 12), 1990 => to_unsigned(649, 12), 1991 => to_unsigned(2162, 12), 1992 => to_unsigned(3443, 12), 1993 => to_unsigned(1884, 12), 1994 => to_unsigned(800, 12), 1995 => to_unsigned(1565, 12), 1996 => to_unsigned(3296, 12), 1997 => to_unsigned(2399, 12), 1998 => to_unsigned(3323, 12), 1999 => to_unsigned(1354, 12), 2000 => to_unsigned(137, 12), 2001 => to_unsigned(2453, 12), 2002 => to_unsigned(317, 12), 2003 => to_unsigned(2618, 12), 2004 => to_unsigned(3767, 12), 2005 => to_unsigned(99, 12), 2006 => to_unsigned(1913, 12), 2007 => to_unsigned(254, 12), 2008 => to_unsigned(1884, 12), 2009 => to_unsigned(905, 12), 2010 => to_unsigned(1456, 12), 2011 => to_unsigned(3370, 12), 2012 => to_unsigned(1372, 12), 2013 => to_unsigned(3653, 12), 2014 => to_unsigned(1860, 12), 2015 => to_unsigned(529, 12), 2016 => to_unsigned(560, 12), 2017 => to_unsigned(3312, 12), 2018 => to_unsigned(3264, 12), 2019 => to_unsigned(1332, 12), 2020 => to_unsigned(889, 12), 2021 => to_unsigned(2820, 12), 2022 => to_unsigned(1200, 12), 2023 => to_unsigned(2943, 12), 2024 => to_unsigned(3976, 12), 2025 => to_unsigned(2279, 12), 2026 => to_unsigned(945, 12), 2027 => to_unsigned(3928, 12), 2028 => to_unsigned(28, 12), 2029 => to_unsigned(1081, 12), 2030 => to_unsigned(3628, 12), 2031 => to_unsigned(731, 12), 2032 => to_unsigned(3947, 12), 2033 => to_unsigned(3750, 12), 2034 => to_unsigned(2116, 12), 2035 => to_unsigned(2650, 12), 2036 => to_unsigned(2200, 12), 2037 => to_unsigned(2123, 12), 2038 => to_unsigned(2348, 12), 2039 => to_unsigned(281, 12), 2040 => to_unsigned(1974, 12), 2041 => to_unsigned(52, 12), 2042 => to_unsigned(215, 12), 2043 => to_unsigned(2395, 12), 2044 => to_unsigned(304, 12), 2045 => to_unsigned(831, 12), 2046 => to_unsigned(3348, 12), 2047 => to_unsigned(1555, 12)),
            6 => (0 => to_unsigned(2876, 12), 1 => to_unsigned(2932, 12), 2 => to_unsigned(3723, 12), 3 => to_unsigned(3290, 12), 4 => to_unsigned(1321, 12), 5 => to_unsigned(1065, 12), 6 => to_unsigned(3846, 12), 7 => to_unsigned(1633, 12), 8 => to_unsigned(2189, 12), 9 => to_unsigned(627, 12), 10 => to_unsigned(3202, 12), 11 => to_unsigned(813, 12), 12 => to_unsigned(2504, 12), 13 => to_unsigned(3613, 12), 14 => to_unsigned(3413, 12), 15 => to_unsigned(1264, 12), 16 => to_unsigned(479, 12), 17 => to_unsigned(3382, 12), 18 => to_unsigned(2615, 12), 19 => to_unsigned(3400, 12), 20 => to_unsigned(1458, 12), 21 => to_unsigned(2863, 12), 22 => to_unsigned(312, 12), 23 => to_unsigned(870, 12), 24 => to_unsigned(2939, 12), 25 => to_unsigned(1876, 12), 26 => to_unsigned(1304, 12), 27 => to_unsigned(2012, 12), 28 => to_unsigned(430, 12), 29 => to_unsigned(239, 12), 30 => to_unsigned(1642, 12), 31 => to_unsigned(1166, 12), 32 => to_unsigned(149, 12), 33 => to_unsigned(857, 12), 34 => to_unsigned(4052, 12), 35 => to_unsigned(1207, 12), 36 => to_unsigned(252, 12), 37 => to_unsigned(1248, 12), 38 => to_unsigned(1620, 12), 39 => to_unsigned(4072, 12), 40 => to_unsigned(2337, 12), 41 => to_unsigned(1164, 12), 42 => to_unsigned(2145, 12), 43 => to_unsigned(327, 12), 44 => to_unsigned(1673, 12), 45 => to_unsigned(2904, 12), 46 => to_unsigned(2702, 12), 47 => to_unsigned(2135, 12), 48 => to_unsigned(357, 12), 49 => to_unsigned(1925, 12), 50 => to_unsigned(1326, 12), 51 => to_unsigned(1257, 12), 52 => to_unsigned(750, 12), 53 => to_unsigned(1668, 12), 54 => to_unsigned(268, 12), 55 => to_unsigned(344, 12), 56 => to_unsigned(3153, 12), 57 => to_unsigned(1486, 12), 58 => to_unsigned(695, 12), 59 => to_unsigned(2126, 12), 60 => to_unsigned(849, 12), 61 => to_unsigned(2398, 12), 62 => to_unsigned(1033, 12), 63 => to_unsigned(677, 12), 64 => to_unsigned(1281, 12), 65 => to_unsigned(1971, 12), 66 => to_unsigned(2496, 12), 67 => to_unsigned(3823, 12), 68 => to_unsigned(4082, 12), 69 => to_unsigned(2586, 12), 70 => to_unsigned(3467, 12), 71 => to_unsigned(1831, 12), 72 => to_unsigned(3241, 12), 73 => to_unsigned(2516, 12), 74 => to_unsigned(2201, 12), 75 => to_unsigned(109, 12), 76 => to_unsigned(801, 12), 77 => to_unsigned(3570, 12), 78 => to_unsigned(2355, 12), 79 => to_unsigned(3830, 12), 80 => to_unsigned(1144, 12), 81 => to_unsigned(3349, 12), 82 => to_unsigned(2685, 12), 83 => to_unsigned(566, 12), 84 => to_unsigned(3663, 12), 85 => to_unsigned(353, 12), 86 => to_unsigned(3440, 12), 87 => to_unsigned(896, 12), 88 => to_unsigned(3851, 12), 89 => to_unsigned(2268, 12), 90 => to_unsigned(2849, 12), 91 => to_unsigned(4090, 12), 92 => to_unsigned(266, 12), 93 => to_unsigned(397, 12), 94 => to_unsigned(2005, 12), 95 => to_unsigned(3082, 12), 96 => to_unsigned(3303, 12), 97 => to_unsigned(2855, 12), 98 => to_unsigned(1824, 12), 99 => to_unsigned(3428, 12), 100 => to_unsigned(964, 12), 101 => to_unsigned(163, 12), 102 => to_unsigned(1736, 12), 103 => to_unsigned(2391, 12), 104 => to_unsigned(1111, 12), 105 => to_unsigned(3277, 12), 106 => to_unsigned(2660, 12), 107 => to_unsigned(2642, 12), 108 => to_unsigned(4031, 12), 109 => to_unsigned(174, 12), 110 => to_unsigned(738, 12), 111 => to_unsigned(338, 12), 112 => to_unsigned(1044, 12), 113 => to_unsigned(3098, 12), 114 => to_unsigned(2460, 12), 115 => to_unsigned(1804, 12), 116 => to_unsigned(2833, 12), 117 => to_unsigned(2434, 12), 118 => to_unsigned(4084, 12), 119 => to_unsigned(1828, 12), 120 => to_unsigned(3018, 12), 121 => to_unsigned(3618, 12), 122 => to_unsigned(935, 12), 123 => to_unsigned(1034, 12), 124 => to_unsigned(2611, 12), 125 => to_unsigned(130, 12), 126 => to_unsigned(193, 12), 127 => to_unsigned(1943, 12), 128 => to_unsigned(2432, 12), 129 => to_unsigned(380, 12), 130 => to_unsigned(1866, 12), 131 => to_unsigned(2555, 12), 132 => to_unsigned(3140, 12), 133 => to_unsigned(1428, 12), 134 => to_unsigned(3769, 12), 135 => to_unsigned(1285, 12), 136 => to_unsigned(3819, 12), 137 => to_unsigned(3940, 12), 138 => to_unsigned(2809, 12), 139 => to_unsigned(750, 12), 140 => to_unsigned(3587, 12), 141 => to_unsigned(365, 12), 142 => to_unsigned(3853, 12), 143 => to_unsigned(2654, 12), 144 => to_unsigned(1195, 12), 145 => to_unsigned(1282, 12), 146 => to_unsigned(2427, 12), 147 => to_unsigned(4001, 12), 148 => to_unsigned(3451, 12), 149 => to_unsigned(3483, 12), 150 => to_unsigned(1541, 12), 151 => to_unsigned(1587, 12), 152 => to_unsigned(1485, 12), 153 => to_unsigned(933, 12), 154 => to_unsigned(3863, 12), 155 => to_unsigned(143, 12), 156 => to_unsigned(1610, 12), 157 => to_unsigned(3804, 12), 158 => to_unsigned(2467, 12), 159 => to_unsigned(1944, 12), 160 => to_unsigned(606, 12), 161 => to_unsigned(1469, 12), 162 => to_unsigned(2357, 12), 163 => to_unsigned(2303, 12), 164 => to_unsigned(1900, 12), 165 => to_unsigned(87, 12), 166 => to_unsigned(3464, 12), 167 => to_unsigned(925, 12), 168 => to_unsigned(1374, 12), 169 => to_unsigned(1123, 12), 170 => to_unsigned(1482, 12), 171 => to_unsigned(878, 12), 172 => to_unsigned(921, 12), 173 => to_unsigned(2437, 12), 174 => to_unsigned(493, 12), 175 => to_unsigned(645, 12), 176 => to_unsigned(1124, 12), 177 => to_unsigned(670, 12), 178 => to_unsigned(1795, 12), 179 => to_unsigned(1400, 12), 180 => to_unsigned(2059, 12), 181 => to_unsigned(2233, 12), 182 => to_unsigned(3099, 12), 183 => to_unsigned(1000, 12), 184 => to_unsigned(3712, 12), 185 => to_unsigned(4059, 12), 186 => to_unsigned(3211, 12), 187 => to_unsigned(1188, 12), 188 => to_unsigned(66, 12), 189 => to_unsigned(2965, 12), 190 => to_unsigned(969, 12), 191 => to_unsigned(2654, 12), 192 => to_unsigned(1850, 12), 193 => to_unsigned(2302, 12), 194 => to_unsigned(1819, 12), 195 => to_unsigned(3986, 12), 196 => to_unsigned(1141, 12), 197 => to_unsigned(2670, 12), 198 => to_unsigned(433, 12), 199 => to_unsigned(890, 12), 200 => to_unsigned(825, 12), 201 => to_unsigned(984, 12), 202 => to_unsigned(2600, 12), 203 => to_unsigned(3123, 12), 204 => to_unsigned(3478, 12), 205 => to_unsigned(626, 12), 206 => to_unsigned(1821, 12), 207 => to_unsigned(2485, 12), 208 => to_unsigned(1704, 12), 209 => to_unsigned(3885, 12), 210 => to_unsigned(2098, 12), 211 => to_unsigned(4021, 12), 212 => to_unsigned(2640, 12), 213 => to_unsigned(231, 12), 214 => to_unsigned(523, 12), 215 => to_unsigned(2848, 12), 216 => to_unsigned(616, 12), 217 => to_unsigned(825, 12), 218 => to_unsigned(895, 12), 219 => to_unsigned(3739, 12), 220 => to_unsigned(3980, 12), 221 => to_unsigned(1358, 12), 222 => to_unsigned(2738, 12), 223 => to_unsigned(1980, 12), 224 => to_unsigned(2893, 12), 225 => to_unsigned(958, 12), 226 => to_unsigned(436, 12), 227 => to_unsigned(3521, 12), 228 => to_unsigned(2236, 12), 229 => to_unsigned(3231, 12), 230 => to_unsigned(3184, 12), 231 => to_unsigned(305, 12), 232 => to_unsigned(1737, 12), 233 => to_unsigned(509, 12), 234 => to_unsigned(2281, 12), 235 => to_unsigned(2958, 12), 236 => to_unsigned(2255, 12), 237 => to_unsigned(523, 12), 238 => to_unsigned(1732, 12), 239 => to_unsigned(801, 12), 240 => to_unsigned(2029, 12), 241 => to_unsigned(2232, 12), 242 => to_unsigned(760, 12), 243 => to_unsigned(425, 12), 244 => to_unsigned(667, 12), 245 => to_unsigned(434, 12), 246 => to_unsigned(2655, 12), 247 => to_unsigned(145, 12), 248 => to_unsigned(1423, 12), 249 => to_unsigned(422, 12), 250 => to_unsigned(1922, 12), 251 => to_unsigned(3925, 12), 252 => to_unsigned(1699, 12), 253 => to_unsigned(529, 12), 254 => to_unsigned(1447, 12), 255 => to_unsigned(734, 12), 256 => to_unsigned(2751, 12), 257 => to_unsigned(2553, 12), 258 => to_unsigned(120, 12), 259 => to_unsigned(305, 12), 260 => to_unsigned(1161, 12), 261 => to_unsigned(2073, 12), 262 => to_unsigned(1693, 12), 263 => to_unsigned(3312, 12), 264 => to_unsigned(2498, 12), 265 => to_unsigned(3696, 12), 266 => to_unsigned(1536, 12), 267 => to_unsigned(433, 12), 268 => to_unsigned(3289, 12), 269 => to_unsigned(3311, 12), 270 => to_unsigned(1797, 12), 271 => to_unsigned(2900, 12), 272 => to_unsigned(653, 12), 273 => to_unsigned(2853, 12), 274 => to_unsigned(2132, 12), 275 => to_unsigned(3691, 12), 276 => to_unsigned(1822, 12), 277 => to_unsigned(444, 12), 278 => to_unsigned(313, 12), 279 => to_unsigned(2555, 12), 280 => to_unsigned(1666, 12), 281 => to_unsigned(3493, 12), 282 => to_unsigned(2484, 12), 283 => to_unsigned(1430, 12), 284 => to_unsigned(3165, 12), 285 => to_unsigned(3924, 12), 286 => to_unsigned(65, 12), 287 => to_unsigned(1065, 12), 288 => to_unsigned(376, 12), 289 => to_unsigned(2134, 12), 290 => to_unsigned(2998, 12), 291 => to_unsigned(1479, 12), 292 => to_unsigned(38, 12), 293 => to_unsigned(400, 12), 294 => to_unsigned(1972, 12), 295 => to_unsigned(2652, 12), 296 => to_unsigned(179, 12), 297 => to_unsigned(237, 12), 298 => to_unsigned(2135, 12), 299 => to_unsigned(540, 12), 300 => to_unsigned(3246, 12), 301 => to_unsigned(2185, 12), 302 => to_unsigned(3497, 12), 303 => to_unsigned(3739, 12), 304 => to_unsigned(3983, 12), 305 => to_unsigned(282, 12), 306 => to_unsigned(4047, 12), 307 => to_unsigned(3058, 12), 308 => to_unsigned(494, 12), 309 => to_unsigned(3065, 12), 310 => to_unsigned(3726, 12), 311 => to_unsigned(2022, 12), 312 => to_unsigned(1680, 12), 313 => to_unsigned(669, 12), 314 => to_unsigned(2493, 12), 315 => to_unsigned(978, 12), 316 => to_unsigned(3590, 12), 317 => to_unsigned(3576, 12), 318 => to_unsigned(3127, 12), 319 => to_unsigned(2625, 12), 320 => to_unsigned(2129, 12), 321 => to_unsigned(3712, 12), 322 => to_unsigned(1438, 12), 323 => to_unsigned(49, 12), 324 => to_unsigned(2036, 12), 325 => to_unsigned(318, 12), 326 => to_unsigned(3073, 12), 327 => to_unsigned(508, 12), 328 => to_unsigned(1995, 12), 329 => to_unsigned(3743, 12), 330 => to_unsigned(3616, 12), 331 => to_unsigned(1354, 12), 332 => to_unsigned(2435, 12), 333 => to_unsigned(1853, 12), 334 => to_unsigned(1880, 12), 335 => to_unsigned(2170, 12), 336 => to_unsigned(2444, 12), 337 => to_unsigned(2586, 12), 338 => to_unsigned(1796, 12), 339 => to_unsigned(3753, 12), 340 => to_unsigned(177, 12), 341 => to_unsigned(4046, 12), 342 => to_unsigned(3988, 12), 343 => to_unsigned(699, 12), 344 => to_unsigned(1066, 12), 345 => to_unsigned(3726, 12), 346 => to_unsigned(310, 12), 347 => to_unsigned(2436, 12), 348 => to_unsigned(59, 12), 349 => to_unsigned(1330, 12), 350 => to_unsigned(2775, 12), 351 => to_unsigned(251, 12), 352 => to_unsigned(2420, 12), 353 => to_unsigned(3594, 12), 354 => to_unsigned(2418, 12), 355 => to_unsigned(267, 12), 356 => to_unsigned(341, 12), 357 => to_unsigned(2489, 12), 358 => to_unsigned(962, 12), 359 => to_unsigned(1661, 12), 360 => to_unsigned(3646, 12), 361 => to_unsigned(3723, 12), 362 => to_unsigned(3967, 12), 363 => to_unsigned(1353, 12), 364 => to_unsigned(2230, 12), 365 => to_unsigned(3509, 12), 366 => to_unsigned(1208, 12), 367 => to_unsigned(414, 12), 368 => to_unsigned(3563, 12), 369 => to_unsigned(1210, 12), 370 => to_unsigned(2984, 12), 371 => to_unsigned(2487, 12), 372 => to_unsigned(1644, 12), 373 => to_unsigned(1247, 12), 374 => to_unsigned(1880, 12), 375 => to_unsigned(1800, 12), 376 => to_unsigned(2000, 12), 377 => to_unsigned(209, 12), 378 => to_unsigned(989, 12), 379 => to_unsigned(3293, 12), 380 => to_unsigned(2319, 12), 381 => to_unsigned(1465, 12), 382 => to_unsigned(889, 12), 383 => to_unsigned(2695, 12), 384 => to_unsigned(1048, 12), 385 => to_unsigned(2250, 12), 386 => to_unsigned(1333, 12), 387 => to_unsigned(1202, 12), 388 => to_unsigned(3656, 12), 389 => to_unsigned(1790, 12), 390 => to_unsigned(1448, 12), 391 => to_unsigned(586, 12), 392 => to_unsigned(679, 12), 393 => to_unsigned(1763, 12), 394 => to_unsigned(2966, 12), 395 => to_unsigned(1535, 12), 396 => to_unsigned(1324, 12), 397 => to_unsigned(1968, 12), 398 => to_unsigned(3765, 12), 399 => to_unsigned(1920, 12), 400 => to_unsigned(1257, 12), 401 => to_unsigned(4049, 12), 402 => to_unsigned(456, 12), 403 => to_unsigned(3187, 12), 404 => to_unsigned(3606, 12), 405 => to_unsigned(2635, 12), 406 => to_unsigned(3293, 12), 407 => to_unsigned(509, 12), 408 => to_unsigned(3177, 12), 409 => to_unsigned(3764, 12), 410 => to_unsigned(160, 12), 411 => to_unsigned(814, 12), 412 => to_unsigned(1427, 12), 413 => to_unsigned(243, 12), 414 => to_unsigned(373, 12), 415 => to_unsigned(3622, 12), 416 => to_unsigned(96, 12), 417 => to_unsigned(1253, 12), 418 => to_unsigned(1071, 12), 419 => to_unsigned(2548, 12), 420 => to_unsigned(1327, 12), 421 => to_unsigned(1737, 12), 422 => to_unsigned(1200, 12), 423 => to_unsigned(3484, 12), 424 => to_unsigned(3282, 12), 425 => to_unsigned(2410, 12), 426 => to_unsigned(3316, 12), 427 => to_unsigned(661, 12), 428 => to_unsigned(542, 12), 429 => to_unsigned(2657, 12), 430 => to_unsigned(672, 12), 431 => to_unsigned(1735, 12), 432 => to_unsigned(2790, 12), 433 => to_unsigned(2147, 12), 434 => to_unsigned(408, 12), 435 => to_unsigned(1601, 12), 436 => to_unsigned(3794, 12), 437 => to_unsigned(822, 12), 438 => to_unsigned(701, 12), 439 => to_unsigned(3200, 12), 440 => to_unsigned(53, 12), 441 => to_unsigned(2644, 12), 442 => to_unsigned(2496, 12), 443 => to_unsigned(3125, 12), 444 => to_unsigned(2184, 12), 445 => to_unsigned(2638, 12), 446 => to_unsigned(3366, 12), 447 => to_unsigned(2002, 12), 448 => to_unsigned(3330, 12), 449 => to_unsigned(771, 12), 450 => to_unsigned(1462, 12), 451 => to_unsigned(658, 12), 452 => to_unsigned(814, 12), 453 => to_unsigned(1778, 12), 454 => to_unsigned(263, 12), 455 => to_unsigned(3832, 12), 456 => to_unsigned(3578, 12), 457 => to_unsigned(3334, 12), 458 => to_unsigned(2560, 12), 459 => to_unsigned(3528, 12), 460 => to_unsigned(1052, 12), 461 => to_unsigned(3088, 12), 462 => to_unsigned(3115, 12), 463 => to_unsigned(2271, 12), 464 => to_unsigned(1848, 12), 465 => to_unsigned(1648, 12), 466 => to_unsigned(489, 12), 467 => to_unsigned(2907, 12), 468 => to_unsigned(329, 12), 469 => to_unsigned(1572, 12), 470 => to_unsigned(359, 12), 471 => to_unsigned(3751, 12), 472 => to_unsigned(2823, 12), 473 => to_unsigned(672, 12), 474 => to_unsigned(782, 12), 475 => to_unsigned(1422, 12), 476 => to_unsigned(383, 12), 477 => to_unsigned(1891, 12), 478 => to_unsigned(2655, 12), 479 => to_unsigned(2939, 12), 480 => to_unsigned(1548, 12), 481 => to_unsigned(2546, 12), 482 => to_unsigned(635, 12), 483 => to_unsigned(2570, 12), 484 => to_unsigned(1444, 12), 485 => to_unsigned(4046, 12), 486 => to_unsigned(3589, 12), 487 => to_unsigned(2191, 12), 488 => to_unsigned(2165, 12), 489 => to_unsigned(626, 12), 490 => to_unsigned(3917, 12), 491 => to_unsigned(2132, 12), 492 => to_unsigned(1768, 12), 493 => to_unsigned(1424, 12), 494 => to_unsigned(80, 12), 495 => to_unsigned(1713, 12), 496 => to_unsigned(3547, 12), 497 => to_unsigned(1900, 12), 498 => to_unsigned(1050, 12), 499 => to_unsigned(1684, 12), 500 => to_unsigned(425, 12), 501 => to_unsigned(2986, 12), 502 => to_unsigned(2734, 12), 503 => to_unsigned(1566, 12), 504 => to_unsigned(929, 12), 505 => to_unsigned(1791, 12), 506 => to_unsigned(3258, 12), 507 => to_unsigned(1971, 12), 508 => to_unsigned(4040, 12), 509 => to_unsigned(3464, 12), 510 => to_unsigned(2075, 12), 511 => to_unsigned(1629, 12), 512 => to_unsigned(323, 12), 513 => to_unsigned(549, 12), 514 => to_unsigned(2872, 12), 515 => to_unsigned(1356, 12), 516 => to_unsigned(2, 12), 517 => to_unsigned(1996, 12), 518 => to_unsigned(3868, 12), 519 => to_unsigned(1907, 12), 520 => to_unsigned(207, 12), 521 => to_unsigned(3208, 12), 522 => to_unsigned(158, 12), 523 => to_unsigned(1626, 12), 524 => to_unsigned(1277, 12), 525 => to_unsigned(2078, 12), 526 => to_unsigned(3376, 12), 527 => to_unsigned(2149, 12), 528 => to_unsigned(40, 12), 529 => to_unsigned(2048, 12), 530 => to_unsigned(875, 12), 531 => to_unsigned(912, 12), 532 => to_unsigned(1808, 12), 533 => to_unsigned(341, 12), 534 => to_unsigned(3525, 12), 535 => to_unsigned(2666, 12), 536 => to_unsigned(142, 12), 537 => to_unsigned(3275, 12), 538 => to_unsigned(3692, 12), 539 => to_unsigned(3705, 12), 540 => to_unsigned(2055, 12), 541 => to_unsigned(3613, 12), 542 => to_unsigned(1191, 12), 543 => to_unsigned(200, 12), 544 => to_unsigned(944, 12), 545 => to_unsigned(1191, 12), 546 => to_unsigned(1423, 12), 547 => to_unsigned(2146, 12), 548 => to_unsigned(564, 12), 549 => to_unsigned(1489, 12), 550 => to_unsigned(3530, 12), 551 => to_unsigned(2374, 12), 552 => to_unsigned(615, 12), 553 => to_unsigned(2729, 12), 554 => to_unsigned(650, 12), 555 => to_unsigned(847, 12), 556 => to_unsigned(2639, 12), 557 => to_unsigned(370, 12), 558 => to_unsigned(2285, 12), 559 => to_unsigned(2038, 12), 560 => to_unsigned(1171, 12), 561 => to_unsigned(3626, 12), 562 => to_unsigned(2989, 12), 563 => to_unsigned(860, 12), 564 => to_unsigned(323, 12), 565 => to_unsigned(3433, 12), 566 => to_unsigned(2862, 12), 567 => to_unsigned(3286, 12), 568 => to_unsigned(1453, 12), 569 => to_unsigned(3611, 12), 570 => to_unsigned(1453, 12), 571 => to_unsigned(585, 12), 572 => to_unsigned(281, 12), 573 => to_unsigned(145, 12), 574 => to_unsigned(3898, 12), 575 => to_unsigned(293, 12), 576 => to_unsigned(68, 12), 577 => to_unsigned(3347, 12), 578 => to_unsigned(1721, 12), 579 => to_unsigned(132, 12), 580 => to_unsigned(1598, 12), 581 => to_unsigned(1393, 12), 582 => to_unsigned(617, 12), 583 => to_unsigned(2192, 12), 584 => to_unsigned(2897, 12), 585 => to_unsigned(384, 12), 586 => to_unsigned(2480, 12), 587 => to_unsigned(287, 12), 588 => to_unsigned(2037, 12), 589 => to_unsigned(1833, 12), 590 => to_unsigned(3999, 12), 591 => to_unsigned(1860, 12), 592 => to_unsigned(1637, 12), 593 => to_unsigned(2972, 12), 594 => to_unsigned(2194, 12), 595 => to_unsigned(2911, 12), 596 => to_unsigned(2687, 12), 597 => to_unsigned(912, 12), 598 => to_unsigned(3910, 12), 599 => to_unsigned(3188, 12), 600 => to_unsigned(3950, 12), 601 => to_unsigned(1748, 12), 602 => to_unsigned(2594, 12), 603 => to_unsigned(3240, 12), 604 => to_unsigned(3790, 12), 605 => to_unsigned(1625, 12), 606 => to_unsigned(614, 12), 607 => to_unsigned(3511, 12), 608 => to_unsigned(2583, 12), 609 => to_unsigned(3926, 12), 610 => to_unsigned(342, 12), 611 => to_unsigned(2623, 12), 612 => to_unsigned(2223, 12), 613 => to_unsigned(2592, 12), 614 => to_unsigned(1655, 12), 615 => to_unsigned(1325, 12), 616 => to_unsigned(85, 12), 617 => to_unsigned(379, 12), 618 => to_unsigned(492, 12), 619 => to_unsigned(394, 12), 620 => to_unsigned(728, 12), 621 => to_unsigned(2890, 12), 622 => to_unsigned(2987, 12), 623 => to_unsigned(2537, 12), 624 => to_unsigned(1215, 12), 625 => to_unsigned(441, 12), 626 => to_unsigned(2668, 12), 627 => to_unsigned(2888, 12), 628 => to_unsigned(923, 12), 629 => to_unsigned(3376, 12), 630 => to_unsigned(3896, 12), 631 => to_unsigned(2855, 12), 632 => to_unsigned(1514, 12), 633 => to_unsigned(1692, 12), 634 => to_unsigned(3726, 12), 635 => to_unsigned(116, 12), 636 => to_unsigned(2078, 12), 637 => to_unsigned(1439, 12), 638 => to_unsigned(3454, 12), 639 => to_unsigned(64, 12), 640 => to_unsigned(3904, 12), 641 => to_unsigned(2187, 12), 642 => to_unsigned(1015, 12), 643 => to_unsigned(2341, 12), 644 => to_unsigned(1664, 12), 645 => to_unsigned(3703, 12), 646 => to_unsigned(2924, 12), 647 => to_unsigned(290, 12), 648 => to_unsigned(3963, 12), 649 => to_unsigned(1042, 12), 650 => to_unsigned(2848, 12), 651 => to_unsigned(422, 12), 652 => to_unsigned(1951, 12), 653 => to_unsigned(1419, 12), 654 => to_unsigned(2941, 12), 655 => to_unsigned(3190, 12), 656 => to_unsigned(3287, 12), 657 => to_unsigned(1234, 12), 658 => to_unsigned(1947, 12), 659 => to_unsigned(2849, 12), 660 => to_unsigned(3849, 12), 661 => to_unsigned(1925, 12), 662 => to_unsigned(2756, 12), 663 => to_unsigned(3582, 12), 664 => to_unsigned(1667, 12), 665 => to_unsigned(1133, 12), 666 => to_unsigned(1483, 12), 667 => to_unsigned(1548, 12), 668 => to_unsigned(1865, 12), 669 => to_unsigned(3211, 12), 670 => to_unsigned(3981, 12), 671 => to_unsigned(3063, 12), 672 => to_unsigned(255, 12), 673 => to_unsigned(933, 12), 674 => to_unsigned(741, 12), 675 => to_unsigned(628, 12), 676 => to_unsigned(3220, 12), 677 => to_unsigned(307, 12), 678 => to_unsigned(1225, 12), 679 => to_unsigned(1957, 12), 680 => to_unsigned(2533, 12), 681 => to_unsigned(762, 12), 682 => to_unsigned(3609, 12), 683 => to_unsigned(557, 12), 684 => to_unsigned(771, 12), 685 => to_unsigned(531, 12), 686 => to_unsigned(2958, 12), 687 => to_unsigned(1203, 12), 688 => to_unsigned(1398, 12), 689 => to_unsigned(3929, 12), 690 => to_unsigned(3458, 12), 691 => to_unsigned(74, 12), 692 => to_unsigned(1590, 12), 693 => to_unsigned(2439, 12), 694 => to_unsigned(708, 12), 695 => to_unsigned(2182, 12), 696 => to_unsigned(3140, 12), 697 => to_unsigned(2600, 12), 698 => to_unsigned(2144, 12), 699 => to_unsigned(1176, 12), 700 => to_unsigned(1935, 12), 701 => to_unsigned(4088, 12), 702 => to_unsigned(1074, 12), 703 => to_unsigned(3990, 12), 704 => to_unsigned(2915, 12), 705 => to_unsigned(2383, 12), 706 => to_unsigned(4054, 12), 707 => to_unsigned(1518, 12), 708 => to_unsigned(714, 12), 709 => to_unsigned(3250, 12), 710 => to_unsigned(2212, 12), 711 => to_unsigned(2194, 12), 712 => to_unsigned(622, 12), 713 => to_unsigned(1717, 12), 714 => to_unsigned(384, 12), 715 => to_unsigned(325, 12), 716 => to_unsigned(2941, 12), 717 => to_unsigned(1604, 12), 718 => to_unsigned(2216, 12), 719 => to_unsigned(1196, 12), 720 => to_unsigned(1036, 12), 721 => to_unsigned(2053, 12), 722 => to_unsigned(3593, 12), 723 => to_unsigned(3868, 12), 724 => to_unsigned(3841, 12), 725 => to_unsigned(3195, 12), 726 => to_unsigned(2526, 12), 727 => to_unsigned(3351, 12), 728 => to_unsigned(1232, 12), 729 => to_unsigned(3599, 12), 730 => to_unsigned(2086, 12), 731 => to_unsigned(450, 12), 732 => to_unsigned(1375, 12), 733 => to_unsigned(3035, 12), 734 => to_unsigned(1634, 12), 735 => to_unsigned(1718, 12), 736 => to_unsigned(1086, 12), 737 => to_unsigned(1248, 12), 738 => to_unsigned(402, 12), 739 => to_unsigned(1868, 12), 740 => to_unsigned(3483, 12), 741 => to_unsigned(3631, 12), 742 => to_unsigned(469, 12), 743 => to_unsigned(601, 12), 744 => to_unsigned(4010, 12), 745 => to_unsigned(1243, 12), 746 => to_unsigned(3121, 12), 747 => to_unsigned(1151, 12), 748 => to_unsigned(2216, 12), 749 => to_unsigned(4080, 12), 750 => to_unsigned(827, 12), 751 => to_unsigned(1542, 12), 752 => to_unsigned(1321, 12), 753 => to_unsigned(774, 12), 754 => to_unsigned(2277, 12), 755 => to_unsigned(1155, 12), 756 => to_unsigned(3795, 12), 757 => to_unsigned(1878, 12), 758 => to_unsigned(3201, 12), 759 => to_unsigned(2868, 12), 760 => to_unsigned(3670, 12), 761 => to_unsigned(3810, 12), 762 => to_unsigned(3133, 12), 763 => to_unsigned(2230, 12), 764 => to_unsigned(445, 12), 765 => to_unsigned(2722, 12), 766 => to_unsigned(978, 12), 767 => to_unsigned(707, 12), 768 => to_unsigned(2306, 12), 769 => to_unsigned(2283, 12), 770 => to_unsigned(619, 12), 771 => to_unsigned(417, 12), 772 => to_unsigned(1408, 12), 773 => to_unsigned(1655, 12), 774 => to_unsigned(2001, 12), 775 => to_unsigned(3812, 12), 776 => to_unsigned(791, 12), 777 => to_unsigned(762, 12), 778 => to_unsigned(1857, 12), 779 => to_unsigned(321, 12), 780 => to_unsigned(257, 12), 781 => to_unsigned(503, 12), 782 => to_unsigned(2580, 12), 783 => to_unsigned(2124, 12), 784 => to_unsigned(1226, 12), 785 => to_unsigned(1887, 12), 786 => to_unsigned(1062, 12), 787 => to_unsigned(1477, 12), 788 => to_unsigned(2232, 12), 789 => to_unsigned(789, 12), 790 => to_unsigned(2906, 12), 791 => to_unsigned(1213, 12), 792 => to_unsigned(1381, 12), 793 => to_unsigned(840, 12), 794 => to_unsigned(1416, 12), 795 => to_unsigned(636, 12), 796 => to_unsigned(1948, 12), 797 => to_unsigned(1279, 12), 798 => to_unsigned(1125, 12), 799 => to_unsigned(3982, 12), 800 => to_unsigned(3839, 12), 801 => to_unsigned(1617, 12), 802 => to_unsigned(2482, 12), 803 => to_unsigned(32, 12), 804 => to_unsigned(2296, 12), 805 => to_unsigned(1591, 12), 806 => to_unsigned(1752, 12), 807 => to_unsigned(1798, 12), 808 => to_unsigned(4085, 12), 809 => to_unsigned(3327, 12), 810 => to_unsigned(15, 12), 811 => to_unsigned(3305, 12), 812 => to_unsigned(1380, 12), 813 => to_unsigned(2831, 12), 814 => to_unsigned(3676, 12), 815 => to_unsigned(3801, 12), 816 => to_unsigned(3470, 12), 817 => to_unsigned(3862, 12), 818 => to_unsigned(3778, 12), 819 => to_unsigned(2010, 12), 820 => to_unsigned(1553, 12), 821 => to_unsigned(3564, 12), 822 => to_unsigned(2095, 12), 823 => to_unsigned(2706, 12), 824 => to_unsigned(88, 12), 825 => to_unsigned(2824, 12), 826 => to_unsigned(1908, 12), 827 => to_unsigned(2710, 12), 828 => to_unsigned(3289, 12), 829 => to_unsigned(3401, 12), 830 => to_unsigned(3855, 12), 831 => to_unsigned(1759, 12), 832 => to_unsigned(2802, 12), 833 => to_unsigned(1004, 12), 834 => to_unsigned(3516, 12), 835 => to_unsigned(2861, 12), 836 => to_unsigned(1562, 12), 837 => to_unsigned(911, 12), 838 => to_unsigned(2244, 12), 839 => to_unsigned(383, 12), 840 => to_unsigned(236, 12), 841 => to_unsigned(1149, 12), 842 => to_unsigned(3722, 12), 843 => to_unsigned(1876, 12), 844 => to_unsigned(3247, 12), 845 => to_unsigned(942, 12), 846 => to_unsigned(2933, 12), 847 => to_unsigned(2351, 12), 848 => to_unsigned(3653, 12), 849 => to_unsigned(2606, 12), 850 => to_unsigned(794, 12), 851 => to_unsigned(3677, 12), 852 => to_unsigned(2549, 12), 853 => to_unsigned(3501, 12), 854 => to_unsigned(2567, 12), 855 => to_unsigned(771, 12), 856 => to_unsigned(1945, 12), 857 => to_unsigned(2753, 12), 858 => to_unsigned(3356, 12), 859 => to_unsigned(847, 12), 860 => to_unsigned(3952, 12), 861 => to_unsigned(3655, 12), 862 => to_unsigned(3120, 12), 863 => to_unsigned(1279, 12), 864 => to_unsigned(3942, 12), 865 => to_unsigned(2759, 12), 866 => to_unsigned(2401, 12), 867 => to_unsigned(1798, 12), 868 => to_unsigned(2552, 12), 869 => to_unsigned(1362, 12), 870 => to_unsigned(546, 12), 871 => to_unsigned(3237, 12), 872 => to_unsigned(1893, 12), 873 => to_unsigned(1635, 12), 874 => to_unsigned(744, 12), 875 => to_unsigned(785, 12), 876 => to_unsigned(107, 12), 877 => to_unsigned(447, 12), 878 => to_unsigned(1430, 12), 879 => to_unsigned(1956, 12), 880 => to_unsigned(1042, 12), 881 => to_unsigned(585, 12), 882 => to_unsigned(3205, 12), 883 => to_unsigned(2183, 12), 884 => to_unsigned(3606, 12), 885 => to_unsigned(2321, 12), 886 => to_unsigned(3240, 12), 887 => to_unsigned(81, 12), 888 => to_unsigned(3164, 12), 889 => to_unsigned(3902, 12), 890 => to_unsigned(216, 12), 891 => to_unsigned(2720, 12), 892 => to_unsigned(891, 12), 893 => to_unsigned(688, 12), 894 => to_unsigned(1763, 12), 895 => to_unsigned(3996, 12), 896 => to_unsigned(1433, 12), 897 => to_unsigned(1693, 12), 898 => to_unsigned(156, 12), 899 => to_unsigned(1239, 12), 900 => to_unsigned(1528, 12), 901 => to_unsigned(958, 12), 902 => to_unsigned(2633, 12), 903 => to_unsigned(1901, 12), 904 => to_unsigned(1609, 12), 905 => to_unsigned(3274, 12), 906 => to_unsigned(1301, 12), 907 => to_unsigned(1942, 12), 908 => to_unsigned(2684, 12), 909 => to_unsigned(1499, 12), 910 => to_unsigned(2564, 12), 911 => to_unsigned(1846, 12), 912 => to_unsigned(2279, 12), 913 => to_unsigned(780, 12), 914 => to_unsigned(3265, 12), 915 => to_unsigned(3724, 12), 916 => to_unsigned(3220, 12), 917 => to_unsigned(1165, 12), 918 => to_unsigned(756, 12), 919 => to_unsigned(1050, 12), 920 => to_unsigned(705, 12), 921 => to_unsigned(883, 12), 922 => to_unsigned(2032, 12), 923 => to_unsigned(2401, 12), 924 => to_unsigned(2565, 12), 925 => to_unsigned(2734, 12), 926 => to_unsigned(1994, 12), 927 => to_unsigned(3363, 12), 928 => to_unsigned(104, 12), 929 => to_unsigned(409, 12), 930 => to_unsigned(3119, 12), 931 => to_unsigned(1536, 12), 932 => to_unsigned(149, 12), 933 => to_unsigned(2695, 12), 934 => to_unsigned(2818, 12), 935 => to_unsigned(1668, 12), 936 => to_unsigned(1720, 12), 937 => to_unsigned(369, 12), 938 => to_unsigned(890, 12), 939 => to_unsigned(3106, 12), 940 => to_unsigned(510, 12), 941 => to_unsigned(54, 12), 942 => to_unsigned(1046, 12), 943 => to_unsigned(1231, 12), 944 => to_unsigned(2453, 12), 945 => to_unsigned(2029, 12), 946 => to_unsigned(3458, 12), 947 => to_unsigned(2895, 12), 948 => to_unsigned(820, 12), 949 => to_unsigned(3351, 12), 950 => to_unsigned(1374, 12), 951 => to_unsigned(1197, 12), 952 => to_unsigned(2812, 12), 953 => to_unsigned(3901, 12), 954 => to_unsigned(246, 12), 955 => to_unsigned(1777, 12), 956 => to_unsigned(786, 12), 957 => to_unsigned(283, 12), 958 => to_unsigned(3282, 12), 959 => to_unsigned(2697, 12), 960 => to_unsigned(3525, 12), 961 => to_unsigned(2530, 12), 962 => to_unsigned(2170, 12), 963 => to_unsigned(23, 12), 964 => to_unsigned(3911, 12), 965 => to_unsigned(2462, 12), 966 => to_unsigned(2407, 12), 967 => to_unsigned(363, 12), 968 => to_unsigned(3209, 12), 969 => to_unsigned(1490, 12), 970 => to_unsigned(276, 12), 971 => to_unsigned(3664, 12), 972 => to_unsigned(1267, 12), 973 => to_unsigned(3181, 12), 974 => to_unsigned(2667, 12), 975 => to_unsigned(2006, 12), 976 => to_unsigned(3985, 12), 977 => to_unsigned(3548, 12), 978 => to_unsigned(476, 12), 979 => to_unsigned(2860, 12), 980 => to_unsigned(401, 12), 981 => to_unsigned(1577, 12), 982 => to_unsigned(2825, 12), 983 => to_unsigned(2071, 12), 984 => to_unsigned(3277, 12), 985 => to_unsigned(455, 12), 986 => to_unsigned(2047, 12), 987 => to_unsigned(3546, 12), 988 => to_unsigned(3482, 12), 989 => to_unsigned(3219, 12), 990 => to_unsigned(3395, 12), 991 => to_unsigned(2744, 12), 992 => to_unsigned(2312, 12), 993 => to_unsigned(3118, 12), 994 => to_unsigned(1275, 12), 995 => to_unsigned(1480, 12), 996 => to_unsigned(642, 12), 997 => to_unsigned(2939, 12), 998 => to_unsigned(3589, 12), 999 => to_unsigned(2446, 12), 1000 => to_unsigned(1185, 12), 1001 => to_unsigned(1092, 12), 1002 => to_unsigned(1270, 12), 1003 => to_unsigned(737, 12), 1004 => to_unsigned(360, 12), 1005 => to_unsigned(2113, 12), 1006 => to_unsigned(819, 12), 1007 => to_unsigned(1835, 12), 1008 => to_unsigned(3320, 12), 1009 => to_unsigned(2926, 12), 1010 => to_unsigned(1411, 12), 1011 => to_unsigned(3433, 12), 1012 => to_unsigned(3124, 12), 1013 => to_unsigned(472, 12), 1014 => to_unsigned(4, 12), 1015 => to_unsigned(538, 12), 1016 => to_unsigned(2462, 12), 1017 => to_unsigned(164, 12), 1018 => to_unsigned(3758, 12), 1019 => to_unsigned(891, 12), 1020 => to_unsigned(969, 12), 1021 => to_unsigned(3591, 12), 1022 => to_unsigned(2460, 12), 1023 => to_unsigned(2156, 12), 1024 => to_unsigned(270, 12), 1025 => to_unsigned(2745, 12), 1026 => to_unsigned(1150, 12), 1027 => to_unsigned(415, 12), 1028 => to_unsigned(1832, 12), 1029 => to_unsigned(2753, 12), 1030 => to_unsigned(3797, 12), 1031 => to_unsigned(405, 12), 1032 => to_unsigned(3174, 12), 1033 => to_unsigned(2527, 12), 1034 => to_unsigned(3794, 12), 1035 => to_unsigned(1020, 12), 1036 => to_unsigned(3103, 12), 1037 => to_unsigned(1761, 12), 1038 => to_unsigned(2950, 12), 1039 => to_unsigned(2972, 12), 1040 => to_unsigned(728, 12), 1041 => to_unsigned(980, 12), 1042 => to_unsigned(3356, 12), 1043 => to_unsigned(17, 12), 1044 => to_unsigned(3111, 12), 1045 => to_unsigned(1168, 12), 1046 => to_unsigned(2106, 12), 1047 => to_unsigned(1025, 12), 1048 => to_unsigned(2921, 12), 1049 => to_unsigned(2357, 12), 1050 => to_unsigned(2885, 12), 1051 => to_unsigned(311, 12), 1052 => to_unsigned(3896, 12), 1053 => to_unsigned(3171, 12), 1054 => to_unsigned(3492, 12), 1055 => to_unsigned(3577, 12), 1056 => to_unsigned(2719, 12), 1057 => to_unsigned(616, 12), 1058 => to_unsigned(3965, 12), 1059 => to_unsigned(577, 12), 1060 => to_unsigned(1384, 12), 1061 => to_unsigned(735, 12), 1062 => to_unsigned(224, 12), 1063 => to_unsigned(2706, 12), 1064 => to_unsigned(3304, 12), 1065 => to_unsigned(1822, 12), 1066 => to_unsigned(1806, 12), 1067 => to_unsigned(725, 12), 1068 => to_unsigned(2271, 12), 1069 => to_unsigned(1440, 12), 1070 => to_unsigned(139, 12), 1071 => to_unsigned(2918, 12), 1072 => to_unsigned(236, 12), 1073 => to_unsigned(1102, 12), 1074 => to_unsigned(783, 12), 1075 => to_unsigned(2695, 12), 1076 => to_unsigned(3015, 12), 1077 => to_unsigned(330, 12), 1078 => to_unsigned(3518, 12), 1079 => to_unsigned(1876, 12), 1080 => to_unsigned(3233, 12), 1081 => to_unsigned(1527, 12), 1082 => to_unsigned(3090, 12), 1083 => to_unsigned(3583, 12), 1084 => to_unsigned(170, 12), 1085 => to_unsigned(4072, 12), 1086 => to_unsigned(155, 12), 1087 => to_unsigned(792, 12), 1088 => to_unsigned(69, 12), 1089 => to_unsigned(3267, 12), 1090 => to_unsigned(3997, 12), 1091 => to_unsigned(2718, 12), 1092 => to_unsigned(1119, 12), 1093 => to_unsigned(802, 12), 1094 => to_unsigned(1050, 12), 1095 => to_unsigned(963, 12), 1096 => to_unsigned(2544, 12), 1097 => to_unsigned(23, 12), 1098 => to_unsigned(1224, 12), 1099 => to_unsigned(490, 12), 1100 => to_unsigned(1944, 12), 1101 => to_unsigned(1002, 12), 1102 => to_unsigned(2438, 12), 1103 => to_unsigned(842, 12), 1104 => to_unsigned(2941, 12), 1105 => to_unsigned(1913, 12), 1106 => to_unsigned(3055, 12), 1107 => to_unsigned(3683, 12), 1108 => to_unsigned(1451, 12), 1109 => to_unsigned(1646, 12), 1110 => to_unsigned(3321, 12), 1111 => to_unsigned(1255, 12), 1112 => to_unsigned(751, 12), 1113 => to_unsigned(241, 12), 1114 => to_unsigned(1588, 12), 1115 => to_unsigned(1754, 12), 1116 => to_unsigned(3117, 12), 1117 => to_unsigned(2532, 12), 1118 => to_unsigned(2511, 12), 1119 => to_unsigned(2962, 12), 1120 => to_unsigned(2819, 12), 1121 => to_unsigned(4060, 12), 1122 => to_unsigned(3391, 12), 1123 => to_unsigned(186, 12), 1124 => to_unsigned(3519, 12), 1125 => to_unsigned(2471, 12), 1126 => to_unsigned(478, 12), 1127 => to_unsigned(1413, 12), 1128 => to_unsigned(1455, 12), 1129 => to_unsigned(3734, 12), 1130 => to_unsigned(3691, 12), 1131 => to_unsigned(51, 12), 1132 => to_unsigned(2609, 12), 1133 => to_unsigned(1609, 12), 1134 => to_unsigned(908, 12), 1135 => to_unsigned(2464, 12), 1136 => to_unsigned(2383, 12), 1137 => to_unsigned(1014, 12), 1138 => to_unsigned(1824, 12), 1139 => to_unsigned(1827, 12), 1140 => to_unsigned(2546, 12), 1141 => to_unsigned(764, 12), 1142 => to_unsigned(2558, 12), 1143 => to_unsigned(1596, 12), 1144 => to_unsigned(3902, 12), 1145 => to_unsigned(1519, 12), 1146 => to_unsigned(1372, 12), 1147 => to_unsigned(2431, 12), 1148 => to_unsigned(3546, 12), 1149 => to_unsigned(739, 12), 1150 => to_unsigned(3666, 12), 1151 => to_unsigned(1452, 12), 1152 => to_unsigned(3306, 12), 1153 => to_unsigned(3507, 12), 1154 => to_unsigned(2616, 12), 1155 => to_unsigned(3548, 12), 1156 => to_unsigned(2312, 12), 1157 => to_unsigned(945, 12), 1158 => to_unsigned(560, 12), 1159 => to_unsigned(4093, 12), 1160 => to_unsigned(2231, 12), 1161 => to_unsigned(3734, 12), 1162 => to_unsigned(3646, 12), 1163 => to_unsigned(479, 12), 1164 => to_unsigned(1849, 12), 1165 => to_unsigned(2773, 12), 1166 => to_unsigned(2338, 12), 1167 => to_unsigned(2999, 12), 1168 => to_unsigned(3881, 12), 1169 => to_unsigned(704, 12), 1170 => to_unsigned(2347, 12), 1171 => to_unsigned(11, 12), 1172 => to_unsigned(1160, 12), 1173 => to_unsigned(2967, 12), 1174 => to_unsigned(568, 12), 1175 => to_unsigned(4053, 12), 1176 => to_unsigned(2041, 12), 1177 => to_unsigned(1592, 12), 1178 => to_unsigned(3312, 12), 1179 => to_unsigned(1335, 12), 1180 => to_unsigned(1902, 12), 1181 => to_unsigned(1117, 12), 1182 => to_unsigned(381, 12), 1183 => to_unsigned(3208, 12), 1184 => to_unsigned(2325, 12), 1185 => to_unsigned(2936, 12), 1186 => to_unsigned(2292, 12), 1187 => to_unsigned(2764, 12), 1188 => to_unsigned(3565, 12), 1189 => to_unsigned(2731, 12), 1190 => to_unsigned(3465, 12), 1191 => to_unsigned(2299, 12), 1192 => to_unsigned(203, 12), 1193 => to_unsigned(2081, 12), 1194 => to_unsigned(45, 12), 1195 => to_unsigned(2025, 12), 1196 => to_unsigned(2099, 12), 1197 => to_unsigned(1776, 12), 1198 => to_unsigned(3800, 12), 1199 => to_unsigned(2375, 12), 1200 => to_unsigned(3797, 12), 1201 => to_unsigned(3869, 12), 1202 => to_unsigned(3818, 12), 1203 => to_unsigned(2279, 12), 1204 => to_unsigned(1382, 12), 1205 => to_unsigned(3031, 12), 1206 => to_unsigned(2114, 12), 1207 => to_unsigned(3242, 12), 1208 => to_unsigned(37, 12), 1209 => to_unsigned(883, 12), 1210 => to_unsigned(753, 12), 1211 => to_unsigned(3398, 12), 1212 => to_unsigned(916, 12), 1213 => to_unsigned(3121, 12), 1214 => to_unsigned(3812, 12), 1215 => to_unsigned(1574, 12), 1216 => to_unsigned(2773, 12), 1217 => to_unsigned(681, 12), 1218 => to_unsigned(2429, 12), 1219 => to_unsigned(1361, 12), 1220 => to_unsigned(2428, 12), 1221 => to_unsigned(160, 12), 1222 => to_unsigned(47, 12), 1223 => to_unsigned(594, 12), 1224 => to_unsigned(2843, 12), 1225 => to_unsigned(1867, 12), 1226 => to_unsigned(1749, 12), 1227 => to_unsigned(328, 12), 1228 => to_unsigned(574, 12), 1229 => to_unsigned(3927, 12), 1230 => to_unsigned(3752, 12), 1231 => to_unsigned(211, 12), 1232 => to_unsigned(660, 12), 1233 => to_unsigned(2779, 12), 1234 => to_unsigned(3325, 12), 1235 => to_unsigned(902, 12), 1236 => to_unsigned(2985, 12), 1237 => to_unsigned(1116, 12), 1238 => to_unsigned(112, 12), 1239 => to_unsigned(1355, 12), 1240 => to_unsigned(6, 12), 1241 => to_unsigned(3408, 12), 1242 => to_unsigned(671, 12), 1243 => to_unsigned(1965, 12), 1244 => to_unsigned(4039, 12), 1245 => to_unsigned(420, 12), 1246 => to_unsigned(3097, 12), 1247 => to_unsigned(2589, 12), 1248 => to_unsigned(502, 12), 1249 => to_unsigned(1150, 12), 1250 => to_unsigned(3711, 12), 1251 => to_unsigned(3502, 12), 1252 => to_unsigned(581, 12), 1253 => to_unsigned(2233, 12), 1254 => to_unsigned(1215, 12), 1255 => to_unsigned(2632, 12), 1256 => to_unsigned(2372, 12), 1257 => to_unsigned(1313, 12), 1258 => to_unsigned(421, 12), 1259 => to_unsigned(2945, 12), 1260 => to_unsigned(1687, 12), 1261 => to_unsigned(3121, 12), 1262 => to_unsigned(524, 12), 1263 => to_unsigned(2049, 12), 1264 => to_unsigned(2631, 12), 1265 => to_unsigned(1372, 12), 1266 => to_unsigned(3720, 12), 1267 => to_unsigned(3246, 12), 1268 => to_unsigned(2980, 12), 1269 => to_unsigned(816, 12), 1270 => to_unsigned(2488, 12), 1271 => to_unsigned(2217, 12), 1272 => to_unsigned(2648, 12), 1273 => to_unsigned(3648, 12), 1274 => to_unsigned(3810, 12), 1275 => to_unsigned(2093, 12), 1276 => to_unsigned(429, 12), 1277 => to_unsigned(3343, 12), 1278 => to_unsigned(551, 12), 1279 => to_unsigned(2818, 12), 1280 => to_unsigned(810, 12), 1281 => to_unsigned(2315, 12), 1282 => to_unsigned(2927, 12), 1283 => to_unsigned(3012, 12), 1284 => to_unsigned(1887, 12), 1285 => to_unsigned(3566, 12), 1286 => to_unsigned(1734, 12), 1287 => to_unsigned(1724, 12), 1288 => to_unsigned(2498, 12), 1289 => to_unsigned(1081, 12), 1290 => to_unsigned(2762, 12), 1291 => to_unsigned(3556, 12), 1292 => to_unsigned(170, 12), 1293 => to_unsigned(1709, 12), 1294 => to_unsigned(2769, 12), 1295 => to_unsigned(110, 12), 1296 => to_unsigned(1484, 12), 1297 => to_unsigned(232, 12), 1298 => to_unsigned(3857, 12), 1299 => to_unsigned(4015, 12), 1300 => to_unsigned(693, 12), 1301 => to_unsigned(391, 12), 1302 => to_unsigned(1867, 12), 1303 => to_unsigned(3482, 12), 1304 => to_unsigned(2326, 12), 1305 => to_unsigned(3300, 12), 1306 => to_unsigned(2673, 12), 1307 => to_unsigned(3547, 12), 1308 => to_unsigned(2684, 12), 1309 => to_unsigned(2124, 12), 1310 => to_unsigned(3271, 12), 1311 => to_unsigned(4050, 12), 1312 => to_unsigned(831, 12), 1313 => to_unsigned(593, 12), 1314 => to_unsigned(1590, 12), 1315 => to_unsigned(3207, 12), 1316 => to_unsigned(182, 12), 1317 => to_unsigned(3271, 12), 1318 => to_unsigned(904, 12), 1319 => to_unsigned(3156, 12), 1320 => to_unsigned(3633, 12), 1321 => to_unsigned(11, 12), 1322 => to_unsigned(2520, 12), 1323 => to_unsigned(1148, 12), 1324 => to_unsigned(3506, 12), 1325 => to_unsigned(410, 12), 1326 => to_unsigned(1805, 12), 1327 => to_unsigned(2160, 12), 1328 => to_unsigned(1580, 12), 1329 => to_unsigned(2188, 12), 1330 => to_unsigned(1611, 12), 1331 => to_unsigned(3278, 12), 1332 => to_unsigned(2323, 12), 1333 => to_unsigned(1186, 12), 1334 => to_unsigned(786, 12), 1335 => to_unsigned(2662, 12), 1336 => to_unsigned(3004, 12), 1337 => to_unsigned(1473, 12), 1338 => to_unsigned(3615, 12), 1339 => to_unsigned(1605, 12), 1340 => to_unsigned(1331, 12), 1341 => to_unsigned(3303, 12), 1342 => to_unsigned(1264, 12), 1343 => to_unsigned(904, 12), 1344 => to_unsigned(416, 12), 1345 => to_unsigned(1146, 12), 1346 => to_unsigned(2310, 12), 1347 => to_unsigned(1953, 12), 1348 => to_unsigned(3584, 12), 1349 => to_unsigned(2682, 12), 1350 => to_unsigned(131, 12), 1351 => to_unsigned(2111, 12), 1352 => to_unsigned(1531, 12), 1353 => to_unsigned(1449, 12), 1354 => to_unsigned(181, 12), 1355 => to_unsigned(3887, 12), 1356 => to_unsigned(570, 12), 1357 => to_unsigned(965, 12), 1358 => to_unsigned(44, 12), 1359 => to_unsigned(3707, 12), 1360 => to_unsigned(3170, 12), 1361 => to_unsigned(385, 12), 1362 => to_unsigned(1127, 12), 1363 => to_unsigned(3723, 12), 1364 => to_unsigned(754, 12), 1365 => to_unsigned(3981, 12), 1366 => to_unsigned(3596, 12), 1367 => to_unsigned(76, 12), 1368 => to_unsigned(1041, 12), 1369 => to_unsigned(443, 12), 1370 => to_unsigned(2473, 12), 1371 => to_unsigned(2356, 12), 1372 => to_unsigned(3417, 12), 1373 => to_unsigned(235, 12), 1374 => to_unsigned(1315, 12), 1375 => to_unsigned(3738, 12), 1376 => to_unsigned(311, 12), 1377 => to_unsigned(446, 12), 1378 => to_unsigned(2018, 12), 1379 => to_unsigned(693, 12), 1380 => to_unsigned(2376, 12), 1381 => to_unsigned(2218, 12), 1382 => to_unsigned(455, 12), 1383 => to_unsigned(1037, 12), 1384 => to_unsigned(392, 12), 1385 => to_unsigned(3610, 12), 1386 => to_unsigned(83, 12), 1387 => to_unsigned(2735, 12), 1388 => to_unsigned(2419, 12), 1389 => to_unsigned(2745, 12), 1390 => to_unsigned(2462, 12), 1391 => to_unsigned(1227, 12), 1392 => to_unsigned(3766, 12), 1393 => to_unsigned(3699, 12), 1394 => to_unsigned(2488, 12), 1395 => to_unsigned(2097, 12), 1396 => to_unsigned(995, 12), 1397 => to_unsigned(3731, 12), 1398 => to_unsigned(150, 12), 1399 => to_unsigned(3684, 12), 1400 => to_unsigned(2963, 12), 1401 => to_unsigned(1908, 12), 1402 => to_unsigned(2991, 12), 1403 => to_unsigned(2482, 12), 1404 => to_unsigned(1506, 12), 1405 => to_unsigned(3067, 12), 1406 => to_unsigned(3145, 12), 1407 => to_unsigned(1323, 12), 1408 => to_unsigned(2066, 12), 1409 => to_unsigned(1588, 12), 1410 => to_unsigned(1132, 12), 1411 => to_unsigned(1541, 12), 1412 => to_unsigned(1562, 12), 1413 => to_unsigned(1295, 12), 1414 => to_unsigned(1439, 12), 1415 => to_unsigned(11, 12), 1416 => to_unsigned(3074, 12), 1417 => to_unsigned(2231, 12), 1418 => to_unsigned(2218, 12), 1419 => to_unsigned(1660, 12), 1420 => to_unsigned(1230, 12), 1421 => to_unsigned(652, 12), 1422 => to_unsigned(458, 12), 1423 => to_unsigned(2759, 12), 1424 => to_unsigned(1430, 12), 1425 => to_unsigned(55, 12), 1426 => to_unsigned(463, 12), 1427 => to_unsigned(948, 12), 1428 => to_unsigned(1347, 12), 1429 => to_unsigned(1999, 12), 1430 => to_unsigned(107, 12), 1431 => to_unsigned(1504, 12), 1432 => to_unsigned(1410, 12), 1433 => to_unsigned(1023, 12), 1434 => to_unsigned(4095, 12), 1435 => to_unsigned(3950, 12), 1436 => to_unsigned(1689, 12), 1437 => to_unsigned(2669, 12), 1438 => to_unsigned(1851, 12), 1439 => to_unsigned(1798, 12), 1440 => to_unsigned(909, 12), 1441 => to_unsigned(2414, 12), 1442 => to_unsigned(1740, 12), 1443 => to_unsigned(754, 12), 1444 => to_unsigned(3193, 12), 1445 => to_unsigned(2681, 12), 1446 => to_unsigned(2654, 12), 1447 => to_unsigned(3033, 12), 1448 => to_unsigned(3374, 12), 1449 => to_unsigned(3713, 12), 1450 => to_unsigned(2871, 12), 1451 => to_unsigned(79, 12), 1452 => to_unsigned(2483, 12), 1453 => to_unsigned(2504, 12), 1454 => to_unsigned(2668, 12), 1455 => to_unsigned(219, 12), 1456 => to_unsigned(64, 12), 1457 => to_unsigned(3115, 12), 1458 => to_unsigned(36, 12), 1459 => to_unsigned(3387, 12), 1460 => to_unsigned(1116, 12), 1461 => to_unsigned(3370, 12), 1462 => to_unsigned(3499, 12), 1463 => to_unsigned(234, 12), 1464 => to_unsigned(211, 12), 1465 => to_unsigned(2850, 12), 1466 => to_unsigned(2885, 12), 1467 => to_unsigned(2146, 12), 1468 => to_unsigned(3362, 12), 1469 => to_unsigned(3009, 12), 1470 => to_unsigned(224, 12), 1471 => to_unsigned(768, 12), 1472 => to_unsigned(1599, 12), 1473 => to_unsigned(869, 12), 1474 => to_unsigned(130, 12), 1475 => to_unsigned(1151, 12), 1476 => to_unsigned(1605, 12), 1477 => to_unsigned(569, 12), 1478 => to_unsigned(2681, 12), 1479 => to_unsigned(3276, 12), 1480 => to_unsigned(1153, 12), 1481 => to_unsigned(775, 12), 1482 => to_unsigned(807, 12), 1483 => to_unsigned(2978, 12), 1484 => to_unsigned(876, 12), 1485 => to_unsigned(2399, 12), 1486 => to_unsigned(3800, 12), 1487 => to_unsigned(590, 12), 1488 => to_unsigned(1720, 12), 1489 => to_unsigned(1075, 12), 1490 => to_unsigned(2930, 12), 1491 => to_unsigned(3551, 12), 1492 => to_unsigned(3446, 12), 1493 => to_unsigned(2837, 12), 1494 => to_unsigned(2003, 12), 1495 => to_unsigned(543, 12), 1496 => to_unsigned(3543, 12), 1497 => to_unsigned(1584, 12), 1498 => to_unsigned(2609, 12), 1499 => to_unsigned(4028, 12), 1500 => to_unsigned(3901, 12), 1501 => to_unsigned(3299, 12), 1502 => to_unsigned(2098, 12), 1503 => to_unsigned(2080, 12), 1504 => to_unsigned(2368, 12), 1505 => to_unsigned(1381, 12), 1506 => to_unsigned(276, 12), 1507 => to_unsigned(4040, 12), 1508 => to_unsigned(3453, 12), 1509 => to_unsigned(683, 12), 1510 => to_unsigned(1477, 12), 1511 => to_unsigned(1448, 12), 1512 => to_unsigned(3440, 12), 1513 => to_unsigned(3452, 12), 1514 => to_unsigned(1945, 12), 1515 => to_unsigned(3191, 12), 1516 => to_unsigned(4038, 12), 1517 => to_unsigned(3837, 12), 1518 => to_unsigned(274, 12), 1519 => to_unsigned(2519, 12), 1520 => to_unsigned(1093, 12), 1521 => to_unsigned(4042, 12), 1522 => to_unsigned(1891, 12), 1523 => to_unsigned(3893, 12), 1524 => to_unsigned(2354, 12), 1525 => to_unsigned(3348, 12), 1526 => to_unsigned(3580, 12), 1527 => to_unsigned(2112, 12), 1528 => to_unsigned(429, 12), 1529 => to_unsigned(2655, 12), 1530 => to_unsigned(2055, 12), 1531 => to_unsigned(592, 12), 1532 => to_unsigned(1635, 12), 1533 => to_unsigned(2661, 12), 1534 => to_unsigned(3409, 12), 1535 => to_unsigned(3006, 12), 1536 => to_unsigned(3255, 12), 1537 => to_unsigned(2896, 12), 1538 => to_unsigned(1940, 12), 1539 => to_unsigned(632, 12), 1540 => to_unsigned(3363, 12), 1541 => to_unsigned(163, 12), 1542 => to_unsigned(23, 12), 1543 => to_unsigned(1496, 12), 1544 => to_unsigned(1849, 12), 1545 => to_unsigned(138, 12), 1546 => to_unsigned(1685, 12), 1547 => to_unsigned(2644, 12), 1548 => to_unsigned(873, 12), 1549 => to_unsigned(2267, 12), 1550 => to_unsigned(2196, 12), 1551 => to_unsigned(2405, 12), 1552 => to_unsigned(3439, 12), 1553 => to_unsigned(2516, 12), 1554 => to_unsigned(594, 12), 1555 => to_unsigned(2067, 12), 1556 => to_unsigned(330, 12), 1557 => to_unsigned(1095, 12), 1558 => to_unsigned(1450, 12), 1559 => to_unsigned(1471, 12), 1560 => to_unsigned(3689, 12), 1561 => to_unsigned(479, 12), 1562 => to_unsigned(2510, 12), 1563 => to_unsigned(349, 12), 1564 => to_unsigned(2739, 12), 1565 => to_unsigned(3187, 12), 1566 => to_unsigned(31, 12), 1567 => to_unsigned(1953, 12), 1568 => to_unsigned(990, 12), 1569 => to_unsigned(2151, 12), 1570 => to_unsigned(374, 12), 1571 => to_unsigned(2027, 12), 1572 => to_unsigned(417, 12), 1573 => to_unsigned(635, 12), 1574 => to_unsigned(29, 12), 1575 => to_unsigned(1928, 12), 1576 => to_unsigned(3491, 12), 1577 => to_unsigned(646, 12), 1578 => to_unsigned(3400, 12), 1579 => to_unsigned(2303, 12), 1580 => to_unsigned(2413, 12), 1581 => to_unsigned(2210, 12), 1582 => to_unsigned(202, 12), 1583 => to_unsigned(3518, 12), 1584 => to_unsigned(954, 12), 1585 => to_unsigned(244, 12), 1586 => to_unsigned(3890, 12), 1587 => to_unsigned(614, 12), 1588 => to_unsigned(1816, 12), 1589 => to_unsigned(2621, 12), 1590 => to_unsigned(921, 12), 1591 => to_unsigned(1246, 12), 1592 => to_unsigned(3657, 12), 1593 => to_unsigned(692, 12), 1594 => to_unsigned(670, 12), 1595 => to_unsigned(2347, 12), 1596 => to_unsigned(3554, 12), 1597 => to_unsigned(1179, 12), 1598 => to_unsigned(3327, 12), 1599 => to_unsigned(775, 12), 1600 => to_unsigned(409, 12), 1601 => to_unsigned(2000, 12), 1602 => to_unsigned(2740, 12), 1603 => to_unsigned(2868, 12), 1604 => to_unsigned(2412, 12), 1605 => to_unsigned(1986, 12), 1606 => to_unsigned(2486, 12), 1607 => to_unsigned(3486, 12), 1608 => to_unsigned(2820, 12), 1609 => to_unsigned(584, 12), 1610 => to_unsigned(2928, 12), 1611 => to_unsigned(2836, 12), 1612 => to_unsigned(431, 12), 1613 => to_unsigned(3297, 12), 1614 => to_unsigned(701, 12), 1615 => to_unsigned(2886, 12), 1616 => to_unsigned(1527, 12), 1617 => to_unsigned(3869, 12), 1618 => to_unsigned(1478, 12), 1619 => to_unsigned(1273, 12), 1620 => to_unsigned(676, 12), 1621 => to_unsigned(2522, 12), 1622 => to_unsigned(545, 12), 1623 => to_unsigned(468, 12), 1624 => to_unsigned(975, 12), 1625 => to_unsigned(1848, 12), 1626 => to_unsigned(2571, 12), 1627 => to_unsigned(1551, 12), 1628 => to_unsigned(3705, 12), 1629 => to_unsigned(2794, 12), 1630 => to_unsigned(2453, 12), 1631 => to_unsigned(1115, 12), 1632 => to_unsigned(1067, 12), 1633 => to_unsigned(1874, 12), 1634 => to_unsigned(650, 12), 1635 => to_unsigned(2316, 12), 1636 => to_unsigned(1712, 12), 1637 => to_unsigned(2806, 12), 1638 => to_unsigned(1398, 12), 1639 => to_unsigned(626, 12), 1640 => to_unsigned(2050, 12), 1641 => to_unsigned(2507, 12), 1642 => to_unsigned(390, 12), 1643 => to_unsigned(3937, 12), 1644 => to_unsigned(215, 12), 1645 => to_unsigned(3957, 12), 1646 => to_unsigned(1257, 12), 1647 => to_unsigned(1246, 12), 1648 => to_unsigned(2237, 12), 1649 => to_unsigned(703, 12), 1650 => to_unsigned(1690, 12), 1651 => to_unsigned(248, 12), 1652 => to_unsigned(3114, 12), 1653 => to_unsigned(3800, 12), 1654 => to_unsigned(1923, 12), 1655 => to_unsigned(1108, 12), 1656 => to_unsigned(2391, 12), 1657 => to_unsigned(2431, 12), 1658 => to_unsigned(843, 12), 1659 => to_unsigned(2564, 12), 1660 => to_unsigned(1973, 12), 1661 => to_unsigned(683, 12), 1662 => to_unsigned(3826, 12), 1663 => to_unsigned(3398, 12), 1664 => to_unsigned(1245, 12), 1665 => to_unsigned(74, 12), 1666 => to_unsigned(88, 12), 1667 => to_unsigned(2047, 12), 1668 => to_unsigned(1210, 12), 1669 => to_unsigned(2261, 12), 1670 => to_unsigned(2761, 12), 1671 => to_unsigned(934, 12), 1672 => to_unsigned(1354, 12), 1673 => to_unsigned(3273, 12), 1674 => to_unsigned(1317, 12), 1675 => to_unsigned(587, 12), 1676 => to_unsigned(3603, 12), 1677 => to_unsigned(2532, 12), 1678 => to_unsigned(2863, 12), 1679 => to_unsigned(821, 12), 1680 => to_unsigned(572, 12), 1681 => to_unsigned(3314, 12), 1682 => to_unsigned(3502, 12), 1683 => to_unsigned(506, 12), 1684 => to_unsigned(157, 12), 1685 => to_unsigned(28, 12), 1686 => to_unsigned(1959, 12), 1687 => to_unsigned(2758, 12), 1688 => to_unsigned(1410, 12), 1689 => to_unsigned(1545, 12), 1690 => to_unsigned(2275, 12), 1691 => to_unsigned(3080, 12), 1692 => to_unsigned(520, 12), 1693 => to_unsigned(3331, 12), 1694 => to_unsigned(2256, 12), 1695 => to_unsigned(2504, 12), 1696 => to_unsigned(1225, 12), 1697 => to_unsigned(1051, 12), 1698 => to_unsigned(3830, 12), 1699 => to_unsigned(279, 12), 1700 => to_unsigned(2813, 12), 1701 => to_unsigned(244, 12), 1702 => to_unsigned(1307, 12), 1703 => to_unsigned(2106, 12), 1704 => to_unsigned(3866, 12), 1705 => to_unsigned(2203, 12), 1706 => to_unsigned(64, 12), 1707 => to_unsigned(3905, 12), 1708 => to_unsigned(3990, 12), 1709 => to_unsigned(3871, 12), 1710 => to_unsigned(658, 12), 1711 => to_unsigned(884, 12), 1712 => to_unsigned(1561, 12), 1713 => to_unsigned(3652, 12), 1714 => to_unsigned(2480, 12), 1715 => to_unsigned(2636, 12), 1716 => to_unsigned(1788, 12), 1717 => to_unsigned(2994, 12), 1718 => to_unsigned(3712, 12), 1719 => to_unsigned(1452, 12), 1720 => to_unsigned(2681, 12), 1721 => to_unsigned(4051, 12), 1722 => to_unsigned(3701, 12), 1723 => to_unsigned(2939, 12), 1724 => to_unsigned(3066, 12), 1725 => to_unsigned(2102, 12), 1726 => to_unsigned(1439, 12), 1727 => to_unsigned(772, 12), 1728 => to_unsigned(3175, 12), 1729 => to_unsigned(105, 12), 1730 => to_unsigned(729, 12), 1731 => to_unsigned(2605, 12), 1732 => to_unsigned(348, 12), 1733 => to_unsigned(1813, 12), 1734 => to_unsigned(2726, 12), 1735 => to_unsigned(919, 12), 1736 => to_unsigned(439, 12), 1737 => to_unsigned(2334, 12), 1738 => to_unsigned(740, 12), 1739 => to_unsigned(2784, 12), 1740 => to_unsigned(1451, 12), 1741 => to_unsigned(3044, 12), 1742 => to_unsigned(143, 12), 1743 => to_unsigned(3612, 12), 1744 => to_unsigned(1271, 12), 1745 => to_unsigned(1673, 12), 1746 => to_unsigned(1958, 12), 1747 => to_unsigned(3565, 12), 1748 => to_unsigned(1613, 12), 1749 => to_unsigned(3866, 12), 1750 => to_unsigned(1149, 12), 1751 => to_unsigned(3523, 12), 1752 => to_unsigned(2411, 12), 1753 => to_unsigned(1831, 12), 1754 => to_unsigned(2659, 12), 1755 => to_unsigned(3096, 12), 1756 => to_unsigned(3555, 12), 1757 => to_unsigned(1305, 12), 1758 => to_unsigned(2404, 12), 1759 => to_unsigned(1865, 12), 1760 => to_unsigned(280, 12), 1761 => to_unsigned(472, 12), 1762 => to_unsigned(2321, 12), 1763 => to_unsigned(802, 12), 1764 => to_unsigned(831, 12), 1765 => to_unsigned(1850, 12), 1766 => to_unsigned(2581, 12), 1767 => to_unsigned(3669, 12), 1768 => to_unsigned(3320, 12), 1769 => to_unsigned(279, 12), 1770 => to_unsigned(1133, 12), 1771 => to_unsigned(1354, 12), 1772 => to_unsigned(2703, 12), 1773 => to_unsigned(2789, 12), 1774 => to_unsigned(421, 12), 1775 => to_unsigned(2142, 12), 1776 => to_unsigned(3718, 12), 1777 => to_unsigned(2526, 12), 1778 => to_unsigned(742, 12), 1779 => to_unsigned(4093, 12), 1780 => to_unsigned(2977, 12), 1781 => to_unsigned(2888, 12), 1782 => to_unsigned(3831, 12), 1783 => to_unsigned(459, 12), 1784 => to_unsigned(3743, 12), 1785 => to_unsigned(362, 12), 1786 => to_unsigned(2293, 12), 1787 => to_unsigned(3101, 12), 1788 => to_unsigned(2174, 12), 1789 => to_unsigned(3546, 12), 1790 => to_unsigned(3749, 12), 1791 => to_unsigned(265, 12), 1792 => to_unsigned(4063, 12), 1793 => to_unsigned(1151, 12), 1794 => to_unsigned(2741, 12), 1795 => to_unsigned(3665, 12), 1796 => to_unsigned(2009, 12), 1797 => to_unsigned(1042, 12), 1798 => to_unsigned(1506, 12), 1799 => to_unsigned(1864, 12), 1800 => to_unsigned(3018, 12), 1801 => to_unsigned(1664, 12), 1802 => to_unsigned(161, 12), 1803 => to_unsigned(1117, 12), 1804 => to_unsigned(971, 12), 1805 => to_unsigned(2914, 12), 1806 => to_unsigned(1022, 12), 1807 => to_unsigned(977, 12), 1808 => to_unsigned(331, 12), 1809 => to_unsigned(975, 12), 1810 => to_unsigned(485, 12), 1811 => to_unsigned(1527, 12), 1812 => to_unsigned(1361, 12), 1813 => to_unsigned(837, 12), 1814 => to_unsigned(1291, 12), 1815 => to_unsigned(1794, 12), 1816 => to_unsigned(3961, 12), 1817 => to_unsigned(1946, 12), 1818 => to_unsigned(4008, 12), 1819 => to_unsigned(2073, 12), 1820 => to_unsigned(3659, 12), 1821 => to_unsigned(3431, 12), 1822 => to_unsigned(2169, 12), 1823 => to_unsigned(2444, 12), 1824 => to_unsigned(3798, 12), 1825 => to_unsigned(2388, 12), 1826 => to_unsigned(1440, 12), 1827 => to_unsigned(57, 12), 1828 => to_unsigned(1590, 12), 1829 => to_unsigned(3073, 12), 1830 => to_unsigned(2613, 12), 1831 => to_unsigned(1811, 12), 1832 => to_unsigned(1614, 12), 1833 => to_unsigned(3837, 12), 1834 => to_unsigned(2091, 12), 1835 => to_unsigned(2131, 12), 1836 => to_unsigned(3273, 12), 1837 => to_unsigned(2993, 12), 1838 => to_unsigned(4004, 12), 1839 => to_unsigned(34, 12), 1840 => to_unsigned(390, 12), 1841 => to_unsigned(763, 12), 1842 => to_unsigned(3962, 12), 1843 => to_unsigned(1045, 12), 1844 => to_unsigned(2981, 12), 1845 => to_unsigned(4050, 12), 1846 => to_unsigned(2896, 12), 1847 => to_unsigned(1222, 12), 1848 => to_unsigned(463, 12), 1849 => to_unsigned(1135, 12), 1850 => to_unsigned(1958, 12), 1851 => to_unsigned(617, 12), 1852 => to_unsigned(3149, 12), 1853 => to_unsigned(3001, 12), 1854 => to_unsigned(2836, 12), 1855 => to_unsigned(769, 12), 1856 => to_unsigned(2480, 12), 1857 => to_unsigned(2478, 12), 1858 => to_unsigned(3381, 12), 1859 => to_unsigned(542, 12), 1860 => to_unsigned(3361, 12), 1861 => to_unsigned(2887, 12), 1862 => to_unsigned(1203, 12), 1863 => to_unsigned(2355, 12), 1864 => to_unsigned(2350, 12), 1865 => to_unsigned(628, 12), 1866 => to_unsigned(1374, 12), 1867 => to_unsigned(1877, 12), 1868 => to_unsigned(3630, 12), 1869 => to_unsigned(963, 12), 1870 => to_unsigned(3304, 12), 1871 => to_unsigned(665, 12), 1872 => to_unsigned(3066, 12), 1873 => to_unsigned(753, 12), 1874 => to_unsigned(2024, 12), 1875 => to_unsigned(2857, 12), 1876 => to_unsigned(342, 12), 1877 => to_unsigned(3777, 12), 1878 => to_unsigned(1635, 12), 1879 => to_unsigned(2624, 12), 1880 => to_unsigned(2083, 12), 1881 => to_unsigned(1612, 12), 1882 => to_unsigned(1302, 12), 1883 => to_unsigned(829, 12), 1884 => to_unsigned(2493, 12), 1885 => to_unsigned(916, 12), 1886 => to_unsigned(2024, 12), 1887 => to_unsigned(2151, 12), 1888 => to_unsigned(558, 12), 1889 => to_unsigned(3632, 12), 1890 => to_unsigned(92, 12), 1891 => to_unsigned(3149, 12), 1892 => to_unsigned(2949, 12), 1893 => to_unsigned(3090, 12), 1894 => to_unsigned(2317, 12), 1895 => to_unsigned(326, 12), 1896 => to_unsigned(3166, 12), 1897 => to_unsigned(1349, 12), 1898 => to_unsigned(1004, 12), 1899 => to_unsigned(1366, 12), 1900 => to_unsigned(1953, 12), 1901 => to_unsigned(3908, 12), 1902 => to_unsigned(782, 12), 1903 => to_unsigned(1214, 12), 1904 => to_unsigned(3758, 12), 1905 => to_unsigned(3749, 12), 1906 => to_unsigned(460, 12), 1907 => to_unsigned(43, 12), 1908 => to_unsigned(3526, 12), 1909 => to_unsigned(2600, 12), 1910 => to_unsigned(1435, 12), 1911 => to_unsigned(1323, 12), 1912 => to_unsigned(1923, 12), 1913 => to_unsigned(17, 12), 1914 => to_unsigned(47, 12), 1915 => to_unsigned(2992, 12), 1916 => to_unsigned(1228, 12), 1917 => to_unsigned(3503, 12), 1918 => to_unsigned(2847, 12), 1919 => to_unsigned(271, 12), 1920 => to_unsigned(3537, 12), 1921 => to_unsigned(2315, 12), 1922 => to_unsigned(1833, 12), 1923 => to_unsigned(2561, 12), 1924 => to_unsigned(2838, 12), 1925 => to_unsigned(102, 12), 1926 => to_unsigned(2103, 12), 1927 => to_unsigned(2821, 12), 1928 => to_unsigned(3947, 12), 1929 => to_unsigned(1987, 12), 1930 => to_unsigned(2321, 12), 1931 => to_unsigned(1841, 12), 1932 => to_unsigned(3440, 12), 1933 => to_unsigned(3864, 12), 1934 => to_unsigned(3259, 12), 1935 => to_unsigned(1715, 12), 1936 => to_unsigned(1617, 12), 1937 => to_unsigned(1109, 12), 1938 => to_unsigned(2362, 12), 1939 => to_unsigned(1280, 12), 1940 => to_unsigned(1618, 12), 1941 => to_unsigned(2001, 12), 1942 => to_unsigned(540, 12), 1943 => to_unsigned(15, 12), 1944 => to_unsigned(3684, 12), 1945 => to_unsigned(2532, 12), 1946 => to_unsigned(2348, 12), 1947 => to_unsigned(351, 12), 1948 => to_unsigned(3777, 12), 1949 => to_unsigned(2318, 12), 1950 => to_unsigned(3104, 12), 1951 => to_unsigned(2096, 12), 1952 => to_unsigned(3458, 12), 1953 => to_unsigned(2155, 12), 1954 => to_unsigned(916, 12), 1955 => to_unsigned(1672, 12), 1956 => to_unsigned(1937, 12), 1957 => to_unsigned(54, 12), 1958 => to_unsigned(2131, 12), 1959 => to_unsigned(3698, 12), 1960 => to_unsigned(674, 12), 1961 => to_unsigned(2632, 12), 1962 => to_unsigned(599, 12), 1963 => to_unsigned(1110, 12), 1964 => to_unsigned(89, 12), 1965 => to_unsigned(2409, 12), 1966 => to_unsigned(3903, 12), 1967 => to_unsigned(1741, 12), 1968 => to_unsigned(3448, 12), 1969 => to_unsigned(4015, 12), 1970 => to_unsigned(1294, 12), 1971 => to_unsigned(696, 12), 1972 => to_unsigned(3752, 12), 1973 => to_unsigned(1718, 12), 1974 => to_unsigned(3664, 12), 1975 => to_unsigned(3878, 12), 1976 => to_unsigned(3097, 12), 1977 => to_unsigned(441, 12), 1978 => to_unsigned(3288, 12), 1979 => to_unsigned(337, 12), 1980 => to_unsigned(3135, 12), 1981 => to_unsigned(1138, 12), 1982 => to_unsigned(3237, 12), 1983 => to_unsigned(1758, 12), 1984 => to_unsigned(1985, 12), 1985 => to_unsigned(2825, 12), 1986 => to_unsigned(621, 12), 1987 => to_unsigned(3899, 12), 1988 => to_unsigned(750, 12), 1989 => to_unsigned(2433, 12), 1990 => to_unsigned(2328, 12), 1991 => to_unsigned(1445, 12), 1992 => to_unsigned(1912, 12), 1993 => to_unsigned(1560, 12), 1994 => to_unsigned(1084, 12), 1995 => to_unsigned(2001, 12), 1996 => to_unsigned(1255, 12), 1997 => to_unsigned(3813, 12), 1998 => to_unsigned(3526, 12), 1999 => to_unsigned(2283, 12), 2000 => to_unsigned(3534, 12), 2001 => to_unsigned(1240, 12), 2002 => to_unsigned(488, 12), 2003 => to_unsigned(4055, 12), 2004 => to_unsigned(2597, 12), 2005 => to_unsigned(2588, 12), 2006 => to_unsigned(130, 12), 2007 => to_unsigned(724, 12), 2008 => to_unsigned(440, 12), 2009 => to_unsigned(2511, 12), 2010 => to_unsigned(1821, 12), 2011 => to_unsigned(1743, 12), 2012 => to_unsigned(3080, 12), 2013 => to_unsigned(2025, 12), 2014 => to_unsigned(1298, 12), 2015 => to_unsigned(1887, 12), 2016 => to_unsigned(3784, 12), 2017 => to_unsigned(699, 12), 2018 => to_unsigned(222, 12), 2019 => to_unsigned(687, 12), 2020 => to_unsigned(3199, 12), 2021 => to_unsigned(3045, 12), 2022 => to_unsigned(2790, 12), 2023 => to_unsigned(592, 12), 2024 => to_unsigned(2437, 12), 2025 => to_unsigned(2220, 12), 2026 => to_unsigned(3670, 12), 2027 => to_unsigned(1525, 12), 2028 => to_unsigned(2596, 12), 2029 => to_unsigned(3886, 12), 2030 => to_unsigned(4086, 12), 2031 => to_unsigned(1805, 12), 2032 => to_unsigned(1137, 12), 2033 => to_unsigned(143, 12), 2034 => to_unsigned(2416, 12), 2035 => to_unsigned(2504, 12), 2036 => to_unsigned(3103, 12), 2037 => to_unsigned(2009, 12), 2038 => to_unsigned(3117, 12), 2039 => to_unsigned(21, 12), 2040 => to_unsigned(3664, 12), 2041 => to_unsigned(1186, 12), 2042 => to_unsigned(649, 12), 2043 => to_unsigned(2441, 12), 2044 => to_unsigned(3421, 12), 2045 => to_unsigned(1822, 12), 2046 => to_unsigned(3338, 12), 2047 => to_unsigned(2022, 12)),
            7 => (0 => to_unsigned(2979, 12), 1 => to_unsigned(376, 12), 2 => to_unsigned(1976, 12), 3 => to_unsigned(1582, 12), 4 => to_unsigned(3166, 12), 5 => to_unsigned(3227, 12), 6 => to_unsigned(2485, 12), 7 => to_unsigned(1604, 12), 8 => to_unsigned(1233, 12), 9 => to_unsigned(1721, 12), 10 => to_unsigned(301, 12), 11 => to_unsigned(2932, 12), 12 => to_unsigned(1290, 12), 13 => to_unsigned(684, 12), 14 => to_unsigned(3223, 12), 15 => to_unsigned(490, 12), 16 => to_unsigned(81, 12), 17 => to_unsigned(2855, 12), 18 => to_unsigned(1784, 12), 19 => to_unsigned(189, 12), 20 => to_unsigned(2486, 12), 21 => to_unsigned(3431, 12), 22 => to_unsigned(3994, 12), 23 => to_unsigned(2165, 12), 24 => to_unsigned(1721, 12), 25 => to_unsigned(2905, 12), 26 => to_unsigned(4018, 12), 27 => to_unsigned(102, 12), 28 => to_unsigned(219, 12), 29 => to_unsigned(1786, 12), 30 => to_unsigned(1047, 12), 31 => to_unsigned(545, 12), 32 => to_unsigned(2846, 12), 33 => to_unsigned(2856, 12), 34 => to_unsigned(420, 12), 35 => to_unsigned(987, 12), 36 => to_unsigned(1401, 12), 37 => to_unsigned(2384, 12), 38 => to_unsigned(2259, 12), 39 => to_unsigned(3566, 12), 40 => to_unsigned(376, 12), 41 => to_unsigned(1406, 12), 42 => to_unsigned(3637, 12), 43 => to_unsigned(1177, 12), 44 => to_unsigned(4095, 12), 45 => to_unsigned(1416, 12), 46 => to_unsigned(3101, 12), 47 => to_unsigned(825, 12), 48 => to_unsigned(1359, 12), 49 => to_unsigned(2671, 12), 50 => to_unsigned(2112, 12), 51 => to_unsigned(1784, 12), 52 => to_unsigned(3763, 12), 53 => to_unsigned(444, 12), 54 => to_unsigned(1269, 12), 55 => to_unsigned(3127, 12), 56 => to_unsigned(1163, 12), 57 => to_unsigned(1522, 12), 58 => to_unsigned(2390, 12), 59 => to_unsigned(3298, 12), 60 => to_unsigned(2521, 12), 61 => to_unsigned(1960, 12), 62 => to_unsigned(1395, 12), 63 => to_unsigned(3296, 12), 64 => to_unsigned(2998, 12), 65 => to_unsigned(3805, 12), 66 => to_unsigned(196, 12), 67 => to_unsigned(1461, 12), 68 => to_unsigned(2215, 12), 69 => to_unsigned(56, 12), 70 => to_unsigned(1134, 12), 71 => to_unsigned(329, 12), 72 => to_unsigned(3395, 12), 73 => to_unsigned(3274, 12), 74 => to_unsigned(3967, 12), 75 => to_unsigned(150, 12), 76 => to_unsigned(284, 12), 77 => to_unsigned(1368, 12), 78 => to_unsigned(1021, 12), 79 => to_unsigned(2902, 12), 80 => to_unsigned(2564, 12), 81 => to_unsigned(852, 12), 82 => to_unsigned(2644, 12), 83 => to_unsigned(2750, 12), 84 => to_unsigned(1117, 12), 85 => to_unsigned(4076, 12), 86 => to_unsigned(3059, 12), 87 => to_unsigned(2159, 12), 88 => to_unsigned(3508, 12), 89 => to_unsigned(3214, 12), 90 => to_unsigned(452, 12), 91 => to_unsigned(3159, 12), 92 => to_unsigned(750, 12), 93 => to_unsigned(2563, 12), 94 => to_unsigned(1465, 12), 95 => to_unsigned(1970, 12), 96 => to_unsigned(983, 12), 97 => to_unsigned(3718, 12), 98 => to_unsigned(586, 12), 99 => to_unsigned(884, 12), 100 => to_unsigned(1486, 12), 101 => to_unsigned(1804, 12), 102 => to_unsigned(3218, 12), 103 => to_unsigned(3519, 12), 104 => to_unsigned(1112, 12), 105 => to_unsigned(3912, 12), 106 => to_unsigned(3356, 12), 107 => to_unsigned(3706, 12), 108 => to_unsigned(3478, 12), 109 => to_unsigned(1208, 12), 110 => to_unsigned(2312, 12), 111 => to_unsigned(210, 12), 112 => to_unsigned(2808, 12), 113 => to_unsigned(2701, 12), 114 => to_unsigned(511, 12), 115 => to_unsigned(2290, 12), 116 => to_unsigned(3995, 12), 117 => to_unsigned(2996, 12), 118 => to_unsigned(1714, 12), 119 => to_unsigned(4046, 12), 120 => to_unsigned(1807, 12), 121 => to_unsigned(905, 12), 122 => to_unsigned(3309, 12), 123 => to_unsigned(2226, 12), 124 => to_unsigned(1119, 12), 125 => to_unsigned(2443, 12), 126 => to_unsigned(3293, 12), 127 => to_unsigned(3913, 12), 128 => to_unsigned(2696, 12), 129 => to_unsigned(431, 12), 130 => to_unsigned(3713, 12), 131 => to_unsigned(281, 12), 132 => to_unsigned(2765, 12), 133 => to_unsigned(3894, 12), 134 => to_unsigned(1600, 12), 135 => to_unsigned(2425, 12), 136 => to_unsigned(3936, 12), 137 => to_unsigned(2633, 12), 138 => to_unsigned(2016, 12), 139 => to_unsigned(3250, 12), 140 => to_unsigned(2363, 12), 141 => to_unsigned(2099, 12), 142 => to_unsigned(2265, 12), 143 => to_unsigned(979, 12), 144 => to_unsigned(3390, 12), 145 => to_unsigned(2275, 12), 146 => to_unsigned(2297, 12), 147 => to_unsigned(4032, 12), 148 => to_unsigned(484, 12), 149 => to_unsigned(2418, 12), 150 => to_unsigned(3363, 12), 151 => to_unsigned(1113, 12), 152 => to_unsigned(2472, 12), 153 => to_unsigned(1070, 12), 154 => to_unsigned(3774, 12), 155 => to_unsigned(1053, 12), 156 => to_unsigned(3385, 12), 157 => to_unsigned(1254, 12), 158 => to_unsigned(3428, 12), 159 => to_unsigned(1079, 12), 160 => to_unsigned(1507, 12), 161 => to_unsigned(1757, 12), 162 => to_unsigned(2196, 12), 163 => to_unsigned(54, 12), 164 => to_unsigned(2424, 12), 165 => to_unsigned(1746, 12), 166 => to_unsigned(891, 12), 167 => to_unsigned(320, 12), 168 => to_unsigned(3329, 12), 169 => to_unsigned(2710, 12), 170 => to_unsigned(3305, 12), 171 => to_unsigned(687, 12), 172 => to_unsigned(1810, 12), 173 => to_unsigned(3186, 12), 174 => to_unsigned(2811, 12), 175 => to_unsigned(8, 12), 176 => to_unsigned(175, 12), 177 => to_unsigned(1648, 12), 178 => to_unsigned(1557, 12), 179 => to_unsigned(4014, 12), 180 => to_unsigned(466, 12), 181 => to_unsigned(4093, 12), 182 => to_unsigned(204, 12), 183 => to_unsigned(2447, 12), 184 => to_unsigned(3805, 12), 185 => to_unsigned(1786, 12), 186 => to_unsigned(3791, 12), 187 => to_unsigned(434, 12), 188 => to_unsigned(135, 12), 189 => to_unsigned(1175, 12), 190 => to_unsigned(3423, 12), 191 => to_unsigned(2542, 12), 192 => to_unsigned(2069, 12), 193 => to_unsigned(3175, 12), 194 => to_unsigned(1166, 12), 195 => to_unsigned(317, 12), 196 => to_unsigned(2969, 12), 197 => to_unsigned(3922, 12), 198 => to_unsigned(1860, 12), 199 => to_unsigned(495, 12), 200 => to_unsigned(2783, 12), 201 => to_unsigned(2657, 12), 202 => to_unsigned(3263, 12), 203 => to_unsigned(1350, 12), 204 => to_unsigned(289, 12), 205 => to_unsigned(1430, 12), 206 => to_unsigned(1788, 12), 207 => to_unsigned(1900, 12), 208 => to_unsigned(2249, 12), 209 => to_unsigned(3863, 12), 210 => to_unsigned(2903, 12), 211 => to_unsigned(2143, 12), 212 => to_unsigned(999, 12), 213 => to_unsigned(2543, 12), 214 => to_unsigned(2062, 12), 215 => to_unsigned(1449, 12), 216 => to_unsigned(1417, 12), 217 => to_unsigned(3300, 12), 218 => to_unsigned(1048, 12), 219 => to_unsigned(883, 12), 220 => to_unsigned(3907, 12), 221 => to_unsigned(1013, 12), 222 => to_unsigned(5, 12), 223 => to_unsigned(1855, 12), 224 => to_unsigned(3658, 12), 225 => to_unsigned(3942, 12), 226 => to_unsigned(412, 12), 227 => to_unsigned(3679, 12), 228 => to_unsigned(22, 12), 229 => to_unsigned(617, 12), 230 => to_unsigned(1526, 12), 231 => to_unsigned(2248, 12), 232 => to_unsigned(1278, 12), 233 => to_unsigned(3530, 12), 234 => to_unsigned(3413, 12), 235 => to_unsigned(1694, 12), 236 => to_unsigned(2002, 12), 237 => to_unsigned(57, 12), 238 => to_unsigned(3038, 12), 239 => to_unsigned(2652, 12), 240 => to_unsigned(3819, 12), 241 => to_unsigned(2591, 12), 242 => to_unsigned(478, 12), 243 => to_unsigned(672, 12), 244 => to_unsigned(2601, 12), 245 => to_unsigned(2168, 12), 246 => to_unsigned(796, 12), 247 => to_unsigned(3652, 12), 248 => to_unsigned(1514, 12), 249 => to_unsigned(833, 12), 250 => to_unsigned(3327, 12), 251 => to_unsigned(354, 12), 252 => to_unsigned(2530, 12), 253 => to_unsigned(1942, 12), 254 => to_unsigned(3312, 12), 255 => to_unsigned(237, 12), 256 => to_unsigned(1478, 12), 257 => to_unsigned(1897, 12), 258 => to_unsigned(2649, 12), 259 => to_unsigned(1388, 12), 260 => to_unsigned(3539, 12), 261 => to_unsigned(1022, 12), 262 => to_unsigned(905, 12), 263 => to_unsigned(994, 12), 264 => to_unsigned(3158, 12), 265 => to_unsigned(3942, 12), 266 => to_unsigned(3753, 12), 267 => to_unsigned(2363, 12), 268 => to_unsigned(3512, 12), 269 => to_unsigned(2229, 12), 270 => to_unsigned(156, 12), 271 => to_unsigned(919, 12), 272 => to_unsigned(2308, 12), 273 => to_unsigned(1405, 12), 274 => to_unsigned(2135, 12), 275 => to_unsigned(2151, 12), 276 => to_unsigned(529, 12), 277 => to_unsigned(1086, 12), 278 => to_unsigned(3208, 12), 279 => to_unsigned(3785, 12), 280 => to_unsigned(756, 12), 281 => to_unsigned(504, 12), 282 => to_unsigned(1729, 12), 283 => to_unsigned(1916, 12), 284 => to_unsigned(3551, 12), 285 => to_unsigned(1423, 12), 286 => to_unsigned(465, 12), 287 => to_unsigned(325, 12), 288 => to_unsigned(647, 12), 289 => to_unsigned(109, 12), 290 => to_unsigned(1730, 12), 291 => to_unsigned(2203, 12), 292 => to_unsigned(2914, 12), 293 => to_unsigned(3270, 12), 294 => to_unsigned(664, 12), 295 => to_unsigned(2034, 12), 296 => to_unsigned(356, 12), 297 => to_unsigned(1389, 12), 298 => to_unsigned(2572, 12), 299 => to_unsigned(4021, 12), 300 => to_unsigned(1549, 12), 301 => to_unsigned(2397, 12), 302 => to_unsigned(2029, 12), 303 => to_unsigned(1437, 12), 304 => to_unsigned(4049, 12), 305 => to_unsigned(2378, 12), 306 => to_unsigned(2728, 12), 307 => to_unsigned(2331, 12), 308 => to_unsigned(30, 12), 309 => to_unsigned(610, 12), 310 => to_unsigned(1176, 12), 311 => to_unsigned(2498, 12), 312 => to_unsigned(826, 12), 313 => to_unsigned(3465, 12), 314 => to_unsigned(1599, 12), 315 => to_unsigned(2021, 12), 316 => to_unsigned(262, 12), 317 => to_unsigned(364, 12), 318 => to_unsigned(3845, 12), 319 => to_unsigned(939, 12), 320 => to_unsigned(1395, 12), 321 => to_unsigned(102, 12), 322 => to_unsigned(1798, 12), 323 => to_unsigned(2679, 12), 324 => to_unsigned(3386, 12), 325 => to_unsigned(545, 12), 326 => to_unsigned(266, 12), 327 => to_unsigned(398, 12), 328 => to_unsigned(3314, 12), 329 => to_unsigned(3672, 12), 330 => to_unsigned(1929, 12), 331 => to_unsigned(2326, 12), 332 => to_unsigned(1960, 12), 333 => to_unsigned(1666, 12), 334 => to_unsigned(243, 12), 335 => to_unsigned(2770, 12), 336 => to_unsigned(3363, 12), 337 => to_unsigned(1960, 12), 338 => to_unsigned(3066, 12), 339 => to_unsigned(2890, 12), 340 => to_unsigned(672, 12), 341 => to_unsigned(4019, 12), 342 => to_unsigned(3734, 12), 343 => to_unsigned(149, 12), 344 => to_unsigned(3384, 12), 345 => to_unsigned(1706, 12), 346 => to_unsigned(3145, 12), 347 => to_unsigned(3954, 12), 348 => to_unsigned(4048, 12), 349 => to_unsigned(2794, 12), 350 => to_unsigned(683, 12), 351 => to_unsigned(855, 12), 352 => to_unsigned(885, 12), 353 => to_unsigned(475, 12), 354 => to_unsigned(2870, 12), 355 => to_unsigned(2810, 12), 356 => to_unsigned(727, 12), 357 => to_unsigned(1406, 12), 358 => to_unsigned(1133, 12), 359 => to_unsigned(2745, 12), 360 => to_unsigned(3406, 12), 361 => to_unsigned(1198, 12), 362 => to_unsigned(800, 12), 363 => to_unsigned(3304, 12), 364 => to_unsigned(1929, 12), 365 => to_unsigned(3552, 12), 366 => to_unsigned(790, 12), 367 => to_unsigned(3127, 12), 368 => to_unsigned(1380, 12), 369 => to_unsigned(493, 12), 370 => to_unsigned(1653, 12), 371 => to_unsigned(1455, 12), 372 => to_unsigned(798, 12), 373 => to_unsigned(1533, 12), 374 => to_unsigned(2056, 12), 375 => to_unsigned(2529, 12), 376 => to_unsigned(3694, 12), 377 => to_unsigned(1036, 12), 378 => to_unsigned(3809, 12), 379 => to_unsigned(2264, 12), 380 => to_unsigned(1704, 12), 381 => to_unsigned(36, 12), 382 => to_unsigned(2851, 12), 383 => to_unsigned(111, 12), 384 => to_unsigned(1158, 12), 385 => to_unsigned(3503, 12), 386 => to_unsigned(1305, 12), 387 => to_unsigned(3310, 12), 388 => to_unsigned(3506, 12), 389 => to_unsigned(2309, 12), 390 => to_unsigned(3239, 12), 391 => to_unsigned(425, 12), 392 => to_unsigned(3644, 12), 393 => to_unsigned(3705, 12), 394 => to_unsigned(191, 12), 395 => to_unsigned(3243, 12), 396 => to_unsigned(1945, 12), 397 => to_unsigned(433, 12), 398 => to_unsigned(2145, 12), 399 => to_unsigned(3130, 12), 400 => to_unsigned(759, 12), 401 => to_unsigned(3661, 12), 402 => to_unsigned(3955, 12), 403 => to_unsigned(3252, 12), 404 => to_unsigned(3629, 12), 405 => to_unsigned(1031, 12), 406 => to_unsigned(207, 12), 407 => to_unsigned(2451, 12), 408 => to_unsigned(2297, 12), 409 => to_unsigned(1532, 12), 410 => to_unsigned(307, 12), 411 => to_unsigned(2739, 12), 412 => to_unsigned(3746, 12), 413 => to_unsigned(1887, 12), 414 => to_unsigned(1690, 12), 415 => to_unsigned(1771, 12), 416 => to_unsigned(2229, 12), 417 => to_unsigned(836, 12), 418 => to_unsigned(1849, 12), 419 => to_unsigned(857, 12), 420 => to_unsigned(2418, 12), 421 => to_unsigned(3289, 12), 422 => to_unsigned(3988, 12), 423 => to_unsigned(1984, 12), 424 => to_unsigned(1463, 12), 425 => to_unsigned(1034, 12), 426 => to_unsigned(158, 12), 427 => to_unsigned(2801, 12), 428 => to_unsigned(715, 12), 429 => to_unsigned(2936, 12), 430 => to_unsigned(3356, 12), 431 => to_unsigned(2956, 12), 432 => to_unsigned(1397, 12), 433 => to_unsigned(818, 12), 434 => to_unsigned(2824, 12), 435 => to_unsigned(2565, 12), 436 => to_unsigned(2629, 12), 437 => to_unsigned(549, 12), 438 => to_unsigned(497, 12), 439 => to_unsigned(2506, 12), 440 => to_unsigned(2863, 12), 441 => to_unsigned(320, 12), 442 => to_unsigned(3828, 12), 443 => to_unsigned(1135, 12), 444 => to_unsigned(403, 12), 445 => to_unsigned(756, 12), 446 => to_unsigned(1971, 12), 447 => to_unsigned(2074, 12), 448 => to_unsigned(1677, 12), 449 => to_unsigned(920, 12), 450 => to_unsigned(1642, 12), 451 => to_unsigned(3858, 12), 452 => to_unsigned(1097, 12), 453 => to_unsigned(1340, 12), 454 => to_unsigned(2700, 12), 455 => to_unsigned(1051, 12), 456 => to_unsigned(2253, 12), 457 => to_unsigned(3848, 12), 458 => to_unsigned(3510, 12), 459 => to_unsigned(375, 12), 460 => to_unsigned(3810, 12), 461 => to_unsigned(1603, 12), 462 => to_unsigned(1030, 12), 463 => to_unsigned(206, 12), 464 => to_unsigned(1361, 12), 465 => to_unsigned(2633, 12), 466 => to_unsigned(2833, 12), 467 => to_unsigned(3796, 12), 468 => to_unsigned(3063, 12), 469 => to_unsigned(873, 12), 470 => to_unsigned(455, 12), 471 => to_unsigned(2062, 12), 472 => to_unsigned(1877, 12), 473 => to_unsigned(3296, 12), 474 => to_unsigned(2018, 12), 475 => to_unsigned(1329, 12), 476 => to_unsigned(1906, 12), 477 => to_unsigned(2179, 12), 478 => to_unsigned(228, 12), 479 => to_unsigned(2653, 12), 480 => to_unsigned(2425, 12), 481 => to_unsigned(1814, 12), 482 => to_unsigned(1551, 12), 483 => to_unsigned(1256, 12), 484 => to_unsigned(3937, 12), 485 => to_unsigned(3173, 12), 486 => to_unsigned(593, 12), 487 => to_unsigned(3150, 12), 488 => to_unsigned(3459, 12), 489 => to_unsigned(480, 12), 490 => to_unsigned(2361, 12), 491 => to_unsigned(400, 12), 492 => to_unsigned(229, 12), 493 => to_unsigned(1220, 12), 494 => to_unsigned(1400, 12), 495 => to_unsigned(691, 12), 496 => to_unsigned(2928, 12), 497 => to_unsigned(3551, 12), 498 => to_unsigned(2072, 12), 499 => to_unsigned(1661, 12), 500 => to_unsigned(2316, 12), 501 => to_unsigned(3607, 12), 502 => to_unsigned(2997, 12), 503 => to_unsigned(1421, 12), 504 => to_unsigned(300, 12), 505 => to_unsigned(2966, 12), 506 => to_unsigned(2743, 12), 507 => to_unsigned(2647, 12), 508 => to_unsigned(3031, 12), 509 => to_unsigned(2902, 12), 510 => to_unsigned(2386, 12), 511 => to_unsigned(3352, 12), 512 => to_unsigned(4089, 12), 513 => to_unsigned(1516, 12), 514 => to_unsigned(2636, 12), 515 => to_unsigned(639, 12), 516 => to_unsigned(2662, 12), 517 => to_unsigned(1390, 12), 518 => to_unsigned(523, 12), 519 => to_unsigned(909, 12), 520 => to_unsigned(1280, 12), 521 => to_unsigned(3135, 12), 522 => to_unsigned(527, 12), 523 => to_unsigned(1598, 12), 524 => to_unsigned(3696, 12), 525 => to_unsigned(2920, 12), 526 => to_unsigned(1531, 12), 527 => to_unsigned(1625, 12), 528 => to_unsigned(3489, 12), 529 => to_unsigned(361, 12), 530 => to_unsigned(346, 12), 531 => to_unsigned(3179, 12), 532 => to_unsigned(3467, 12), 533 => to_unsigned(1373, 12), 534 => to_unsigned(1335, 12), 535 => to_unsigned(202, 12), 536 => to_unsigned(277, 12), 537 => to_unsigned(344, 12), 538 => to_unsigned(3533, 12), 539 => to_unsigned(545, 12), 540 => to_unsigned(3308, 12), 541 => to_unsigned(3593, 12), 542 => to_unsigned(429, 12), 543 => to_unsigned(2723, 12), 544 => to_unsigned(1378, 12), 545 => to_unsigned(1317, 12), 546 => to_unsigned(3287, 12), 547 => to_unsigned(2154, 12), 548 => to_unsigned(1387, 12), 549 => to_unsigned(3005, 12), 550 => to_unsigned(1653, 12), 551 => to_unsigned(107, 12), 552 => to_unsigned(3778, 12), 553 => to_unsigned(1318, 12), 554 => to_unsigned(3819, 12), 555 => to_unsigned(686, 12), 556 => to_unsigned(3457, 12), 557 => to_unsigned(1258, 12), 558 => to_unsigned(349, 12), 559 => to_unsigned(1594, 12), 560 => to_unsigned(2271, 12), 561 => to_unsigned(1604, 12), 562 => to_unsigned(430, 12), 563 => to_unsigned(3673, 12), 564 => to_unsigned(2167, 12), 565 => to_unsigned(1645, 12), 566 => to_unsigned(1833, 12), 567 => to_unsigned(2424, 12), 568 => to_unsigned(3847, 12), 569 => to_unsigned(3564, 12), 570 => to_unsigned(2115, 12), 571 => to_unsigned(2170, 12), 572 => to_unsigned(2215, 12), 573 => to_unsigned(391, 12), 574 => to_unsigned(1812, 12), 575 => to_unsigned(856, 12), 576 => to_unsigned(1944, 12), 577 => to_unsigned(1313, 12), 578 => to_unsigned(3506, 12), 579 => to_unsigned(2768, 12), 580 => to_unsigned(1659, 12), 581 => to_unsigned(1865, 12), 582 => to_unsigned(1052, 12), 583 => to_unsigned(2894, 12), 584 => to_unsigned(1438, 12), 585 => to_unsigned(2477, 12), 586 => to_unsigned(3786, 12), 587 => to_unsigned(3041, 12), 588 => to_unsigned(1948, 12), 589 => to_unsigned(3007, 12), 590 => to_unsigned(573, 12), 591 => to_unsigned(966, 12), 592 => to_unsigned(2216, 12), 593 => to_unsigned(454, 12), 594 => to_unsigned(2536, 12), 595 => to_unsigned(469, 12), 596 => to_unsigned(2417, 12), 597 => to_unsigned(408, 12), 598 => to_unsigned(2097, 12), 599 => to_unsigned(951, 12), 600 => to_unsigned(2063, 12), 601 => to_unsigned(2187, 12), 602 => to_unsigned(1326, 12), 603 => to_unsigned(2584, 12), 604 => to_unsigned(594, 12), 605 => to_unsigned(2264, 12), 606 => to_unsigned(1367, 12), 607 => to_unsigned(2658, 12), 608 => to_unsigned(517, 12), 609 => to_unsigned(2382, 12), 610 => to_unsigned(4087, 12), 611 => to_unsigned(1055, 12), 612 => to_unsigned(2159, 12), 613 => to_unsigned(1977, 12), 614 => to_unsigned(3367, 12), 615 => to_unsigned(3455, 12), 616 => to_unsigned(2546, 12), 617 => to_unsigned(3960, 12), 618 => to_unsigned(3814, 12), 619 => to_unsigned(1462, 12), 620 => to_unsigned(2292, 12), 621 => to_unsigned(1617, 12), 622 => to_unsigned(3902, 12), 623 => to_unsigned(3426, 12), 624 => to_unsigned(1448, 12), 625 => to_unsigned(2432, 12), 626 => to_unsigned(2835, 12), 627 => to_unsigned(2662, 12), 628 => to_unsigned(2715, 12), 629 => to_unsigned(3676, 12), 630 => to_unsigned(1157, 12), 631 => to_unsigned(921, 12), 632 => to_unsigned(3779, 12), 633 => to_unsigned(1286, 12), 634 => to_unsigned(2580, 12), 635 => to_unsigned(1546, 12), 636 => to_unsigned(1793, 12), 637 => to_unsigned(1063, 12), 638 => to_unsigned(3449, 12), 639 => to_unsigned(3605, 12), 640 => to_unsigned(3789, 12), 641 => to_unsigned(1701, 12), 642 => to_unsigned(1291, 12), 643 => to_unsigned(3766, 12), 644 => to_unsigned(1305, 12), 645 => to_unsigned(1015, 12), 646 => to_unsigned(4086, 12), 647 => to_unsigned(1781, 12), 648 => to_unsigned(2628, 12), 649 => to_unsigned(745, 12), 650 => to_unsigned(128, 12), 651 => to_unsigned(2782, 12), 652 => to_unsigned(3316, 12), 653 => to_unsigned(3429, 12), 654 => to_unsigned(3804, 12), 655 => to_unsigned(9, 12), 656 => to_unsigned(127, 12), 657 => to_unsigned(2257, 12), 658 => to_unsigned(3774, 12), 659 => to_unsigned(1807, 12), 660 => to_unsigned(2357, 12), 661 => to_unsigned(307, 12), 662 => to_unsigned(885, 12), 663 => to_unsigned(423, 12), 664 => to_unsigned(2640, 12), 665 => to_unsigned(2283, 12), 666 => to_unsigned(2041, 12), 667 => to_unsigned(280, 12), 668 => to_unsigned(762, 12), 669 => to_unsigned(1702, 12), 670 => to_unsigned(3046, 12), 671 => to_unsigned(2731, 12), 672 => to_unsigned(3089, 12), 673 => to_unsigned(2348, 12), 674 => to_unsigned(3509, 12), 675 => to_unsigned(2580, 12), 676 => to_unsigned(1033, 12), 677 => to_unsigned(1439, 12), 678 => to_unsigned(3207, 12), 679 => to_unsigned(3162, 12), 680 => to_unsigned(55, 12), 681 => to_unsigned(3414, 12), 682 => to_unsigned(4090, 12), 683 => to_unsigned(4095, 12), 684 => to_unsigned(480, 12), 685 => to_unsigned(1796, 12), 686 => to_unsigned(530, 12), 687 => to_unsigned(2387, 12), 688 => to_unsigned(557, 12), 689 => to_unsigned(650, 12), 690 => to_unsigned(607, 12), 691 => to_unsigned(1158, 12), 692 => to_unsigned(2539, 12), 693 => to_unsigned(4092, 12), 694 => to_unsigned(115, 12), 695 => to_unsigned(361, 12), 696 => to_unsigned(2822, 12), 697 => to_unsigned(1765, 12), 698 => to_unsigned(1387, 12), 699 => to_unsigned(357, 12), 700 => to_unsigned(2479, 12), 701 => to_unsigned(3801, 12), 702 => to_unsigned(2962, 12), 703 => to_unsigned(3343, 12), 704 => to_unsigned(753, 12), 705 => to_unsigned(1244, 12), 706 => to_unsigned(1263, 12), 707 => to_unsigned(773, 12), 708 => to_unsigned(2695, 12), 709 => to_unsigned(3468, 12), 710 => to_unsigned(187, 12), 711 => to_unsigned(996, 12), 712 => to_unsigned(1712, 12), 713 => to_unsigned(1299, 12), 714 => to_unsigned(3175, 12), 715 => to_unsigned(4000, 12), 716 => to_unsigned(2357, 12), 717 => to_unsigned(1604, 12), 718 => to_unsigned(1533, 12), 719 => to_unsigned(690, 12), 720 => to_unsigned(3626, 12), 721 => to_unsigned(2365, 12), 722 => to_unsigned(2357, 12), 723 => to_unsigned(4039, 12), 724 => to_unsigned(1716, 12), 725 => to_unsigned(2690, 12), 726 => to_unsigned(746, 12), 727 => to_unsigned(3863, 12), 728 => to_unsigned(2661, 12), 729 => to_unsigned(1164, 12), 730 => to_unsigned(108, 12), 731 => to_unsigned(3360, 12), 732 => to_unsigned(1641, 12), 733 => to_unsigned(352, 12), 734 => to_unsigned(3011, 12), 735 => to_unsigned(21, 12), 736 => to_unsigned(1691, 12), 737 => to_unsigned(1370, 12), 738 => to_unsigned(1853, 12), 739 => to_unsigned(771, 12), 740 => to_unsigned(1781, 12), 741 => to_unsigned(118, 12), 742 => to_unsigned(298, 12), 743 => to_unsigned(485, 12), 744 => to_unsigned(462, 12), 745 => to_unsigned(1500, 12), 746 => to_unsigned(3541, 12), 747 => to_unsigned(821, 12), 748 => to_unsigned(2401, 12), 749 => to_unsigned(1942, 12), 750 => to_unsigned(1580, 12), 751 => to_unsigned(2964, 12), 752 => to_unsigned(2951, 12), 753 => to_unsigned(1308, 12), 754 => to_unsigned(1226, 12), 755 => to_unsigned(1738, 12), 756 => to_unsigned(3153, 12), 757 => to_unsigned(12, 12), 758 => to_unsigned(1505, 12), 759 => to_unsigned(1950, 12), 760 => to_unsigned(558, 12), 761 => to_unsigned(3029, 12), 762 => to_unsigned(1266, 12), 763 => to_unsigned(2766, 12), 764 => to_unsigned(3878, 12), 765 => to_unsigned(3068, 12), 766 => to_unsigned(2881, 12), 767 => to_unsigned(3517, 12), 768 => to_unsigned(2934, 12), 769 => to_unsigned(2499, 12), 770 => to_unsigned(1318, 12), 771 => to_unsigned(3103, 12), 772 => to_unsigned(4092, 12), 773 => to_unsigned(3931, 12), 774 => to_unsigned(1979, 12), 775 => to_unsigned(2198, 12), 776 => to_unsigned(1680, 12), 777 => to_unsigned(1140, 12), 778 => to_unsigned(245, 12), 779 => to_unsigned(2345, 12), 780 => to_unsigned(1742, 12), 781 => to_unsigned(1393, 12), 782 => to_unsigned(3425, 12), 783 => to_unsigned(2595, 12), 784 => to_unsigned(1996, 12), 785 => to_unsigned(632, 12), 786 => to_unsigned(1010, 12), 787 => to_unsigned(3232, 12), 788 => to_unsigned(2885, 12), 789 => to_unsigned(2469, 12), 790 => to_unsigned(657, 12), 791 => to_unsigned(968, 12), 792 => to_unsigned(1150, 12), 793 => to_unsigned(693, 12), 794 => to_unsigned(1107, 12), 795 => to_unsigned(1849, 12), 796 => to_unsigned(2429, 12), 797 => to_unsigned(2568, 12), 798 => to_unsigned(2701, 12), 799 => to_unsigned(3381, 12), 800 => to_unsigned(2568, 12), 801 => to_unsigned(354, 12), 802 => to_unsigned(2733, 12), 803 => to_unsigned(1477, 12), 804 => to_unsigned(401, 12), 805 => to_unsigned(2559, 12), 806 => to_unsigned(2962, 12), 807 => to_unsigned(1089, 12), 808 => to_unsigned(3334, 12), 809 => to_unsigned(2266, 12), 810 => to_unsigned(3448, 12), 811 => to_unsigned(267, 12), 812 => to_unsigned(762, 12), 813 => to_unsigned(169, 12), 814 => to_unsigned(2300, 12), 815 => to_unsigned(716, 12), 816 => to_unsigned(3042, 12), 817 => to_unsigned(2440, 12), 818 => to_unsigned(3165, 12), 819 => to_unsigned(3325, 12), 820 => to_unsigned(1114, 12), 821 => to_unsigned(2366, 12), 822 => to_unsigned(787, 12), 823 => to_unsigned(3335, 12), 824 => to_unsigned(1017, 12), 825 => to_unsigned(3260, 12), 826 => to_unsigned(1745, 12), 827 => to_unsigned(1615, 12), 828 => to_unsigned(1350, 12), 829 => to_unsigned(353, 12), 830 => to_unsigned(3362, 12), 831 => to_unsigned(552, 12), 832 => to_unsigned(2817, 12), 833 => to_unsigned(78, 12), 834 => to_unsigned(1688, 12), 835 => to_unsigned(99, 12), 836 => to_unsigned(3525, 12), 837 => to_unsigned(4059, 12), 838 => to_unsigned(3647, 12), 839 => to_unsigned(3613, 12), 840 => to_unsigned(2797, 12), 841 => to_unsigned(2368, 12), 842 => to_unsigned(3655, 12), 843 => to_unsigned(2490, 12), 844 => to_unsigned(3375, 12), 845 => to_unsigned(66, 12), 846 => to_unsigned(1578, 12), 847 => to_unsigned(84, 12), 848 => to_unsigned(2398, 12), 849 => to_unsigned(1283, 12), 850 => to_unsigned(3046, 12), 851 => to_unsigned(2127, 12), 852 => to_unsigned(2131, 12), 853 => to_unsigned(3661, 12), 854 => to_unsigned(1953, 12), 855 => to_unsigned(1768, 12), 856 => to_unsigned(3100, 12), 857 => to_unsigned(3005, 12), 858 => to_unsigned(3734, 12), 859 => to_unsigned(2500, 12), 860 => to_unsigned(2006, 12), 861 => to_unsigned(2689, 12), 862 => to_unsigned(2480, 12), 863 => to_unsigned(1262, 12), 864 => to_unsigned(3490, 12), 865 => to_unsigned(1729, 12), 866 => to_unsigned(1874, 12), 867 => to_unsigned(994, 12), 868 => to_unsigned(559, 12), 869 => to_unsigned(3573, 12), 870 => to_unsigned(1125, 12), 871 => to_unsigned(2578, 12), 872 => to_unsigned(3746, 12), 873 => to_unsigned(1397, 12), 874 => to_unsigned(819, 12), 875 => to_unsigned(2085, 12), 876 => to_unsigned(2373, 12), 877 => to_unsigned(3889, 12), 878 => to_unsigned(453, 12), 879 => to_unsigned(2244, 12), 880 => to_unsigned(1456, 12), 881 => to_unsigned(2603, 12), 882 => to_unsigned(769, 12), 883 => to_unsigned(778, 12), 884 => to_unsigned(2835, 12), 885 => to_unsigned(584, 12), 886 => to_unsigned(3866, 12), 887 => to_unsigned(1841, 12), 888 => to_unsigned(363, 12), 889 => to_unsigned(1890, 12), 890 => to_unsigned(195, 12), 891 => to_unsigned(1930, 12), 892 => to_unsigned(2423, 12), 893 => to_unsigned(898, 12), 894 => to_unsigned(1042, 12), 895 => to_unsigned(2847, 12), 896 => to_unsigned(1571, 12), 897 => to_unsigned(3548, 12), 898 => to_unsigned(1584, 12), 899 => to_unsigned(3885, 12), 900 => to_unsigned(3430, 12), 901 => to_unsigned(1029, 12), 902 => to_unsigned(1093, 12), 903 => to_unsigned(315, 12), 904 => to_unsigned(3550, 12), 905 => to_unsigned(3313, 12), 906 => to_unsigned(1318, 12), 907 => to_unsigned(1005, 12), 908 => to_unsigned(3039, 12), 909 => to_unsigned(1352, 12), 910 => to_unsigned(1968, 12), 911 => to_unsigned(1734, 12), 912 => to_unsigned(718, 12), 913 => to_unsigned(1410, 12), 914 => to_unsigned(3349, 12), 915 => to_unsigned(193, 12), 916 => to_unsigned(2195, 12), 917 => to_unsigned(1626, 12), 918 => to_unsigned(2199, 12), 919 => to_unsigned(3949, 12), 920 => to_unsigned(887, 12), 921 => to_unsigned(2375, 12), 922 => to_unsigned(3609, 12), 923 => to_unsigned(1177, 12), 924 => to_unsigned(1928, 12), 925 => to_unsigned(825, 12), 926 => to_unsigned(1228, 12), 927 => to_unsigned(2393, 12), 928 => to_unsigned(2271, 12), 929 => to_unsigned(262, 12), 930 => to_unsigned(1268, 12), 931 => to_unsigned(98, 12), 932 => to_unsigned(1959, 12), 933 => to_unsigned(3275, 12), 934 => to_unsigned(3483, 12), 935 => to_unsigned(1196, 12), 936 => to_unsigned(2416, 12), 937 => to_unsigned(1079, 12), 938 => to_unsigned(627, 12), 939 => to_unsigned(1177, 12), 940 => to_unsigned(803, 12), 941 => to_unsigned(2991, 12), 942 => to_unsigned(2290, 12), 943 => to_unsigned(3097, 12), 944 => to_unsigned(3823, 12), 945 => to_unsigned(938, 12), 946 => to_unsigned(1463, 12), 947 => to_unsigned(4021, 12), 948 => to_unsigned(2235, 12), 949 => to_unsigned(2344, 12), 950 => to_unsigned(1073, 12), 951 => to_unsigned(3149, 12), 952 => to_unsigned(1626, 12), 953 => to_unsigned(2460, 12), 954 => to_unsigned(1474, 12), 955 => to_unsigned(2628, 12), 956 => to_unsigned(2380, 12), 957 => to_unsigned(720, 12), 958 => to_unsigned(2348, 12), 959 => to_unsigned(591, 12), 960 => to_unsigned(2785, 12), 961 => to_unsigned(3171, 12), 962 => to_unsigned(2815, 12), 963 => to_unsigned(590, 12), 964 => to_unsigned(3730, 12), 965 => to_unsigned(3349, 12), 966 => to_unsigned(3233, 12), 967 => to_unsigned(412, 12), 968 => to_unsigned(2057, 12), 969 => to_unsigned(3345, 12), 970 => to_unsigned(2824, 12), 971 => to_unsigned(2670, 12), 972 => to_unsigned(2388, 12), 973 => to_unsigned(537, 12), 974 => to_unsigned(3367, 12), 975 => to_unsigned(3927, 12), 976 => to_unsigned(2821, 12), 977 => to_unsigned(3706, 12), 978 => to_unsigned(56, 12), 979 => to_unsigned(2886, 12), 980 => to_unsigned(3873, 12), 981 => to_unsigned(682, 12), 982 => to_unsigned(2786, 12), 983 => to_unsigned(1020, 12), 984 => to_unsigned(2033, 12), 985 => to_unsigned(1126, 12), 986 => to_unsigned(3356, 12), 987 => to_unsigned(1162, 12), 988 => to_unsigned(2217, 12), 989 => to_unsigned(877, 12), 990 => to_unsigned(4068, 12), 991 => to_unsigned(2652, 12), 992 => to_unsigned(3846, 12), 993 => to_unsigned(3379, 12), 994 => to_unsigned(13, 12), 995 => to_unsigned(2446, 12), 996 => to_unsigned(3141, 12), 997 => to_unsigned(4016, 12), 998 => to_unsigned(850, 12), 999 => to_unsigned(2594, 12), 1000 => to_unsigned(1324, 12), 1001 => to_unsigned(1146, 12), 1002 => to_unsigned(2330, 12), 1003 => to_unsigned(561, 12), 1004 => to_unsigned(3203, 12), 1005 => to_unsigned(1441, 12), 1006 => to_unsigned(1118, 12), 1007 => to_unsigned(2977, 12), 1008 => to_unsigned(2010, 12), 1009 => to_unsigned(434, 12), 1010 => to_unsigned(678, 12), 1011 => to_unsigned(1210, 12), 1012 => to_unsigned(2025, 12), 1013 => to_unsigned(3405, 12), 1014 => to_unsigned(2685, 12), 1015 => to_unsigned(2583, 12), 1016 => to_unsigned(3145, 12), 1017 => to_unsigned(3555, 12), 1018 => to_unsigned(1852, 12), 1019 => to_unsigned(1325, 12), 1020 => to_unsigned(685, 12), 1021 => to_unsigned(913, 12), 1022 => to_unsigned(2762, 12), 1023 => to_unsigned(2137, 12), 1024 => to_unsigned(3440, 12), 1025 => to_unsigned(582, 12), 1026 => to_unsigned(889, 12), 1027 => to_unsigned(2297, 12), 1028 => to_unsigned(1390, 12), 1029 => to_unsigned(3712, 12), 1030 => to_unsigned(2027, 12), 1031 => to_unsigned(1327, 12), 1032 => to_unsigned(737, 12), 1033 => to_unsigned(1496, 12), 1034 => to_unsigned(997, 12), 1035 => to_unsigned(3935, 12), 1036 => to_unsigned(2927, 12), 1037 => to_unsigned(2344, 12), 1038 => to_unsigned(101, 12), 1039 => to_unsigned(3632, 12), 1040 => to_unsigned(1475, 12), 1041 => to_unsigned(1776, 12), 1042 => to_unsigned(2343, 12), 1043 => to_unsigned(3140, 12), 1044 => to_unsigned(3111, 12), 1045 => to_unsigned(3846, 12), 1046 => to_unsigned(1074, 12), 1047 => to_unsigned(3172, 12), 1048 => to_unsigned(4015, 12), 1049 => to_unsigned(1881, 12), 1050 => to_unsigned(523, 12), 1051 => to_unsigned(1159, 12), 1052 => to_unsigned(3101, 12), 1053 => to_unsigned(1975, 12), 1054 => to_unsigned(1966, 12), 1055 => to_unsigned(3085, 12), 1056 => to_unsigned(2243, 12), 1057 => to_unsigned(2151, 12), 1058 => to_unsigned(2067, 12), 1059 => to_unsigned(657, 12), 1060 => to_unsigned(4008, 12), 1061 => to_unsigned(1161, 12), 1062 => to_unsigned(1736, 12), 1063 => to_unsigned(2768, 12), 1064 => to_unsigned(844, 12), 1065 => to_unsigned(4056, 12), 1066 => to_unsigned(3145, 12), 1067 => to_unsigned(2920, 12), 1068 => to_unsigned(1925, 12), 1069 => to_unsigned(3325, 12), 1070 => to_unsigned(889, 12), 1071 => to_unsigned(319, 12), 1072 => to_unsigned(2547, 12), 1073 => to_unsigned(1572, 12), 1074 => to_unsigned(46, 12), 1075 => to_unsigned(2520, 12), 1076 => to_unsigned(631, 12), 1077 => to_unsigned(659, 12), 1078 => to_unsigned(2367, 12), 1079 => to_unsigned(2131, 12), 1080 => to_unsigned(2295, 12), 1081 => to_unsigned(2489, 12), 1082 => to_unsigned(2567, 12), 1083 => to_unsigned(483, 12), 1084 => to_unsigned(3367, 12), 1085 => to_unsigned(451, 12), 1086 => to_unsigned(1616, 12), 1087 => to_unsigned(2789, 12), 1088 => to_unsigned(2442, 12), 1089 => to_unsigned(3280, 12), 1090 => to_unsigned(1498, 12), 1091 => to_unsigned(1830, 12), 1092 => to_unsigned(2891, 12), 1093 => to_unsigned(2130, 12), 1094 => to_unsigned(2787, 12), 1095 => to_unsigned(3288, 12), 1096 => to_unsigned(3249, 12), 1097 => to_unsigned(2418, 12), 1098 => to_unsigned(1620, 12), 1099 => to_unsigned(2511, 12), 1100 => to_unsigned(2313, 12), 1101 => to_unsigned(2694, 12), 1102 => to_unsigned(1922, 12), 1103 => to_unsigned(3031, 12), 1104 => to_unsigned(2621, 12), 1105 => to_unsigned(1459, 12), 1106 => to_unsigned(839, 12), 1107 => to_unsigned(1475, 12), 1108 => to_unsigned(3443, 12), 1109 => to_unsigned(1235, 12), 1110 => to_unsigned(3437, 12), 1111 => to_unsigned(2599, 12), 1112 => to_unsigned(910, 12), 1113 => to_unsigned(2181, 12), 1114 => to_unsigned(3603, 12), 1115 => to_unsigned(3438, 12), 1116 => to_unsigned(3447, 12), 1117 => to_unsigned(3816, 12), 1118 => to_unsigned(194, 12), 1119 => to_unsigned(3825, 12), 1120 => to_unsigned(1706, 12), 1121 => to_unsigned(2026, 12), 1122 => to_unsigned(1997, 12), 1123 => to_unsigned(1432, 12), 1124 => to_unsigned(544, 12), 1125 => to_unsigned(614, 12), 1126 => to_unsigned(2373, 12), 1127 => to_unsigned(811, 12), 1128 => to_unsigned(951, 12), 1129 => to_unsigned(1051, 12), 1130 => to_unsigned(618, 12), 1131 => to_unsigned(2048, 12), 1132 => to_unsigned(273, 12), 1133 => to_unsigned(122, 12), 1134 => to_unsigned(1896, 12), 1135 => to_unsigned(1382, 12), 1136 => to_unsigned(1615, 12), 1137 => to_unsigned(2458, 12), 1138 => to_unsigned(3662, 12), 1139 => to_unsigned(1432, 12), 1140 => to_unsigned(2754, 12), 1141 => to_unsigned(89, 12), 1142 => to_unsigned(1800, 12), 1143 => to_unsigned(1974, 12), 1144 => to_unsigned(1214, 12), 1145 => to_unsigned(460, 12), 1146 => to_unsigned(2651, 12), 1147 => to_unsigned(2576, 12), 1148 => to_unsigned(882, 12), 1149 => to_unsigned(2579, 12), 1150 => to_unsigned(3050, 12), 1151 => to_unsigned(2102, 12), 1152 => to_unsigned(1208, 12), 1153 => to_unsigned(1914, 12), 1154 => to_unsigned(632, 12), 1155 => to_unsigned(2928, 12), 1156 => to_unsigned(1403, 12), 1157 => to_unsigned(232, 12), 1158 => to_unsigned(1214, 12), 1159 => to_unsigned(3209, 12), 1160 => to_unsigned(3212, 12), 1161 => to_unsigned(949, 12), 1162 => to_unsigned(4046, 12), 1163 => to_unsigned(959, 12), 1164 => to_unsigned(849, 12), 1165 => to_unsigned(1264, 12), 1166 => to_unsigned(3844, 12), 1167 => to_unsigned(1431, 12), 1168 => to_unsigned(4082, 12), 1169 => to_unsigned(359, 12), 1170 => to_unsigned(3130, 12), 1171 => to_unsigned(3489, 12), 1172 => to_unsigned(3845, 12), 1173 => to_unsigned(3163, 12), 1174 => to_unsigned(3597, 12), 1175 => to_unsigned(3388, 12), 1176 => to_unsigned(4053, 12), 1177 => to_unsigned(3756, 12), 1178 => to_unsigned(547, 12), 1179 => to_unsigned(78, 12), 1180 => to_unsigned(1042, 12), 1181 => to_unsigned(1965, 12), 1182 => to_unsigned(3128, 12), 1183 => to_unsigned(2935, 12), 1184 => to_unsigned(1079, 12), 1185 => to_unsigned(1359, 12), 1186 => to_unsigned(3517, 12), 1187 => to_unsigned(3818, 12), 1188 => to_unsigned(2991, 12), 1189 => to_unsigned(2110, 12), 1190 => to_unsigned(2576, 12), 1191 => to_unsigned(2410, 12), 1192 => to_unsigned(2852, 12), 1193 => to_unsigned(3292, 12), 1194 => to_unsigned(1718, 12), 1195 => to_unsigned(3392, 12), 1196 => to_unsigned(3946, 12), 1197 => to_unsigned(3678, 12), 1198 => to_unsigned(3112, 12), 1199 => to_unsigned(2664, 12), 1200 => to_unsigned(2477, 12), 1201 => to_unsigned(1930, 12), 1202 => to_unsigned(3832, 12), 1203 => to_unsigned(3736, 12), 1204 => to_unsigned(1170, 12), 1205 => to_unsigned(3062, 12), 1206 => to_unsigned(1313, 12), 1207 => to_unsigned(1321, 12), 1208 => to_unsigned(774, 12), 1209 => to_unsigned(995, 12), 1210 => to_unsigned(2745, 12), 1211 => to_unsigned(3583, 12), 1212 => to_unsigned(749, 12), 1213 => to_unsigned(450, 12), 1214 => to_unsigned(1398, 12), 1215 => to_unsigned(1647, 12), 1216 => to_unsigned(3408, 12), 1217 => to_unsigned(1694, 12), 1218 => to_unsigned(2301, 12), 1219 => to_unsigned(3698, 12), 1220 => to_unsigned(1596, 12), 1221 => to_unsigned(2158, 12), 1222 => to_unsigned(3826, 12), 1223 => to_unsigned(1343, 12), 1224 => to_unsigned(1361, 12), 1225 => to_unsigned(1311, 12), 1226 => to_unsigned(2747, 12), 1227 => to_unsigned(2552, 12), 1228 => to_unsigned(1685, 12), 1229 => to_unsigned(2784, 12), 1230 => to_unsigned(1469, 12), 1231 => to_unsigned(1111, 12), 1232 => to_unsigned(2545, 12), 1233 => to_unsigned(3261, 12), 1234 => to_unsigned(2683, 12), 1235 => to_unsigned(2972, 12), 1236 => to_unsigned(731, 12), 1237 => to_unsigned(779, 12), 1238 => to_unsigned(3913, 12), 1239 => to_unsigned(899, 12), 1240 => to_unsigned(720, 12), 1241 => to_unsigned(2995, 12), 1242 => to_unsigned(841, 12), 1243 => to_unsigned(3987, 12), 1244 => to_unsigned(2115, 12), 1245 => to_unsigned(2848, 12), 1246 => to_unsigned(3440, 12), 1247 => to_unsigned(1097, 12), 1248 => to_unsigned(3178, 12), 1249 => to_unsigned(2792, 12), 1250 => to_unsigned(3854, 12), 1251 => to_unsigned(3129, 12), 1252 => to_unsigned(229, 12), 1253 => to_unsigned(303, 12), 1254 => to_unsigned(1851, 12), 1255 => to_unsigned(3288, 12), 1256 => to_unsigned(2708, 12), 1257 => to_unsigned(2401, 12), 1258 => to_unsigned(2900, 12), 1259 => to_unsigned(728, 12), 1260 => to_unsigned(4070, 12), 1261 => to_unsigned(2567, 12), 1262 => to_unsigned(1484, 12), 1263 => to_unsigned(1534, 12), 1264 => to_unsigned(3210, 12), 1265 => to_unsigned(456, 12), 1266 => to_unsigned(2547, 12), 1267 => to_unsigned(2561, 12), 1268 => to_unsigned(3036, 12), 1269 => to_unsigned(3826, 12), 1270 => to_unsigned(2140, 12), 1271 => to_unsigned(2086, 12), 1272 => to_unsigned(464, 12), 1273 => to_unsigned(3228, 12), 1274 => to_unsigned(2926, 12), 1275 => to_unsigned(2117, 12), 1276 => to_unsigned(1825, 12), 1277 => to_unsigned(1348, 12), 1278 => to_unsigned(1574, 12), 1279 => to_unsigned(1660, 12), 1280 => to_unsigned(2923, 12), 1281 => to_unsigned(1582, 12), 1282 => to_unsigned(3850, 12), 1283 => to_unsigned(255, 12), 1284 => to_unsigned(1439, 12), 1285 => to_unsigned(3732, 12), 1286 => to_unsigned(747, 12), 1287 => to_unsigned(2524, 12), 1288 => to_unsigned(3847, 12), 1289 => to_unsigned(796, 12), 1290 => to_unsigned(790, 12), 1291 => to_unsigned(906, 12), 1292 => to_unsigned(3205, 12), 1293 => to_unsigned(756, 12), 1294 => to_unsigned(893, 12), 1295 => to_unsigned(446, 12), 1296 => to_unsigned(3150, 12), 1297 => to_unsigned(2370, 12), 1298 => to_unsigned(1759, 12), 1299 => to_unsigned(2900, 12), 1300 => to_unsigned(1030, 12), 1301 => to_unsigned(74, 12), 1302 => to_unsigned(300, 12), 1303 => to_unsigned(114, 12), 1304 => to_unsigned(3960, 12), 1305 => to_unsigned(900, 12), 1306 => to_unsigned(835, 12), 1307 => to_unsigned(3820, 12), 1308 => to_unsigned(252, 12), 1309 => to_unsigned(3695, 12), 1310 => to_unsigned(2243, 12), 1311 => to_unsigned(3164, 12), 1312 => to_unsigned(3408, 12), 1313 => to_unsigned(3407, 12), 1314 => to_unsigned(1659, 12), 1315 => to_unsigned(3987, 12), 1316 => to_unsigned(1607, 12), 1317 => to_unsigned(1610, 12), 1318 => to_unsigned(1850, 12), 1319 => to_unsigned(451, 12), 1320 => to_unsigned(1147, 12), 1321 => to_unsigned(3108, 12), 1322 => to_unsigned(2320, 12), 1323 => to_unsigned(2938, 12), 1324 => to_unsigned(2801, 12), 1325 => to_unsigned(1996, 12), 1326 => to_unsigned(3613, 12), 1327 => to_unsigned(364, 12), 1328 => to_unsigned(1701, 12), 1329 => to_unsigned(2224, 12), 1330 => to_unsigned(2526, 12), 1331 => to_unsigned(862, 12), 1332 => to_unsigned(1386, 12), 1333 => to_unsigned(3529, 12), 1334 => to_unsigned(462, 12), 1335 => to_unsigned(3855, 12), 1336 => to_unsigned(3271, 12), 1337 => to_unsigned(870, 12), 1338 => to_unsigned(2262, 12), 1339 => to_unsigned(3498, 12), 1340 => to_unsigned(3858, 12), 1341 => to_unsigned(23, 12), 1342 => to_unsigned(208, 12), 1343 => to_unsigned(4020, 12), 1344 => to_unsigned(702, 12), 1345 => to_unsigned(3896, 12), 1346 => to_unsigned(3334, 12), 1347 => to_unsigned(1706, 12), 1348 => to_unsigned(3761, 12), 1349 => to_unsigned(3180, 12), 1350 => to_unsigned(696, 12), 1351 => to_unsigned(3773, 12), 1352 => to_unsigned(2235, 12), 1353 => to_unsigned(633, 12), 1354 => to_unsigned(1622, 12), 1355 => to_unsigned(1438, 12), 1356 => to_unsigned(1822, 12), 1357 => to_unsigned(171, 12), 1358 => to_unsigned(1766, 12), 1359 => to_unsigned(1802, 12), 1360 => to_unsigned(3697, 12), 1361 => to_unsigned(510, 12), 1362 => to_unsigned(1333, 12), 1363 => to_unsigned(3009, 12), 1364 => to_unsigned(1383, 12), 1365 => to_unsigned(1109, 12), 1366 => to_unsigned(1590, 12), 1367 => to_unsigned(2733, 12), 1368 => to_unsigned(3676, 12), 1369 => to_unsigned(455, 12), 1370 => to_unsigned(1258, 12), 1371 => to_unsigned(3925, 12), 1372 => to_unsigned(1056, 12), 1373 => to_unsigned(2126, 12), 1374 => to_unsigned(1769, 12), 1375 => to_unsigned(1752, 12), 1376 => to_unsigned(2226, 12), 1377 => to_unsigned(3082, 12), 1378 => to_unsigned(2475, 12), 1379 => to_unsigned(1032, 12), 1380 => to_unsigned(2744, 12), 1381 => to_unsigned(140, 12), 1382 => to_unsigned(2546, 12), 1383 => to_unsigned(3258, 12), 1384 => to_unsigned(1562, 12), 1385 => to_unsigned(2053, 12), 1386 => to_unsigned(3058, 12), 1387 => to_unsigned(1532, 12), 1388 => to_unsigned(3891, 12), 1389 => to_unsigned(4034, 12), 1390 => to_unsigned(1689, 12), 1391 => to_unsigned(3163, 12), 1392 => to_unsigned(548, 12), 1393 => to_unsigned(1899, 12), 1394 => to_unsigned(2675, 12), 1395 => to_unsigned(3127, 12), 1396 => to_unsigned(116, 12), 1397 => to_unsigned(1209, 12), 1398 => to_unsigned(2293, 12), 1399 => to_unsigned(3509, 12), 1400 => to_unsigned(2210, 12), 1401 => to_unsigned(749, 12), 1402 => to_unsigned(111, 12), 1403 => to_unsigned(2941, 12), 1404 => to_unsigned(2078, 12), 1405 => to_unsigned(3705, 12), 1406 => to_unsigned(3583, 12), 1407 => to_unsigned(1770, 12), 1408 => to_unsigned(1100, 12), 1409 => to_unsigned(3264, 12), 1410 => to_unsigned(4084, 12), 1411 => to_unsigned(915, 12), 1412 => to_unsigned(1602, 12), 1413 => to_unsigned(2892, 12), 1414 => to_unsigned(542, 12), 1415 => to_unsigned(3095, 12), 1416 => to_unsigned(705, 12), 1417 => to_unsigned(2886, 12), 1418 => to_unsigned(2061, 12), 1419 => to_unsigned(408, 12), 1420 => to_unsigned(785, 12), 1421 => to_unsigned(309, 12), 1422 => to_unsigned(3121, 12), 1423 => to_unsigned(3879, 12), 1424 => to_unsigned(1971, 12), 1425 => to_unsigned(2962, 12), 1426 => to_unsigned(2674, 12), 1427 => to_unsigned(1564, 12), 1428 => to_unsigned(1101, 12), 1429 => to_unsigned(987, 12), 1430 => to_unsigned(2550, 12), 1431 => to_unsigned(2220, 12), 1432 => to_unsigned(2826, 12), 1433 => to_unsigned(3427, 12), 1434 => to_unsigned(2882, 12), 1435 => to_unsigned(3391, 12), 1436 => to_unsigned(3275, 12), 1437 => to_unsigned(2776, 12), 1438 => to_unsigned(2344, 12), 1439 => to_unsigned(1266, 12), 1440 => to_unsigned(2429, 12), 1441 => to_unsigned(147, 12), 1442 => to_unsigned(375, 12), 1443 => to_unsigned(148, 12), 1444 => to_unsigned(3168, 12), 1445 => to_unsigned(2735, 12), 1446 => to_unsigned(1148, 12), 1447 => to_unsigned(2271, 12), 1448 => to_unsigned(3200, 12), 1449 => to_unsigned(1326, 12), 1450 => to_unsigned(1126, 12), 1451 => to_unsigned(4042, 12), 1452 => to_unsigned(2316, 12), 1453 => to_unsigned(3279, 12), 1454 => to_unsigned(2879, 12), 1455 => to_unsigned(1518, 12), 1456 => to_unsigned(1133, 12), 1457 => to_unsigned(3821, 12), 1458 => to_unsigned(3022, 12), 1459 => to_unsigned(3526, 12), 1460 => to_unsigned(1299, 12), 1461 => to_unsigned(1134, 12), 1462 => to_unsigned(2624, 12), 1463 => to_unsigned(1611, 12), 1464 => to_unsigned(2073, 12), 1465 => to_unsigned(783, 12), 1466 => to_unsigned(2724, 12), 1467 => to_unsigned(1744, 12), 1468 => to_unsigned(621, 12), 1469 => to_unsigned(363, 12), 1470 => to_unsigned(3034, 12), 1471 => to_unsigned(937, 12), 1472 => to_unsigned(3966, 12), 1473 => to_unsigned(2081, 12), 1474 => to_unsigned(2638, 12), 1475 => to_unsigned(3334, 12), 1476 => to_unsigned(3811, 12), 1477 => to_unsigned(2212, 12), 1478 => to_unsigned(1750, 12), 1479 => to_unsigned(3738, 12), 1480 => to_unsigned(2075, 12), 1481 => to_unsigned(3131, 12), 1482 => to_unsigned(1867, 12), 1483 => to_unsigned(2463, 12), 1484 => to_unsigned(259, 12), 1485 => to_unsigned(2275, 12), 1486 => to_unsigned(781, 12), 1487 => to_unsigned(1503, 12), 1488 => to_unsigned(1550, 12), 1489 => to_unsigned(831, 12), 1490 => to_unsigned(2166, 12), 1491 => to_unsigned(555, 12), 1492 => to_unsigned(658, 12), 1493 => to_unsigned(394, 12), 1494 => to_unsigned(2427, 12), 1495 => to_unsigned(2874, 12), 1496 => to_unsigned(3622, 12), 1497 => to_unsigned(2495, 12), 1498 => to_unsigned(2368, 12), 1499 => to_unsigned(1056, 12), 1500 => to_unsigned(993, 12), 1501 => to_unsigned(4072, 12), 1502 => to_unsigned(2997, 12), 1503 => to_unsigned(2753, 12), 1504 => to_unsigned(751, 12), 1505 => to_unsigned(1102, 12), 1506 => to_unsigned(1725, 12), 1507 => to_unsigned(3039, 12), 1508 => to_unsigned(242, 12), 1509 => to_unsigned(1859, 12), 1510 => to_unsigned(2197, 12), 1511 => to_unsigned(131, 12), 1512 => to_unsigned(3800, 12), 1513 => to_unsigned(266, 12), 1514 => to_unsigned(836, 12), 1515 => to_unsigned(1223, 12), 1516 => to_unsigned(2318, 12), 1517 => to_unsigned(4027, 12), 1518 => to_unsigned(4002, 12), 1519 => to_unsigned(1643, 12), 1520 => to_unsigned(3143, 12), 1521 => to_unsigned(1582, 12), 1522 => to_unsigned(3304, 12), 1523 => to_unsigned(2404, 12), 1524 => to_unsigned(1171, 12), 1525 => to_unsigned(2314, 12), 1526 => to_unsigned(473, 12), 1527 => to_unsigned(2789, 12), 1528 => to_unsigned(707, 12), 1529 => to_unsigned(535, 12), 1530 => to_unsigned(1873, 12), 1531 => to_unsigned(2398, 12), 1532 => to_unsigned(2326, 12), 1533 => to_unsigned(2298, 12), 1534 => to_unsigned(3182, 12), 1535 => to_unsigned(1027, 12), 1536 => to_unsigned(892, 12), 1537 => to_unsigned(1832, 12), 1538 => to_unsigned(8, 12), 1539 => to_unsigned(1770, 12), 1540 => to_unsigned(149, 12), 1541 => to_unsigned(3004, 12), 1542 => to_unsigned(1710, 12), 1543 => to_unsigned(582, 12), 1544 => to_unsigned(2382, 12), 1545 => to_unsigned(1300, 12), 1546 => to_unsigned(2278, 12), 1547 => to_unsigned(944, 12), 1548 => to_unsigned(2801, 12), 1549 => to_unsigned(2258, 12), 1550 => to_unsigned(2124, 12), 1551 => to_unsigned(445, 12), 1552 => to_unsigned(2707, 12), 1553 => to_unsigned(226, 12), 1554 => to_unsigned(1879, 12), 1555 => to_unsigned(440, 12), 1556 => to_unsigned(2278, 12), 1557 => to_unsigned(2955, 12), 1558 => to_unsigned(50, 12), 1559 => to_unsigned(2674, 12), 1560 => to_unsigned(233, 12), 1561 => to_unsigned(2863, 12), 1562 => to_unsigned(3083, 12), 1563 => to_unsigned(1006, 12), 1564 => to_unsigned(3813, 12), 1565 => to_unsigned(2352, 12), 1566 => to_unsigned(1458, 12), 1567 => to_unsigned(2897, 12), 1568 => to_unsigned(4072, 12), 1569 => to_unsigned(2219, 12), 1570 => to_unsigned(2328, 12), 1571 => to_unsigned(1293, 12), 1572 => to_unsigned(1139, 12), 1573 => to_unsigned(1848, 12), 1574 => to_unsigned(655, 12), 1575 => to_unsigned(1711, 12), 1576 => to_unsigned(147, 12), 1577 => to_unsigned(882, 12), 1578 => to_unsigned(2342, 12), 1579 => to_unsigned(2427, 12), 1580 => to_unsigned(3519, 12), 1581 => to_unsigned(1072, 12), 1582 => to_unsigned(1364, 12), 1583 => to_unsigned(2966, 12), 1584 => to_unsigned(1064, 12), 1585 => to_unsigned(3365, 12), 1586 => to_unsigned(1064, 12), 1587 => to_unsigned(3792, 12), 1588 => to_unsigned(684, 12), 1589 => to_unsigned(182, 12), 1590 => to_unsigned(3166, 12), 1591 => to_unsigned(392, 12), 1592 => to_unsigned(3447, 12), 1593 => to_unsigned(3518, 12), 1594 => to_unsigned(208, 12), 1595 => to_unsigned(3050, 12), 1596 => to_unsigned(1198, 12), 1597 => to_unsigned(1821, 12), 1598 => to_unsigned(841, 12), 1599 => to_unsigned(260, 12), 1600 => to_unsigned(1668, 12), 1601 => to_unsigned(32, 12), 1602 => to_unsigned(2311, 12), 1603 => to_unsigned(140, 12), 1604 => to_unsigned(3182, 12), 1605 => to_unsigned(2774, 12), 1606 => to_unsigned(3462, 12), 1607 => to_unsigned(20, 12), 1608 => to_unsigned(1003, 12), 1609 => to_unsigned(2973, 12), 1610 => to_unsigned(209, 12), 1611 => to_unsigned(3396, 12), 1612 => to_unsigned(2413, 12), 1613 => to_unsigned(2429, 12), 1614 => to_unsigned(2985, 12), 1615 => to_unsigned(2804, 12), 1616 => to_unsigned(3967, 12), 1617 => to_unsigned(2210, 12), 1618 => to_unsigned(2001, 12), 1619 => to_unsigned(387, 12), 1620 => to_unsigned(3390, 12), 1621 => to_unsigned(2892, 12), 1622 => to_unsigned(4015, 12), 1623 => to_unsigned(1503, 12), 1624 => to_unsigned(1928, 12), 1625 => to_unsigned(302, 12), 1626 => to_unsigned(2716, 12), 1627 => to_unsigned(3692, 12), 1628 => to_unsigned(3085, 12), 1629 => to_unsigned(500, 12), 1630 => to_unsigned(3553, 12), 1631 => to_unsigned(1372, 12), 1632 => to_unsigned(3737, 12), 1633 => to_unsigned(3021, 12), 1634 => to_unsigned(1883, 12), 1635 => to_unsigned(29, 12), 1636 => to_unsigned(7, 12), 1637 => to_unsigned(2522, 12), 1638 => to_unsigned(2, 12), 1639 => to_unsigned(1482, 12), 1640 => to_unsigned(388, 12), 1641 => to_unsigned(1981, 12), 1642 => to_unsigned(377, 12), 1643 => to_unsigned(730, 12), 1644 => to_unsigned(435, 12), 1645 => to_unsigned(706, 12), 1646 => to_unsigned(1564, 12), 1647 => to_unsigned(440, 12), 1648 => to_unsigned(1738, 12), 1649 => to_unsigned(3412, 12), 1650 => to_unsigned(3780, 12), 1651 => to_unsigned(1208, 12), 1652 => to_unsigned(2554, 12), 1653 => to_unsigned(1550, 12), 1654 => to_unsigned(4038, 12), 1655 => to_unsigned(349, 12), 1656 => to_unsigned(2135, 12), 1657 => to_unsigned(2114, 12), 1658 => to_unsigned(3254, 12), 1659 => to_unsigned(2846, 12), 1660 => to_unsigned(323, 12), 1661 => to_unsigned(3677, 12), 1662 => to_unsigned(1044, 12), 1663 => to_unsigned(182, 12), 1664 => to_unsigned(3407, 12), 1665 => to_unsigned(2970, 12), 1666 => to_unsigned(3518, 12), 1667 => to_unsigned(2042, 12), 1668 => to_unsigned(3129, 12), 1669 => to_unsigned(1272, 12), 1670 => to_unsigned(347, 12), 1671 => to_unsigned(2520, 12), 1672 => to_unsigned(3049, 12), 1673 => to_unsigned(2757, 12), 1674 => to_unsigned(3021, 12), 1675 => to_unsigned(2701, 12), 1676 => to_unsigned(193, 12), 1677 => to_unsigned(249, 12), 1678 => to_unsigned(2790, 12), 1679 => to_unsigned(2061, 12), 1680 => to_unsigned(2106, 12), 1681 => to_unsigned(2728, 12), 1682 => to_unsigned(3016, 12), 1683 => to_unsigned(484, 12), 1684 => to_unsigned(4090, 12), 1685 => to_unsigned(2171, 12), 1686 => to_unsigned(1415, 12), 1687 => to_unsigned(151, 12), 1688 => to_unsigned(1355, 12), 1689 => to_unsigned(580, 12), 1690 => to_unsigned(689, 12), 1691 => to_unsigned(2626, 12), 1692 => to_unsigned(3800, 12), 1693 => to_unsigned(1724, 12), 1694 => to_unsigned(445, 12), 1695 => to_unsigned(2527, 12), 1696 => to_unsigned(816, 12), 1697 => to_unsigned(3886, 12), 1698 => to_unsigned(3053, 12), 1699 => to_unsigned(2680, 12), 1700 => to_unsigned(2624, 12), 1701 => to_unsigned(1757, 12), 1702 => to_unsigned(617, 12), 1703 => to_unsigned(2013, 12), 1704 => to_unsigned(2891, 12), 1705 => to_unsigned(25, 12), 1706 => to_unsigned(3791, 12), 1707 => to_unsigned(471, 12), 1708 => to_unsigned(2825, 12), 1709 => to_unsigned(2243, 12), 1710 => to_unsigned(2475, 12), 1711 => to_unsigned(3399, 12), 1712 => to_unsigned(2172, 12), 1713 => to_unsigned(990, 12), 1714 => to_unsigned(2033, 12), 1715 => to_unsigned(3338, 12), 1716 => to_unsigned(3728, 12), 1717 => to_unsigned(1218, 12), 1718 => to_unsigned(218, 12), 1719 => to_unsigned(802, 12), 1720 => to_unsigned(307, 12), 1721 => to_unsigned(2100, 12), 1722 => to_unsigned(3037, 12), 1723 => to_unsigned(2877, 12), 1724 => to_unsigned(809, 12), 1725 => to_unsigned(3339, 12), 1726 => to_unsigned(2206, 12), 1727 => to_unsigned(180, 12), 1728 => to_unsigned(1716, 12), 1729 => to_unsigned(68, 12), 1730 => to_unsigned(799, 12), 1731 => to_unsigned(3071, 12), 1732 => to_unsigned(4004, 12), 1733 => to_unsigned(3478, 12), 1734 => to_unsigned(2918, 12), 1735 => to_unsigned(2741, 12), 1736 => to_unsigned(1823, 12), 1737 => to_unsigned(2840, 12), 1738 => to_unsigned(3423, 12), 1739 => to_unsigned(1192, 12), 1740 => to_unsigned(2054, 12), 1741 => to_unsigned(3963, 12), 1742 => to_unsigned(833, 12), 1743 => to_unsigned(1777, 12), 1744 => to_unsigned(2437, 12), 1745 => to_unsigned(3763, 12), 1746 => to_unsigned(433, 12), 1747 => to_unsigned(515, 12), 1748 => to_unsigned(247, 12), 1749 => to_unsigned(3609, 12), 1750 => to_unsigned(3077, 12), 1751 => to_unsigned(738, 12), 1752 => to_unsigned(382, 12), 1753 => to_unsigned(2848, 12), 1754 => to_unsigned(1774, 12), 1755 => to_unsigned(2827, 12), 1756 => to_unsigned(3916, 12), 1757 => to_unsigned(2263, 12), 1758 => to_unsigned(1989, 12), 1759 => to_unsigned(2694, 12), 1760 => to_unsigned(2895, 12), 1761 => to_unsigned(2233, 12), 1762 => to_unsigned(1339, 12), 1763 => to_unsigned(1522, 12), 1764 => to_unsigned(967, 12), 1765 => to_unsigned(1706, 12), 1766 => to_unsigned(647, 12), 1767 => to_unsigned(56, 12), 1768 => to_unsigned(3334, 12), 1769 => to_unsigned(413, 12), 1770 => to_unsigned(2222, 12), 1771 => to_unsigned(1291, 12), 1772 => to_unsigned(2659, 12), 1773 => to_unsigned(2305, 12), 1774 => to_unsigned(3116, 12), 1775 => to_unsigned(2238, 12), 1776 => to_unsigned(1298, 12), 1777 => to_unsigned(687, 12), 1778 => to_unsigned(4094, 12), 1779 => to_unsigned(998, 12), 1780 => to_unsigned(1804, 12), 1781 => to_unsigned(2914, 12), 1782 => to_unsigned(1590, 12), 1783 => to_unsigned(441, 12), 1784 => to_unsigned(2496, 12), 1785 => to_unsigned(3355, 12), 1786 => to_unsigned(2874, 12), 1787 => to_unsigned(391, 12), 1788 => to_unsigned(3754, 12), 1789 => to_unsigned(2019, 12), 1790 => to_unsigned(2000, 12), 1791 => to_unsigned(3186, 12), 1792 => to_unsigned(583, 12), 1793 => to_unsigned(2479, 12), 1794 => to_unsigned(2335, 12), 1795 => to_unsigned(3732, 12), 1796 => to_unsigned(2409, 12), 1797 => to_unsigned(2352, 12), 1798 => to_unsigned(1284, 12), 1799 => to_unsigned(514, 12), 1800 => to_unsigned(3296, 12), 1801 => to_unsigned(2923, 12), 1802 => to_unsigned(669, 12), 1803 => to_unsigned(2008, 12), 1804 => to_unsigned(3557, 12), 1805 => to_unsigned(3466, 12), 1806 => to_unsigned(1945, 12), 1807 => to_unsigned(1532, 12), 1808 => to_unsigned(2179, 12), 1809 => to_unsigned(1088, 12), 1810 => to_unsigned(4041, 12), 1811 => to_unsigned(57, 12), 1812 => to_unsigned(2628, 12), 1813 => to_unsigned(504, 12), 1814 => to_unsigned(2520, 12), 1815 => to_unsigned(2948, 12), 1816 => to_unsigned(3425, 12), 1817 => to_unsigned(1504, 12), 1818 => to_unsigned(3083, 12), 1819 => to_unsigned(2333, 12), 1820 => to_unsigned(226, 12), 1821 => to_unsigned(703, 12), 1822 => to_unsigned(3120, 12), 1823 => to_unsigned(3683, 12), 1824 => to_unsigned(2593, 12), 1825 => to_unsigned(1532, 12), 1826 => to_unsigned(3451, 12), 1827 => to_unsigned(2587, 12), 1828 => to_unsigned(1568, 12), 1829 => to_unsigned(3980, 12), 1830 => to_unsigned(524, 12), 1831 => to_unsigned(3843, 12), 1832 => to_unsigned(3043, 12), 1833 => to_unsigned(1017, 12), 1834 => to_unsigned(118, 12), 1835 => to_unsigned(1717, 12), 1836 => to_unsigned(1925, 12), 1837 => to_unsigned(3975, 12), 1838 => to_unsigned(2144, 12), 1839 => to_unsigned(1252, 12), 1840 => to_unsigned(2646, 12), 1841 => to_unsigned(978, 12), 1842 => to_unsigned(1115, 12), 1843 => to_unsigned(3231, 12), 1844 => to_unsigned(717, 12), 1845 => to_unsigned(582, 12), 1846 => to_unsigned(1946, 12), 1847 => to_unsigned(2567, 12), 1848 => to_unsigned(1245, 12), 1849 => to_unsigned(1123, 12), 1850 => to_unsigned(285, 12), 1851 => to_unsigned(2301, 12), 1852 => to_unsigned(2326, 12), 1853 => to_unsigned(1708, 12), 1854 => to_unsigned(1328, 12), 1855 => to_unsigned(1762, 12), 1856 => to_unsigned(3297, 12), 1857 => to_unsigned(1892, 12), 1858 => to_unsigned(1966, 12), 1859 => to_unsigned(1327, 12), 1860 => to_unsigned(2522, 12), 1861 => to_unsigned(631, 12), 1862 => to_unsigned(1999, 12), 1863 => to_unsigned(3635, 12), 1864 => to_unsigned(1237, 12), 1865 => to_unsigned(3720, 12), 1866 => to_unsigned(1139, 12), 1867 => to_unsigned(3112, 12), 1868 => to_unsigned(2003, 12), 1869 => to_unsigned(3234, 12), 1870 => to_unsigned(633, 12), 1871 => to_unsigned(2470, 12), 1872 => to_unsigned(283, 12), 1873 => to_unsigned(626, 12), 1874 => to_unsigned(846, 12), 1875 => to_unsigned(2597, 12), 1876 => to_unsigned(1098, 12), 1877 => to_unsigned(355, 12), 1878 => to_unsigned(1441, 12), 1879 => to_unsigned(3558, 12), 1880 => to_unsigned(1621, 12), 1881 => to_unsigned(2815, 12), 1882 => to_unsigned(2872, 12), 1883 => to_unsigned(2382, 12), 1884 => to_unsigned(1146, 12), 1885 => to_unsigned(1386, 12), 1886 => to_unsigned(2807, 12), 1887 => to_unsigned(1678, 12), 1888 => to_unsigned(1842, 12), 1889 => to_unsigned(630, 12), 1890 => to_unsigned(226, 12), 1891 => to_unsigned(2071, 12), 1892 => to_unsigned(1755, 12), 1893 => to_unsigned(2663, 12), 1894 => to_unsigned(144, 12), 1895 => to_unsigned(1855, 12), 1896 => to_unsigned(739, 12), 1897 => to_unsigned(209, 12), 1898 => to_unsigned(1117, 12), 1899 => to_unsigned(3752, 12), 1900 => to_unsigned(3845, 12), 1901 => to_unsigned(1463, 12), 1902 => to_unsigned(1693, 12), 1903 => to_unsigned(2940, 12), 1904 => to_unsigned(2273, 12), 1905 => to_unsigned(3117, 12), 1906 => to_unsigned(1551, 12), 1907 => to_unsigned(2149, 12), 1908 => to_unsigned(2806, 12), 1909 => to_unsigned(4027, 12), 1910 => to_unsigned(2837, 12), 1911 => to_unsigned(3335, 12), 1912 => to_unsigned(3306, 12), 1913 => to_unsigned(341, 12), 1914 => to_unsigned(3091, 12), 1915 => to_unsigned(1619, 12), 1916 => to_unsigned(67, 12), 1917 => to_unsigned(3441, 12), 1918 => to_unsigned(3276, 12), 1919 => to_unsigned(3151, 12), 1920 => to_unsigned(3270, 12), 1921 => to_unsigned(3590, 12), 1922 => to_unsigned(718, 12), 1923 => to_unsigned(1474, 12), 1924 => to_unsigned(1941, 12), 1925 => to_unsigned(1530, 12), 1926 => to_unsigned(195, 12), 1927 => to_unsigned(2995, 12), 1928 => to_unsigned(731, 12), 1929 => to_unsigned(606, 12), 1930 => to_unsigned(2079, 12), 1931 => to_unsigned(627, 12), 1932 => to_unsigned(2529, 12), 1933 => to_unsigned(2663, 12), 1934 => to_unsigned(2409, 12), 1935 => to_unsigned(2877, 12), 1936 => to_unsigned(3447, 12), 1937 => to_unsigned(3509, 12), 1938 => to_unsigned(3744, 12), 1939 => to_unsigned(3728, 12), 1940 => to_unsigned(4021, 12), 1941 => to_unsigned(1351, 12), 1942 => to_unsigned(1881, 12), 1943 => to_unsigned(435, 12), 1944 => to_unsigned(2930, 12), 1945 => to_unsigned(889, 12), 1946 => to_unsigned(1289, 12), 1947 => to_unsigned(1928, 12), 1948 => to_unsigned(3239, 12), 1949 => to_unsigned(3052, 12), 1950 => to_unsigned(1106, 12), 1951 => to_unsigned(522, 12), 1952 => to_unsigned(2957, 12), 1953 => to_unsigned(1695, 12), 1954 => to_unsigned(2604, 12), 1955 => to_unsigned(352, 12), 1956 => to_unsigned(607, 12), 1957 => to_unsigned(1478, 12), 1958 => to_unsigned(322, 12), 1959 => to_unsigned(2728, 12), 1960 => to_unsigned(1469, 12), 1961 => to_unsigned(1016, 12), 1962 => to_unsigned(238, 12), 1963 => to_unsigned(3803, 12), 1964 => to_unsigned(3541, 12), 1965 => to_unsigned(1780, 12), 1966 => to_unsigned(1964, 12), 1967 => to_unsigned(603, 12), 1968 => to_unsigned(2016, 12), 1969 => to_unsigned(3839, 12), 1970 => to_unsigned(552, 12), 1971 => to_unsigned(3210, 12), 1972 => to_unsigned(3252, 12), 1973 => to_unsigned(2757, 12), 1974 => to_unsigned(394, 12), 1975 => to_unsigned(90, 12), 1976 => to_unsigned(1014, 12), 1977 => to_unsigned(886, 12), 1978 => to_unsigned(917, 12), 1979 => to_unsigned(3748, 12), 1980 => to_unsigned(3762, 12), 1981 => to_unsigned(3823, 12), 1982 => to_unsigned(3348, 12), 1983 => to_unsigned(440, 12), 1984 => to_unsigned(3455, 12), 1985 => to_unsigned(2149, 12), 1986 => to_unsigned(3768, 12), 1987 => to_unsigned(1465, 12), 1988 => to_unsigned(3730, 12), 1989 => to_unsigned(1426, 12), 1990 => to_unsigned(3612, 12), 1991 => to_unsigned(898, 12), 1992 => to_unsigned(1585, 12), 1993 => to_unsigned(1327, 12), 1994 => to_unsigned(1203, 12), 1995 => to_unsigned(2531, 12), 1996 => to_unsigned(1782, 12), 1997 => to_unsigned(2768, 12), 1998 => to_unsigned(113, 12), 1999 => to_unsigned(1486, 12), 2000 => to_unsigned(1422, 12), 2001 => to_unsigned(2824, 12), 2002 => to_unsigned(958, 12), 2003 => to_unsigned(1797, 12), 2004 => to_unsigned(324, 12), 2005 => to_unsigned(1579, 12), 2006 => to_unsigned(2469, 12), 2007 => to_unsigned(2501, 12), 2008 => to_unsigned(2862, 12), 2009 => to_unsigned(2244, 12), 2010 => to_unsigned(1065, 12), 2011 => to_unsigned(1934, 12), 2012 => to_unsigned(528, 12), 2013 => to_unsigned(2264, 12), 2014 => to_unsigned(1205, 12), 2015 => to_unsigned(2842, 12), 2016 => to_unsigned(1081, 12), 2017 => to_unsigned(1801, 12), 2018 => to_unsigned(1584, 12), 2019 => to_unsigned(2132, 12), 2020 => to_unsigned(3162, 12), 2021 => to_unsigned(0, 12), 2022 => to_unsigned(205, 12), 2023 => to_unsigned(2179, 12), 2024 => to_unsigned(3394, 12), 2025 => to_unsigned(10, 12), 2026 => to_unsigned(3053, 12), 2027 => to_unsigned(2768, 12), 2028 => to_unsigned(3771, 12), 2029 => to_unsigned(1538, 12), 2030 => to_unsigned(3014, 12), 2031 => to_unsigned(3516, 12), 2032 => to_unsigned(4080, 12), 2033 => to_unsigned(316, 12), 2034 => to_unsigned(1887, 12), 2035 => to_unsigned(2204, 12), 2036 => to_unsigned(501, 12), 2037 => to_unsigned(184, 12), 2038 => to_unsigned(1876, 12), 2039 => to_unsigned(3334, 12), 2040 => to_unsigned(17, 12), 2041 => to_unsigned(1019, 12), 2042 => to_unsigned(1971, 12), 2043 => to_unsigned(788, 12), 2044 => to_unsigned(347, 12), 2045 => to_unsigned(2706, 12), 2046 => to_unsigned(1522, 12), 2047 => to_unsigned(197, 12)),
            8 => (0 => to_unsigned(3795, 12), 1 => to_unsigned(2609, 12), 2 => to_unsigned(1537, 12), 3 => to_unsigned(1167, 12), 4 => to_unsigned(336, 12), 5 => to_unsigned(1421, 12), 6 => to_unsigned(1864, 12), 7 => to_unsigned(810, 12), 8 => to_unsigned(613, 12), 9 => to_unsigned(3827, 12), 10 => to_unsigned(2308, 12), 11 => to_unsigned(3614, 12), 12 => to_unsigned(934, 12), 13 => to_unsigned(1656, 12), 14 => to_unsigned(966, 12), 15 => to_unsigned(3955, 12), 16 => to_unsigned(945, 12), 17 => to_unsigned(427, 12), 18 => to_unsigned(3929, 12), 19 => to_unsigned(1662, 12), 20 => to_unsigned(4000, 12), 21 => to_unsigned(3295, 12), 22 => to_unsigned(3370, 12), 23 => to_unsigned(3389, 12), 24 => to_unsigned(117, 12), 25 => to_unsigned(2369, 12), 26 => to_unsigned(987, 12), 27 => to_unsigned(448, 12), 28 => to_unsigned(2492, 12), 29 => to_unsigned(2816, 12), 30 => to_unsigned(1935, 12), 31 => to_unsigned(1664, 12), 32 => to_unsigned(226, 12), 33 => to_unsigned(4071, 12), 34 => to_unsigned(1306, 12), 35 => to_unsigned(225, 12), 36 => to_unsigned(753, 12), 37 => to_unsigned(3201, 12), 38 => to_unsigned(572, 12), 39 => to_unsigned(2271, 12), 40 => to_unsigned(1434, 12), 41 => to_unsigned(3709, 12), 42 => to_unsigned(2467, 12), 43 => to_unsigned(1194, 12), 44 => to_unsigned(91, 12), 45 => to_unsigned(3796, 12), 46 => to_unsigned(1980, 12), 47 => to_unsigned(2323, 12), 48 => to_unsigned(723, 12), 49 => to_unsigned(1417, 12), 50 => to_unsigned(124, 12), 51 => to_unsigned(3013, 12), 52 => to_unsigned(2863, 12), 53 => to_unsigned(3006, 12), 54 => to_unsigned(3458, 12), 55 => to_unsigned(4063, 12), 56 => to_unsigned(1931, 12), 57 => to_unsigned(2929, 12), 58 => to_unsigned(273, 12), 59 => to_unsigned(1220, 12), 60 => to_unsigned(1487, 12), 61 => to_unsigned(3001, 12), 62 => to_unsigned(1409, 12), 63 => to_unsigned(384, 12), 64 => to_unsigned(2563, 12), 65 => to_unsigned(3128, 12), 66 => to_unsigned(3394, 12), 67 => to_unsigned(198, 12), 68 => to_unsigned(1728, 12), 69 => to_unsigned(322, 12), 70 => to_unsigned(1998, 12), 71 => to_unsigned(118, 12), 72 => to_unsigned(1570, 12), 73 => to_unsigned(1004, 12), 74 => to_unsigned(2399, 12), 75 => to_unsigned(3960, 12), 76 => to_unsigned(2876, 12), 77 => to_unsigned(2175, 12), 78 => to_unsigned(30, 12), 79 => to_unsigned(1501, 12), 80 => to_unsigned(1918, 12), 81 => to_unsigned(2321, 12), 82 => to_unsigned(2372, 12), 83 => to_unsigned(3264, 12), 84 => to_unsigned(2300, 12), 85 => to_unsigned(1731, 12), 86 => to_unsigned(951, 12), 87 => to_unsigned(699, 12), 88 => to_unsigned(1125, 12), 89 => to_unsigned(2263, 12), 90 => to_unsigned(259, 12), 91 => to_unsigned(871, 12), 92 => to_unsigned(1286, 12), 93 => to_unsigned(3273, 12), 94 => to_unsigned(3344, 12), 95 => to_unsigned(1656, 12), 96 => to_unsigned(1811, 12), 97 => to_unsigned(3155, 12), 98 => to_unsigned(3860, 12), 99 => to_unsigned(3305, 12), 100 => to_unsigned(1857, 12), 101 => to_unsigned(286, 12), 102 => to_unsigned(4020, 12), 103 => to_unsigned(351, 12), 104 => to_unsigned(679, 12), 105 => to_unsigned(3995, 12), 106 => to_unsigned(2464, 12), 107 => to_unsigned(3669, 12), 108 => to_unsigned(2157, 12), 109 => to_unsigned(3620, 12), 110 => to_unsigned(1665, 12), 111 => to_unsigned(999, 12), 112 => to_unsigned(3587, 12), 113 => to_unsigned(3754, 12), 114 => to_unsigned(1556, 12), 115 => to_unsigned(107, 12), 116 => to_unsigned(1109, 12), 117 => to_unsigned(2256, 12), 118 => to_unsigned(3834, 12), 119 => to_unsigned(2954, 12), 120 => to_unsigned(2112, 12), 121 => to_unsigned(989, 12), 122 => to_unsigned(648, 12), 123 => to_unsigned(104, 12), 124 => to_unsigned(4045, 12), 125 => to_unsigned(2996, 12), 126 => to_unsigned(3332, 12), 127 => to_unsigned(3587, 12), 128 => to_unsigned(2370, 12), 129 => to_unsigned(3330, 12), 130 => to_unsigned(1285, 12), 131 => to_unsigned(2866, 12), 132 => to_unsigned(693, 12), 133 => to_unsigned(3625, 12), 134 => to_unsigned(2697, 12), 135 => to_unsigned(880, 12), 136 => to_unsigned(266, 12), 137 => to_unsigned(2499, 12), 138 => to_unsigned(3355, 12), 139 => to_unsigned(3687, 12), 140 => to_unsigned(4059, 12), 141 => to_unsigned(407, 12), 142 => to_unsigned(1697, 12), 143 => to_unsigned(3583, 12), 144 => to_unsigned(3065, 12), 145 => to_unsigned(1108, 12), 146 => to_unsigned(2567, 12), 147 => to_unsigned(1242, 12), 148 => to_unsigned(3962, 12), 149 => to_unsigned(1622, 12), 150 => to_unsigned(7, 12), 151 => to_unsigned(623, 12), 152 => to_unsigned(2274, 12), 153 => to_unsigned(2862, 12), 154 => to_unsigned(751, 12), 155 => to_unsigned(1134, 12), 156 => to_unsigned(2828, 12), 157 => to_unsigned(1811, 12), 158 => to_unsigned(2935, 12), 159 => to_unsigned(2387, 12), 160 => to_unsigned(1516, 12), 161 => to_unsigned(364, 12), 162 => to_unsigned(2070, 12), 163 => to_unsigned(3522, 12), 164 => to_unsigned(3406, 12), 165 => to_unsigned(3908, 12), 166 => to_unsigned(1230, 12), 167 => to_unsigned(1502, 12), 168 => to_unsigned(2270, 12), 169 => to_unsigned(1301, 12), 170 => to_unsigned(373, 12), 171 => to_unsigned(2042, 12), 172 => to_unsigned(3792, 12), 173 => to_unsigned(3730, 12), 174 => to_unsigned(1376, 12), 175 => to_unsigned(369, 12), 176 => to_unsigned(1617, 12), 177 => to_unsigned(970, 12), 178 => to_unsigned(1289, 12), 179 => to_unsigned(1466, 12), 180 => to_unsigned(2654, 12), 181 => to_unsigned(1284, 12), 182 => to_unsigned(3756, 12), 183 => to_unsigned(161, 12), 184 => to_unsigned(3041, 12), 185 => to_unsigned(1679, 12), 186 => to_unsigned(2302, 12), 187 => to_unsigned(2754, 12), 188 => to_unsigned(445, 12), 189 => to_unsigned(680, 12), 190 => to_unsigned(3728, 12), 191 => to_unsigned(2125, 12), 192 => to_unsigned(149, 12), 193 => to_unsigned(3965, 12), 194 => to_unsigned(2379, 12), 195 => to_unsigned(3577, 12), 196 => to_unsigned(3665, 12), 197 => to_unsigned(4082, 12), 198 => to_unsigned(2671, 12), 199 => to_unsigned(1593, 12), 200 => to_unsigned(3046, 12), 201 => to_unsigned(1573, 12), 202 => to_unsigned(714, 12), 203 => to_unsigned(361, 12), 204 => to_unsigned(770, 12), 205 => to_unsigned(2168, 12), 206 => to_unsigned(3799, 12), 207 => to_unsigned(2246, 12), 208 => to_unsigned(3604, 12), 209 => to_unsigned(3092, 12), 210 => to_unsigned(2237, 12), 211 => to_unsigned(3430, 12), 212 => to_unsigned(2949, 12), 213 => to_unsigned(1073, 12), 214 => to_unsigned(3397, 12), 215 => to_unsigned(2421, 12), 216 => to_unsigned(3920, 12), 217 => to_unsigned(3020, 12), 218 => to_unsigned(918, 12), 219 => to_unsigned(2804, 12), 220 => to_unsigned(3762, 12), 221 => to_unsigned(207, 12), 222 => to_unsigned(3367, 12), 223 => to_unsigned(964, 12), 224 => to_unsigned(2983, 12), 225 => to_unsigned(3345, 12), 226 => to_unsigned(2480, 12), 227 => to_unsigned(351, 12), 228 => to_unsigned(2074, 12), 229 => to_unsigned(1053, 12), 230 => to_unsigned(3723, 12), 231 => to_unsigned(383, 12), 232 => to_unsigned(2790, 12), 233 => to_unsigned(2369, 12), 234 => to_unsigned(3450, 12), 235 => to_unsigned(1010, 12), 236 => to_unsigned(1949, 12), 237 => to_unsigned(3886, 12), 238 => to_unsigned(3325, 12), 239 => to_unsigned(3819, 12), 240 => to_unsigned(2096, 12), 241 => to_unsigned(3191, 12), 242 => to_unsigned(2278, 12), 243 => to_unsigned(3635, 12), 244 => to_unsigned(2943, 12), 245 => to_unsigned(3, 12), 246 => to_unsigned(2897, 12), 247 => to_unsigned(1342, 12), 248 => to_unsigned(465, 12), 249 => to_unsigned(2052, 12), 250 => to_unsigned(3026, 12), 251 => to_unsigned(1105, 12), 252 => to_unsigned(2786, 12), 253 => to_unsigned(3779, 12), 254 => to_unsigned(1949, 12), 255 => to_unsigned(1585, 12), 256 => to_unsigned(3185, 12), 257 => to_unsigned(659, 12), 258 => to_unsigned(814, 12), 259 => to_unsigned(338, 12), 260 => to_unsigned(1831, 12), 261 => to_unsigned(330, 12), 262 => to_unsigned(2685, 12), 263 => to_unsigned(3293, 12), 264 => to_unsigned(1736, 12), 265 => to_unsigned(638, 12), 266 => to_unsigned(2472, 12), 267 => to_unsigned(2008, 12), 268 => to_unsigned(1122, 12), 269 => to_unsigned(1390, 12), 270 => to_unsigned(1211, 12), 271 => to_unsigned(3285, 12), 272 => to_unsigned(1774, 12), 273 => to_unsigned(1029, 12), 274 => to_unsigned(3140, 12), 275 => to_unsigned(1572, 12), 276 => to_unsigned(2684, 12), 277 => to_unsigned(551, 12), 278 => to_unsigned(2166, 12), 279 => to_unsigned(2645, 12), 280 => to_unsigned(2809, 12), 281 => to_unsigned(676, 12), 282 => to_unsigned(1198, 12), 283 => to_unsigned(3788, 12), 284 => to_unsigned(3789, 12), 285 => to_unsigned(195, 12), 286 => to_unsigned(173, 12), 287 => to_unsigned(2600, 12), 288 => to_unsigned(2979, 12), 289 => to_unsigned(617, 12), 290 => to_unsigned(487, 12), 291 => to_unsigned(696, 12), 292 => to_unsigned(4082, 12), 293 => to_unsigned(2334, 12), 294 => to_unsigned(3498, 12), 295 => to_unsigned(2897, 12), 296 => to_unsigned(3419, 12), 297 => to_unsigned(323, 12), 298 => to_unsigned(1306, 12), 299 => to_unsigned(1931, 12), 300 => to_unsigned(42, 12), 301 => to_unsigned(3787, 12), 302 => to_unsigned(3193, 12), 303 => to_unsigned(3219, 12), 304 => to_unsigned(883, 12), 305 => to_unsigned(341, 12), 306 => to_unsigned(3971, 12), 307 => to_unsigned(100, 12), 308 => to_unsigned(1076, 12), 309 => to_unsigned(1406, 12), 310 => to_unsigned(1941, 12), 311 => to_unsigned(1402, 12), 312 => to_unsigned(3817, 12), 313 => to_unsigned(3313, 12), 314 => to_unsigned(1260, 12), 315 => to_unsigned(3815, 12), 316 => to_unsigned(1498, 12), 317 => to_unsigned(3693, 12), 318 => to_unsigned(2781, 12), 319 => to_unsigned(1873, 12), 320 => to_unsigned(3597, 12), 321 => to_unsigned(190, 12), 322 => to_unsigned(3393, 12), 323 => to_unsigned(2678, 12), 324 => to_unsigned(3861, 12), 325 => to_unsigned(3659, 12), 326 => to_unsigned(1364, 12), 327 => to_unsigned(3273, 12), 328 => to_unsigned(3964, 12), 329 => to_unsigned(2827, 12), 330 => to_unsigned(2695, 12), 331 => to_unsigned(1692, 12), 332 => to_unsigned(655, 12), 333 => to_unsigned(3429, 12), 334 => to_unsigned(1883, 12), 335 => to_unsigned(149, 12), 336 => to_unsigned(1305, 12), 337 => to_unsigned(3800, 12), 338 => to_unsigned(1510, 12), 339 => to_unsigned(2249, 12), 340 => to_unsigned(73, 12), 341 => to_unsigned(1275, 12), 342 => to_unsigned(929, 12), 343 => to_unsigned(1484, 12), 344 => to_unsigned(1153, 12), 345 => to_unsigned(1884, 12), 346 => to_unsigned(2168, 12), 347 => to_unsigned(1767, 12), 348 => to_unsigned(2029, 12), 349 => to_unsigned(3364, 12), 350 => to_unsigned(2268, 12), 351 => to_unsigned(4003, 12), 352 => to_unsigned(1067, 12), 353 => to_unsigned(2243, 12), 354 => to_unsigned(1436, 12), 355 => to_unsigned(3081, 12), 356 => to_unsigned(3235, 12), 357 => to_unsigned(2566, 12), 358 => to_unsigned(3471, 12), 359 => to_unsigned(886, 12), 360 => to_unsigned(3543, 12), 361 => to_unsigned(2513, 12), 362 => to_unsigned(1766, 12), 363 => to_unsigned(985, 12), 364 => to_unsigned(1414, 12), 365 => to_unsigned(1617, 12), 366 => to_unsigned(999, 12), 367 => to_unsigned(85, 12), 368 => to_unsigned(1661, 12), 369 => to_unsigned(2251, 12), 370 => to_unsigned(409, 12), 371 => to_unsigned(2856, 12), 372 => to_unsigned(2311, 12), 373 => to_unsigned(3052, 12), 374 => to_unsigned(2075, 12), 375 => to_unsigned(3565, 12), 376 => to_unsigned(3978, 12), 377 => to_unsigned(297, 12), 378 => to_unsigned(3532, 12), 379 => to_unsigned(2879, 12), 380 => to_unsigned(1882, 12), 381 => to_unsigned(3786, 12), 382 => to_unsigned(740, 12), 383 => to_unsigned(805, 12), 384 => to_unsigned(1632, 12), 385 => to_unsigned(1029, 12), 386 => to_unsigned(3836, 12), 387 => to_unsigned(953, 12), 388 => to_unsigned(3385, 12), 389 => to_unsigned(3785, 12), 390 => to_unsigned(2394, 12), 391 => to_unsigned(1067, 12), 392 => to_unsigned(294, 12), 393 => to_unsigned(1624, 12), 394 => to_unsigned(1668, 12), 395 => to_unsigned(3658, 12), 396 => to_unsigned(3550, 12), 397 => to_unsigned(2265, 12), 398 => to_unsigned(2684, 12), 399 => to_unsigned(2357, 12), 400 => to_unsigned(2223, 12), 401 => to_unsigned(928, 12), 402 => to_unsigned(3099, 12), 403 => to_unsigned(2137, 12), 404 => to_unsigned(2075, 12), 405 => to_unsigned(3714, 12), 406 => to_unsigned(1342, 12), 407 => to_unsigned(2493, 12), 408 => to_unsigned(2446, 12), 409 => to_unsigned(3947, 12), 410 => to_unsigned(3009, 12), 411 => to_unsigned(1537, 12), 412 => to_unsigned(1800, 12), 413 => to_unsigned(3962, 12), 414 => to_unsigned(2407, 12), 415 => to_unsigned(1592, 12), 416 => to_unsigned(310, 12), 417 => to_unsigned(923, 12), 418 => to_unsigned(3132, 12), 419 => to_unsigned(825, 12), 420 => to_unsigned(3464, 12), 421 => to_unsigned(21, 12), 422 => to_unsigned(3201, 12), 423 => to_unsigned(1085, 12), 424 => to_unsigned(3588, 12), 425 => to_unsigned(273, 12), 426 => to_unsigned(1155, 12), 427 => to_unsigned(1310, 12), 428 => to_unsigned(172, 12), 429 => to_unsigned(3378, 12), 430 => to_unsigned(3159, 12), 431 => to_unsigned(2640, 12), 432 => to_unsigned(1151, 12), 433 => to_unsigned(345, 12), 434 => to_unsigned(1627, 12), 435 => to_unsigned(1039, 12), 436 => to_unsigned(2584, 12), 437 => to_unsigned(1793, 12), 438 => to_unsigned(3059, 12), 439 => to_unsigned(1716, 12), 440 => to_unsigned(2314, 12), 441 => to_unsigned(2377, 12), 442 => to_unsigned(941, 12), 443 => to_unsigned(2889, 12), 444 => to_unsigned(3713, 12), 445 => to_unsigned(3658, 12), 446 => to_unsigned(1577, 12), 447 => to_unsigned(1130, 12), 448 => to_unsigned(3613, 12), 449 => to_unsigned(3026, 12), 450 => to_unsigned(3660, 12), 451 => to_unsigned(3581, 12), 452 => to_unsigned(192, 12), 453 => to_unsigned(1467, 12), 454 => to_unsigned(2909, 12), 455 => to_unsigned(1090, 12), 456 => to_unsigned(581, 12), 457 => to_unsigned(1552, 12), 458 => to_unsigned(2062, 12), 459 => to_unsigned(2058, 12), 460 => to_unsigned(2180, 12), 461 => to_unsigned(1532, 12), 462 => to_unsigned(1470, 12), 463 => to_unsigned(1030, 12), 464 => to_unsigned(2668, 12), 465 => to_unsigned(3223, 12), 466 => to_unsigned(1109, 12), 467 => to_unsigned(2820, 12), 468 => to_unsigned(55, 12), 469 => to_unsigned(2152, 12), 470 => to_unsigned(1793, 12), 471 => to_unsigned(3535, 12), 472 => to_unsigned(2765, 12), 473 => to_unsigned(683, 12), 474 => to_unsigned(1010, 12), 475 => to_unsigned(3625, 12), 476 => to_unsigned(1456, 12), 477 => to_unsigned(1374, 12), 478 => to_unsigned(1128, 12), 479 => to_unsigned(2531, 12), 480 => to_unsigned(3661, 12), 481 => to_unsigned(1371, 12), 482 => to_unsigned(39, 12), 483 => to_unsigned(4044, 12), 484 => to_unsigned(3497, 12), 485 => to_unsigned(2822, 12), 486 => to_unsigned(3880, 12), 487 => to_unsigned(17, 12), 488 => to_unsigned(2981, 12), 489 => to_unsigned(130, 12), 490 => to_unsigned(1980, 12), 491 => to_unsigned(2425, 12), 492 => to_unsigned(106, 12), 493 => to_unsigned(1731, 12), 494 => to_unsigned(1276, 12), 495 => to_unsigned(428, 12), 496 => to_unsigned(637, 12), 497 => to_unsigned(1578, 12), 498 => to_unsigned(4044, 12), 499 => to_unsigned(1240, 12), 500 => to_unsigned(3708, 12), 501 => to_unsigned(1529, 12), 502 => to_unsigned(878, 12), 503 => to_unsigned(1869, 12), 504 => to_unsigned(515, 12), 505 => to_unsigned(4009, 12), 506 => to_unsigned(3154, 12), 507 => to_unsigned(500, 12), 508 => to_unsigned(2389, 12), 509 => to_unsigned(231, 12), 510 => to_unsigned(2661, 12), 511 => to_unsigned(1211, 12), 512 => to_unsigned(475, 12), 513 => to_unsigned(3981, 12), 514 => to_unsigned(1303, 12), 515 => to_unsigned(2420, 12), 516 => to_unsigned(2894, 12), 517 => to_unsigned(1105, 12), 518 => to_unsigned(600, 12), 519 => to_unsigned(866, 12), 520 => to_unsigned(1038, 12), 521 => to_unsigned(644, 12), 522 => to_unsigned(3192, 12), 523 => to_unsigned(2590, 12), 524 => to_unsigned(2140, 12), 525 => to_unsigned(2229, 12), 526 => to_unsigned(2786, 12), 527 => to_unsigned(849, 12), 528 => to_unsigned(289, 12), 529 => to_unsigned(1994, 12), 530 => to_unsigned(3106, 12), 531 => to_unsigned(3006, 12), 532 => to_unsigned(2745, 12), 533 => to_unsigned(661, 12), 534 => to_unsigned(593, 12), 535 => to_unsigned(4036, 12), 536 => to_unsigned(3598, 12), 537 => to_unsigned(1888, 12), 538 => to_unsigned(2020, 12), 539 => to_unsigned(3819, 12), 540 => to_unsigned(1048, 12), 541 => to_unsigned(1376, 12), 542 => to_unsigned(970, 12), 543 => to_unsigned(3006, 12), 544 => to_unsigned(1279, 12), 545 => to_unsigned(3838, 12), 546 => to_unsigned(2820, 12), 547 => to_unsigned(1390, 12), 548 => to_unsigned(2304, 12), 549 => to_unsigned(3152, 12), 550 => to_unsigned(1314, 12), 551 => to_unsigned(337, 12), 552 => to_unsigned(1123, 12), 553 => to_unsigned(3193, 12), 554 => to_unsigned(3656, 12), 555 => to_unsigned(1117, 12), 556 => to_unsigned(2957, 12), 557 => to_unsigned(3611, 12), 558 => to_unsigned(585, 12), 559 => to_unsigned(4017, 12), 560 => to_unsigned(2741, 12), 561 => to_unsigned(2213, 12), 562 => to_unsigned(2229, 12), 563 => to_unsigned(3070, 12), 564 => to_unsigned(3557, 12), 565 => to_unsigned(2100, 12), 566 => to_unsigned(661, 12), 567 => to_unsigned(1173, 12), 568 => to_unsigned(684, 12), 569 => to_unsigned(3446, 12), 570 => to_unsigned(1835, 12), 571 => to_unsigned(2723, 12), 572 => to_unsigned(3944, 12), 573 => to_unsigned(28, 12), 574 => to_unsigned(2541, 12), 575 => to_unsigned(3018, 12), 576 => to_unsigned(2136, 12), 577 => to_unsigned(3482, 12), 578 => to_unsigned(3204, 12), 579 => to_unsigned(2113, 12), 580 => to_unsigned(1305, 12), 581 => to_unsigned(2072, 12), 582 => to_unsigned(3515, 12), 583 => to_unsigned(1454, 12), 584 => to_unsigned(2724, 12), 585 => to_unsigned(3558, 12), 586 => to_unsigned(2898, 12), 587 => to_unsigned(298, 12), 588 => to_unsigned(15, 12), 589 => to_unsigned(2088, 12), 590 => to_unsigned(3943, 12), 591 => to_unsigned(0, 12), 592 => to_unsigned(1164, 12), 593 => to_unsigned(1793, 12), 594 => to_unsigned(3632, 12), 595 => to_unsigned(2236, 12), 596 => to_unsigned(1441, 12), 597 => to_unsigned(2046, 12), 598 => to_unsigned(2251, 12), 599 => to_unsigned(1149, 12), 600 => to_unsigned(2983, 12), 601 => to_unsigned(1611, 12), 602 => to_unsigned(1259, 12), 603 => to_unsigned(2754, 12), 604 => to_unsigned(411, 12), 605 => to_unsigned(724, 12), 606 => to_unsigned(384, 12), 607 => to_unsigned(1689, 12), 608 => to_unsigned(1316, 12), 609 => to_unsigned(2017, 12), 610 => to_unsigned(1280, 12), 611 => to_unsigned(226, 12), 612 => to_unsigned(1360, 12), 613 => to_unsigned(3928, 12), 614 => to_unsigned(2744, 12), 615 => to_unsigned(1559, 12), 616 => to_unsigned(1877, 12), 617 => to_unsigned(2457, 12), 618 => to_unsigned(3245, 12), 619 => to_unsigned(144, 12), 620 => to_unsigned(988, 12), 621 => to_unsigned(1083, 12), 622 => to_unsigned(915, 12), 623 => to_unsigned(2629, 12), 624 => to_unsigned(1548, 12), 625 => to_unsigned(3842, 12), 626 => to_unsigned(2731, 12), 627 => to_unsigned(3633, 12), 628 => to_unsigned(3682, 12), 629 => to_unsigned(63, 12), 630 => to_unsigned(248, 12), 631 => to_unsigned(982, 12), 632 => to_unsigned(674, 12), 633 => to_unsigned(1413, 12), 634 => to_unsigned(2335, 12), 635 => to_unsigned(2615, 12), 636 => to_unsigned(2984, 12), 637 => to_unsigned(83, 12), 638 => to_unsigned(2854, 12), 639 => to_unsigned(1528, 12), 640 => to_unsigned(3770, 12), 641 => to_unsigned(2872, 12), 642 => to_unsigned(1956, 12), 643 => to_unsigned(2623, 12), 644 => to_unsigned(87, 12), 645 => to_unsigned(3544, 12), 646 => to_unsigned(3060, 12), 647 => to_unsigned(2046, 12), 648 => to_unsigned(935, 12), 649 => to_unsigned(2633, 12), 650 => to_unsigned(1004, 12), 651 => to_unsigned(574, 12), 652 => to_unsigned(3222, 12), 653 => to_unsigned(3922, 12), 654 => to_unsigned(2863, 12), 655 => to_unsigned(3889, 12), 656 => to_unsigned(1338, 12), 657 => to_unsigned(1889, 12), 658 => to_unsigned(1143, 12), 659 => to_unsigned(1774, 12), 660 => to_unsigned(3921, 12), 661 => to_unsigned(1372, 12), 662 => to_unsigned(1085, 12), 663 => to_unsigned(1421, 12), 664 => to_unsigned(2765, 12), 665 => to_unsigned(1689, 12), 666 => to_unsigned(1058, 12), 667 => to_unsigned(3597, 12), 668 => to_unsigned(3290, 12), 669 => to_unsigned(3617, 12), 670 => to_unsigned(894, 12), 671 => to_unsigned(849, 12), 672 => to_unsigned(2744, 12), 673 => to_unsigned(3064, 12), 674 => to_unsigned(1265, 12), 675 => to_unsigned(473, 12), 676 => to_unsigned(373, 12), 677 => to_unsigned(4075, 12), 678 => to_unsigned(2229, 12), 679 => to_unsigned(3824, 12), 680 => to_unsigned(2991, 12), 681 => to_unsigned(4077, 12), 682 => to_unsigned(1588, 12), 683 => to_unsigned(2410, 12), 684 => to_unsigned(3172, 12), 685 => to_unsigned(477, 12), 686 => to_unsigned(1862, 12), 687 => to_unsigned(1512, 12), 688 => to_unsigned(1744, 12), 689 => to_unsigned(1181, 12), 690 => to_unsigned(1475, 12), 691 => to_unsigned(1678, 12), 692 => to_unsigned(403, 12), 693 => to_unsigned(2012, 12), 694 => to_unsigned(1390, 12), 695 => to_unsigned(895, 12), 696 => to_unsigned(291, 12), 697 => to_unsigned(931, 12), 698 => to_unsigned(3297, 12), 699 => to_unsigned(447, 12), 700 => to_unsigned(4093, 12), 701 => to_unsigned(2057, 12), 702 => to_unsigned(1957, 12), 703 => to_unsigned(3165, 12), 704 => to_unsigned(4083, 12), 705 => to_unsigned(2882, 12), 706 => to_unsigned(2034, 12), 707 => to_unsigned(2126, 12), 708 => to_unsigned(2183, 12), 709 => to_unsigned(1793, 12), 710 => to_unsigned(746, 12), 711 => to_unsigned(237, 12), 712 => to_unsigned(2250, 12), 713 => to_unsigned(425, 12), 714 => to_unsigned(1166, 12), 715 => to_unsigned(1922, 12), 716 => to_unsigned(1364, 12), 717 => to_unsigned(1116, 12), 718 => to_unsigned(1200, 12), 719 => to_unsigned(3813, 12), 720 => to_unsigned(1898, 12), 721 => to_unsigned(1862, 12), 722 => to_unsigned(3820, 12), 723 => to_unsigned(1996, 12), 724 => to_unsigned(1652, 12), 725 => to_unsigned(1990, 12), 726 => to_unsigned(623, 12), 727 => to_unsigned(1867, 12), 728 => to_unsigned(1302, 12), 729 => to_unsigned(1046, 12), 730 => to_unsigned(1046, 12), 731 => to_unsigned(3697, 12), 732 => to_unsigned(354, 12), 733 => to_unsigned(3727, 12), 734 => to_unsigned(1277, 12), 735 => to_unsigned(668, 12), 736 => to_unsigned(1688, 12), 737 => to_unsigned(822, 12), 738 => to_unsigned(2483, 12), 739 => to_unsigned(2891, 12), 740 => to_unsigned(429, 12), 741 => to_unsigned(2857, 12), 742 => to_unsigned(2045, 12), 743 => to_unsigned(4042, 12), 744 => to_unsigned(3847, 12), 745 => to_unsigned(1008, 12), 746 => to_unsigned(549, 12), 747 => to_unsigned(2514, 12), 748 => to_unsigned(1493, 12), 749 => to_unsigned(1372, 12), 750 => to_unsigned(1287, 12), 751 => to_unsigned(2741, 12), 752 => to_unsigned(2464, 12), 753 => to_unsigned(2429, 12), 754 => to_unsigned(1664, 12), 755 => to_unsigned(418, 12), 756 => to_unsigned(2418, 12), 757 => to_unsigned(3819, 12), 758 => to_unsigned(1381, 12), 759 => to_unsigned(1756, 12), 760 => to_unsigned(1662, 12), 761 => to_unsigned(2205, 12), 762 => to_unsigned(3014, 12), 763 => to_unsigned(1604, 12), 764 => to_unsigned(3081, 12), 765 => to_unsigned(2183, 12), 766 => to_unsigned(1362, 12), 767 => to_unsigned(3436, 12), 768 => to_unsigned(3678, 12), 769 => to_unsigned(1869, 12), 770 => to_unsigned(3693, 12), 771 => to_unsigned(1791, 12), 772 => to_unsigned(3545, 12), 773 => to_unsigned(359, 12), 774 => to_unsigned(2082, 12), 775 => to_unsigned(1135, 12), 776 => to_unsigned(3689, 12), 777 => to_unsigned(173, 12), 778 => to_unsigned(3476, 12), 779 => to_unsigned(2795, 12), 780 => to_unsigned(2776, 12), 781 => to_unsigned(143, 12), 782 => to_unsigned(2895, 12), 783 => to_unsigned(3925, 12), 784 => to_unsigned(1451, 12), 785 => to_unsigned(55, 12), 786 => to_unsigned(4038, 12), 787 => to_unsigned(1438, 12), 788 => to_unsigned(662, 12), 789 => to_unsigned(4000, 12), 790 => to_unsigned(3953, 12), 791 => to_unsigned(3218, 12), 792 => to_unsigned(1546, 12), 793 => to_unsigned(3549, 12), 794 => to_unsigned(767, 12), 795 => to_unsigned(3418, 12), 796 => to_unsigned(4043, 12), 797 => to_unsigned(538, 12), 798 => to_unsigned(3997, 12), 799 => to_unsigned(1488, 12), 800 => to_unsigned(840, 12), 801 => to_unsigned(8, 12), 802 => to_unsigned(1698, 12), 803 => to_unsigned(2908, 12), 804 => to_unsigned(678, 12), 805 => to_unsigned(127, 12), 806 => to_unsigned(360, 12), 807 => to_unsigned(2944, 12), 808 => to_unsigned(2404, 12), 809 => to_unsigned(1533, 12), 810 => to_unsigned(1562, 12), 811 => to_unsigned(2190, 12), 812 => to_unsigned(378, 12), 813 => to_unsigned(2875, 12), 814 => to_unsigned(482, 12), 815 => to_unsigned(2720, 12), 816 => to_unsigned(1075, 12), 817 => to_unsigned(2279, 12), 818 => to_unsigned(1636, 12), 819 => to_unsigned(3796, 12), 820 => to_unsigned(2745, 12), 821 => to_unsigned(2558, 12), 822 => to_unsigned(3, 12), 823 => to_unsigned(3708, 12), 824 => to_unsigned(2335, 12), 825 => to_unsigned(3726, 12), 826 => to_unsigned(3329, 12), 827 => to_unsigned(3039, 12), 828 => to_unsigned(544, 12), 829 => to_unsigned(2428, 12), 830 => to_unsigned(758, 12), 831 => to_unsigned(625, 12), 832 => to_unsigned(4065, 12), 833 => to_unsigned(139, 12), 834 => to_unsigned(970, 12), 835 => to_unsigned(3576, 12), 836 => to_unsigned(2546, 12), 837 => to_unsigned(1329, 12), 838 => to_unsigned(3468, 12), 839 => to_unsigned(834, 12), 840 => to_unsigned(2821, 12), 841 => to_unsigned(2191, 12), 842 => to_unsigned(1559, 12), 843 => to_unsigned(3453, 12), 844 => to_unsigned(306, 12), 845 => to_unsigned(3996, 12), 846 => to_unsigned(270, 12), 847 => to_unsigned(1258, 12), 848 => to_unsigned(2485, 12), 849 => to_unsigned(2367, 12), 850 => to_unsigned(660, 12), 851 => to_unsigned(104, 12), 852 => to_unsigned(254, 12), 853 => to_unsigned(2437, 12), 854 => to_unsigned(51, 12), 855 => to_unsigned(532, 12), 856 => to_unsigned(2532, 12), 857 => to_unsigned(3294, 12), 858 => to_unsigned(3900, 12), 859 => to_unsigned(2099, 12), 860 => to_unsigned(2881, 12), 861 => to_unsigned(421, 12), 862 => to_unsigned(726, 12), 863 => to_unsigned(2232, 12), 864 => to_unsigned(2966, 12), 865 => to_unsigned(293, 12), 866 => to_unsigned(1999, 12), 867 => to_unsigned(2324, 12), 868 => to_unsigned(1786, 12), 869 => to_unsigned(2999, 12), 870 => to_unsigned(1328, 12), 871 => to_unsigned(2991, 12), 872 => to_unsigned(1772, 12), 873 => to_unsigned(1321, 12), 874 => to_unsigned(3146, 12), 875 => to_unsigned(228, 12), 876 => to_unsigned(2787, 12), 877 => to_unsigned(170, 12), 878 => to_unsigned(14, 12), 879 => to_unsigned(2334, 12), 880 => to_unsigned(175, 12), 881 => to_unsigned(2011, 12), 882 => to_unsigned(2240, 12), 883 => to_unsigned(2914, 12), 884 => to_unsigned(1029, 12), 885 => to_unsigned(1850, 12), 886 => to_unsigned(691, 12), 887 => to_unsigned(1742, 12), 888 => to_unsigned(1760, 12), 889 => to_unsigned(256, 12), 890 => to_unsigned(67, 12), 891 => to_unsigned(3148, 12), 892 => to_unsigned(3673, 12), 893 => to_unsigned(2207, 12), 894 => to_unsigned(259, 12), 895 => to_unsigned(1771, 12), 896 => to_unsigned(327, 12), 897 => to_unsigned(2908, 12), 898 => to_unsigned(1007, 12), 899 => to_unsigned(2484, 12), 900 => to_unsigned(2189, 12), 901 => to_unsigned(2735, 12), 902 => to_unsigned(1037, 12), 903 => to_unsigned(954, 12), 904 => to_unsigned(1470, 12), 905 => to_unsigned(3559, 12), 906 => to_unsigned(3214, 12), 907 => to_unsigned(3802, 12), 908 => to_unsigned(936, 12), 909 => to_unsigned(3260, 12), 910 => to_unsigned(150, 12), 911 => to_unsigned(1518, 12), 912 => to_unsigned(960, 12), 913 => to_unsigned(2158, 12), 914 => to_unsigned(2203, 12), 915 => to_unsigned(3824, 12), 916 => to_unsigned(899, 12), 917 => to_unsigned(2011, 12), 918 => to_unsigned(3903, 12), 919 => to_unsigned(2588, 12), 920 => to_unsigned(1040, 12), 921 => to_unsigned(1436, 12), 922 => to_unsigned(2101, 12), 923 => to_unsigned(3699, 12), 924 => to_unsigned(1685, 12), 925 => to_unsigned(602, 12), 926 => to_unsigned(3177, 12), 927 => to_unsigned(953, 12), 928 => to_unsigned(3524, 12), 929 => to_unsigned(3243, 12), 930 => to_unsigned(2239, 12), 931 => to_unsigned(1868, 12), 932 => to_unsigned(2484, 12), 933 => to_unsigned(3134, 12), 934 => to_unsigned(983, 12), 935 => to_unsigned(85, 12), 936 => to_unsigned(162, 12), 937 => to_unsigned(2694, 12), 938 => to_unsigned(2388, 12), 939 => to_unsigned(438, 12), 940 => to_unsigned(568, 12), 941 => to_unsigned(1829, 12), 942 => to_unsigned(2319, 12), 943 => to_unsigned(3454, 12), 944 => to_unsigned(1806, 12), 945 => to_unsigned(3005, 12), 946 => to_unsigned(354, 12), 947 => to_unsigned(2329, 12), 948 => to_unsigned(908, 12), 949 => to_unsigned(3524, 12), 950 => to_unsigned(2153, 12), 951 => to_unsigned(1466, 12), 952 => to_unsigned(2701, 12), 953 => to_unsigned(2746, 12), 954 => to_unsigned(683, 12), 955 => to_unsigned(2720, 12), 956 => to_unsigned(82, 12), 957 => to_unsigned(3406, 12), 958 => to_unsigned(2854, 12), 959 => to_unsigned(893, 12), 960 => to_unsigned(1854, 12), 961 => to_unsigned(2532, 12), 962 => to_unsigned(680, 12), 963 => to_unsigned(3034, 12), 964 => to_unsigned(734, 12), 965 => to_unsigned(2855, 12), 966 => to_unsigned(955, 12), 967 => to_unsigned(3072, 12), 968 => to_unsigned(161, 12), 969 => to_unsigned(180, 12), 970 => to_unsigned(1752, 12), 971 => to_unsigned(3792, 12), 972 => to_unsigned(264, 12), 973 => to_unsigned(2144, 12), 974 => to_unsigned(3777, 12), 975 => to_unsigned(2320, 12), 976 => to_unsigned(2455, 12), 977 => to_unsigned(3933, 12), 978 => to_unsigned(263, 12), 979 => to_unsigned(2653, 12), 980 => to_unsigned(3237, 12), 981 => to_unsigned(1665, 12), 982 => to_unsigned(688, 12), 983 => to_unsigned(3384, 12), 984 => to_unsigned(3753, 12), 985 => to_unsigned(3694, 12), 986 => to_unsigned(3943, 12), 987 => to_unsigned(3088, 12), 988 => to_unsigned(2858, 12), 989 => to_unsigned(1721, 12), 990 => to_unsigned(637, 12), 991 => to_unsigned(3748, 12), 992 => to_unsigned(794, 12), 993 => to_unsigned(288, 12), 994 => to_unsigned(4080, 12), 995 => to_unsigned(1044, 12), 996 => to_unsigned(3754, 12), 997 => to_unsigned(701, 12), 998 => to_unsigned(2185, 12), 999 => to_unsigned(1810, 12), 1000 => to_unsigned(4004, 12), 1001 => to_unsigned(2897, 12), 1002 => to_unsigned(3190, 12), 1003 => to_unsigned(1913, 12), 1004 => to_unsigned(1043, 12), 1005 => to_unsigned(3528, 12), 1006 => to_unsigned(3262, 12), 1007 => to_unsigned(281, 12), 1008 => to_unsigned(2457, 12), 1009 => to_unsigned(1675, 12), 1010 => to_unsigned(2851, 12), 1011 => to_unsigned(945, 12), 1012 => to_unsigned(868, 12), 1013 => to_unsigned(2005, 12), 1014 => to_unsigned(381, 12), 1015 => to_unsigned(1423, 12), 1016 => to_unsigned(1203, 12), 1017 => to_unsigned(2010, 12), 1018 => to_unsigned(284, 12), 1019 => to_unsigned(2786, 12), 1020 => to_unsigned(3986, 12), 1021 => to_unsigned(1630, 12), 1022 => to_unsigned(1116, 12), 1023 => to_unsigned(3049, 12), 1024 => to_unsigned(2456, 12), 1025 => to_unsigned(837, 12), 1026 => to_unsigned(1111, 12), 1027 => to_unsigned(2394, 12), 1028 => to_unsigned(276, 12), 1029 => to_unsigned(3015, 12), 1030 => to_unsigned(2626, 12), 1031 => to_unsigned(2064, 12), 1032 => to_unsigned(3827, 12), 1033 => to_unsigned(347, 12), 1034 => to_unsigned(2613, 12), 1035 => to_unsigned(413, 12), 1036 => to_unsigned(199, 12), 1037 => to_unsigned(1763, 12), 1038 => to_unsigned(2213, 12), 1039 => to_unsigned(2086, 12), 1040 => to_unsigned(2698, 12), 1041 => to_unsigned(546, 12), 1042 => to_unsigned(3412, 12), 1043 => to_unsigned(2830, 12), 1044 => to_unsigned(3614, 12), 1045 => to_unsigned(2102, 12), 1046 => to_unsigned(601, 12), 1047 => to_unsigned(3238, 12), 1048 => to_unsigned(3808, 12), 1049 => to_unsigned(3515, 12), 1050 => to_unsigned(865, 12), 1051 => to_unsigned(440, 12), 1052 => to_unsigned(275, 12), 1053 => to_unsigned(3923, 12), 1054 => to_unsigned(3485, 12), 1055 => to_unsigned(3301, 12), 1056 => to_unsigned(3966, 12), 1057 => to_unsigned(897, 12), 1058 => to_unsigned(1278, 12), 1059 => to_unsigned(3637, 12), 1060 => to_unsigned(1224, 12), 1061 => to_unsigned(3716, 12), 1062 => to_unsigned(3237, 12), 1063 => to_unsigned(2483, 12), 1064 => to_unsigned(2918, 12), 1065 => to_unsigned(1625, 12), 1066 => to_unsigned(473, 12), 1067 => to_unsigned(1782, 12), 1068 => to_unsigned(3109, 12), 1069 => to_unsigned(3388, 12), 1070 => to_unsigned(3814, 12), 1071 => to_unsigned(3700, 12), 1072 => to_unsigned(279, 12), 1073 => to_unsigned(2681, 12), 1074 => to_unsigned(4094, 12), 1075 => to_unsigned(3441, 12), 1076 => to_unsigned(439, 12), 1077 => to_unsigned(3405, 12), 1078 => to_unsigned(3442, 12), 1079 => to_unsigned(2208, 12), 1080 => to_unsigned(3604, 12), 1081 => to_unsigned(1916, 12), 1082 => to_unsigned(2332, 12), 1083 => to_unsigned(2673, 12), 1084 => to_unsigned(2469, 12), 1085 => to_unsigned(3014, 12), 1086 => to_unsigned(2803, 12), 1087 => to_unsigned(576, 12), 1088 => to_unsigned(1509, 12), 1089 => to_unsigned(3921, 12), 1090 => to_unsigned(2558, 12), 1091 => to_unsigned(2640, 12), 1092 => to_unsigned(3797, 12), 1093 => to_unsigned(2377, 12), 1094 => to_unsigned(2164, 12), 1095 => to_unsigned(3691, 12), 1096 => to_unsigned(1346, 12), 1097 => to_unsigned(2689, 12), 1098 => to_unsigned(2177, 12), 1099 => to_unsigned(871, 12), 1100 => to_unsigned(726, 12), 1101 => to_unsigned(2452, 12), 1102 => to_unsigned(3198, 12), 1103 => to_unsigned(1354, 12), 1104 => to_unsigned(1004, 12), 1105 => to_unsigned(1929, 12), 1106 => to_unsigned(3716, 12), 1107 => to_unsigned(2605, 12), 1108 => to_unsigned(311, 12), 1109 => to_unsigned(2647, 12), 1110 => to_unsigned(63, 12), 1111 => to_unsigned(624, 12), 1112 => to_unsigned(328, 12), 1113 => to_unsigned(887, 12), 1114 => to_unsigned(2960, 12), 1115 => to_unsigned(2338, 12), 1116 => to_unsigned(813, 12), 1117 => to_unsigned(2974, 12), 1118 => to_unsigned(3976, 12), 1119 => to_unsigned(163, 12), 1120 => to_unsigned(1210, 12), 1121 => to_unsigned(700, 12), 1122 => to_unsigned(4060, 12), 1123 => to_unsigned(182, 12), 1124 => to_unsigned(1559, 12), 1125 => to_unsigned(901, 12), 1126 => to_unsigned(3939, 12), 1127 => to_unsigned(632, 12), 1128 => to_unsigned(3164, 12), 1129 => to_unsigned(972, 12), 1130 => to_unsigned(2596, 12), 1131 => to_unsigned(90, 12), 1132 => to_unsigned(660, 12), 1133 => to_unsigned(1507, 12), 1134 => to_unsigned(3287, 12), 1135 => to_unsigned(1277, 12), 1136 => to_unsigned(1858, 12), 1137 => to_unsigned(3786, 12), 1138 => to_unsigned(1924, 12), 1139 => to_unsigned(125, 12), 1140 => to_unsigned(2289, 12), 1141 => to_unsigned(3555, 12), 1142 => to_unsigned(2339, 12), 1143 => to_unsigned(563, 12), 1144 => to_unsigned(274, 12), 1145 => to_unsigned(3346, 12), 1146 => to_unsigned(3866, 12), 1147 => to_unsigned(2303, 12), 1148 => to_unsigned(2618, 12), 1149 => to_unsigned(3562, 12), 1150 => to_unsigned(2849, 12), 1151 => to_unsigned(2215, 12), 1152 => to_unsigned(851, 12), 1153 => to_unsigned(2899, 12), 1154 => to_unsigned(1540, 12), 1155 => to_unsigned(2958, 12), 1156 => to_unsigned(1227, 12), 1157 => to_unsigned(1637, 12), 1158 => to_unsigned(1109, 12), 1159 => to_unsigned(3077, 12), 1160 => to_unsigned(4073, 12), 1161 => to_unsigned(1678, 12), 1162 => to_unsigned(4038, 12), 1163 => to_unsigned(2126, 12), 1164 => to_unsigned(1414, 12), 1165 => to_unsigned(586, 12), 1166 => to_unsigned(3217, 12), 1167 => to_unsigned(109, 12), 1168 => to_unsigned(3287, 12), 1169 => to_unsigned(2242, 12), 1170 => to_unsigned(726, 12), 1171 => to_unsigned(2876, 12), 1172 => to_unsigned(3218, 12), 1173 => to_unsigned(208, 12), 1174 => to_unsigned(1143, 12), 1175 => to_unsigned(1072, 12), 1176 => to_unsigned(2370, 12), 1177 => to_unsigned(840, 12), 1178 => to_unsigned(213, 12), 1179 => to_unsigned(2659, 12), 1180 => to_unsigned(2955, 12), 1181 => to_unsigned(2857, 12), 1182 => to_unsigned(1615, 12), 1183 => to_unsigned(3251, 12), 1184 => to_unsigned(1940, 12), 1185 => to_unsigned(1140, 12), 1186 => to_unsigned(3158, 12), 1187 => to_unsigned(2021, 12), 1188 => to_unsigned(345, 12), 1189 => to_unsigned(1863, 12), 1190 => to_unsigned(728, 12), 1191 => to_unsigned(3948, 12), 1192 => to_unsigned(299, 12), 1193 => to_unsigned(1551, 12), 1194 => to_unsigned(1263, 12), 1195 => to_unsigned(1355, 12), 1196 => to_unsigned(3607, 12), 1197 => to_unsigned(2730, 12), 1198 => to_unsigned(2137, 12), 1199 => to_unsigned(1120, 12), 1200 => to_unsigned(885, 12), 1201 => to_unsigned(3031, 12), 1202 => to_unsigned(2279, 12), 1203 => to_unsigned(1518, 12), 1204 => to_unsigned(1170, 12), 1205 => to_unsigned(3565, 12), 1206 => to_unsigned(429, 12), 1207 => to_unsigned(3491, 12), 1208 => to_unsigned(929, 12), 1209 => to_unsigned(2353, 12), 1210 => to_unsigned(2860, 12), 1211 => to_unsigned(3275, 12), 1212 => to_unsigned(3517, 12), 1213 => to_unsigned(2603, 12), 1214 => to_unsigned(2338, 12), 1215 => to_unsigned(539, 12), 1216 => to_unsigned(1934, 12), 1217 => to_unsigned(899, 12), 1218 => to_unsigned(840, 12), 1219 => to_unsigned(961, 12), 1220 => to_unsigned(2312, 12), 1221 => to_unsigned(847, 12), 1222 => to_unsigned(3149, 12), 1223 => to_unsigned(3638, 12), 1224 => to_unsigned(3067, 12), 1225 => to_unsigned(1325, 12), 1226 => to_unsigned(4034, 12), 1227 => to_unsigned(3124, 12), 1228 => to_unsigned(4040, 12), 1229 => to_unsigned(3709, 12), 1230 => to_unsigned(3063, 12), 1231 => to_unsigned(2792, 12), 1232 => to_unsigned(2746, 12), 1233 => to_unsigned(3283, 12), 1234 => to_unsigned(396, 12), 1235 => to_unsigned(2680, 12), 1236 => to_unsigned(2450, 12), 1237 => to_unsigned(254, 12), 1238 => to_unsigned(2352, 12), 1239 => to_unsigned(3931, 12), 1240 => to_unsigned(3547, 12), 1241 => to_unsigned(3093, 12), 1242 => to_unsigned(144, 12), 1243 => to_unsigned(1702, 12), 1244 => to_unsigned(1220, 12), 1245 => to_unsigned(2911, 12), 1246 => to_unsigned(3863, 12), 1247 => to_unsigned(1709, 12), 1248 => to_unsigned(1251, 12), 1249 => to_unsigned(911, 12), 1250 => to_unsigned(2577, 12), 1251 => to_unsigned(108, 12), 1252 => to_unsigned(2507, 12), 1253 => to_unsigned(1916, 12), 1254 => to_unsigned(1825, 12), 1255 => to_unsigned(1429, 12), 1256 => to_unsigned(2072, 12), 1257 => to_unsigned(334, 12), 1258 => to_unsigned(3537, 12), 1259 => to_unsigned(228, 12), 1260 => to_unsigned(2717, 12), 1261 => to_unsigned(2975, 12), 1262 => to_unsigned(2541, 12), 1263 => to_unsigned(1642, 12), 1264 => to_unsigned(965, 12), 1265 => to_unsigned(485, 12), 1266 => to_unsigned(2946, 12), 1267 => to_unsigned(3892, 12), 1268 => to_unsigned(3357, 12), 1269 => to_unsigned(3702, 12), 1270 => to_unsigned(799, 12), 1271 => to_unsigned(2530, 12), 1272 => to_unsigned(2115, 12), 1273 => to_unsigned(2678, 12), 1274 => to_unsigned(1676, 12), 1275 => to_unsigned(2275, 12), 1276 => to_unsigned(660, 12), 1277 => to_unsigned(3622, 12), 1278 => to_unsigned(2865, 12), 1279 => to_unsigned(374, 12), 1280 => to_unsigned(812, 12), 1281 => to_unsigned(796, 12), 1282 => to_unsigned(1672, 12), 1283 => to_unsigned(210, 12), 1284 => to_unsigned(3210, 12), 1285 => to_unsigned(81, 12), 1286 => to_unsigned(2977, 12), 1287 => to_unsigned(3817, 12), 1288 => to_unsigned(2392, 12), 1289 => to_unsigned(3129, 12), 1290 => to_unsigned(566, 12), 1291 => to_unsigned(2188, 12), 1292 => to_unsigned(205, 12), 1293 => to_unsigned(2050, 12), 1294 => to_unsigned(91, 12), 1295 => to_unsigned(3100, 12), 1296 => to_unsigned(2836, 12), 1297 => to_unsigned(3264, 12), 1298 => to_unsigned(3624, 12), 1299 => to_unsigned(2792, 12), 1300 => to_unsigned(3306, 12), 1301 => to_unsigned(1045, 12), 1302 => to_unsigned(373, 12), 1303 => to_unsigned(3607, 12), 1304 => to_unsigned(1105, 12), 1305 => to_unsigned(3741, 12), 1306 => to_unsigned(738, 12), 1307 => to_unsigned(3450, 12), 1308 => to_unsigned(1514, 12), 1309 => to_unsigned(1450, 12), 1310 => to_unsigned(2203, 12), 1311 => to_unsigned(1702, 12), 1312 => to_unsigned(3318, 12), 1313 => to_unsigned(2935, 12), 1314 => to_unsigned(3593, 12), 1315 => to_unsigned(2874, 12), 1316 => to_unsigned(3837, 12), 1317 => to_unsigned(1522, 12), 1318 => to_unsigned(2338, 12), 1319 => to_unsigned(2810, 12), 1320 => to_unsigned(1079, 12), 1321 => to_unsigned(933, 12), 1322 => to_unsigned(687, 12), 1323 => to_unsigned(2777, 12), 1324 => to_unsigned(1685, 12), 1325 => to_unsigned(4078, 12), 1326 => to_unsigned(1965, 12), 1327 => to_unsigned(2079, 12), 1328 => to_unsigned(3595, 12), 1329 => to_unsigned(3725, 12), 1330 => to_unsigned(692, 12), 1331 => to_unsigned(1551, 12), 1332 => to_unsigned(3092, 12), 1333 => to_unsigned(3977, 12), 1334 => to_unsigned(3944, 12), 1335 => to_unsigned(3216, 12), 1336 => to_unsigned(1574, 12), 1337 => to_unsigned(1960, 12), 1338 => to_unsigned(46, 12), 1339 => to_unsigned(507, 12), 1340 => to_unsigned(83, 12), 1341 => to_unsigned(2424, 12), 1342 => to_unsigned(1936, 12), 1343 => to_unsigned(1093, 12), 1344 => to_unsigned(3858, 12), 1345 => to_unsigned(1114, 12), 1346 => to_unsigned(2279, 12), 1347 => to_unsigned(3680, 12), 1348 => to_unsigned(3627, 12), 1349 => to_unsigned(4075, 12), 1350 => to_unsigned(3752, 12), 1351 => to_unsigned(569, 12), 1352 => to_unsigned(3658, 12), 1353 => to_unsigned(1759, 12), 1354 => to_unsigned(3910, 12), 1355 => to_unsigned(2342, 12), 1356 => to_unsigned(2713, 12), 1357 => to_unsigned(1659, 12), 1358 => to_unsigned(3145, 12), 1359 => to_unsigned(1852, 12), 1360 => to_unsigned(3172, 12), 1361 => to_unsigned(1095, 12), 1362 => to_unsigned(3731, 12), 1363 => to_unsigned(1797, 12), 1364 => to_unsigned(3846, 12), 1365 => to_unsigned(2203, 12), 1366 => to_unsigned(3481, 12), 1367 => to_unsigned(752, 12), 1368 => to_unsigned(2387, 12), 1369 => to_unsigned(2215, 12), 1370 => to_unsigned(1530, 12), 1371 => to_unsigned(3989, 12), 1372 => to_unsigned(2808, 12), 1373 => to_unsigned(1510, 12), 1374 => to_unsigned(1356, 12), 1375 => to_unsigned(408, 12), 1376 => to_unsigned(3295, 12), 1377 => to_unsigned(2289, 12), 1378 => to_unsigned(91, 12), 1379 => to_unsigned(1146, 12), 1380 => to_unsigned(3134, 12), 1381 => to_unsigned(3633, 12), 1382 => to_unsigned(819, 12), 1383 => to_unsigned(3149, 12), 1384 => to_unsigned(781, 12), 1385 => to_unsigned(3648, 12), 1386 => to_unsigned(1868, 12), 1387 => to_unsigned(1683, 12), 1388 => to_unsigned(2743, 12), 1389 => to_unsigned(1099, 12), 1390 => to_unsigned(1340, 12), 1391 => to_unsigned(1225, 12), 1392 => to_unsigned(3163, 12), 1393 => to_unsigned(1000, 12), 1394 => to_unsigned(3570, 12), 1395 => to_unsigned(4007, 12), 1396 => to_unsigned(55, 12), 1397 => to_unsigned(867, 12), 1398 => to_unsigned(2471, 12), 1399 => to_unsigned(1850, 12), 1400 => to_unsigned(943, 12), 1401 => to_unsigned(4087, 12), 1402 => to_unsigned(2220, 12), 1403 => to_unsigned(635, 12), 1404 => to_unsigned(1039, 12), 1405 => to_unsigned(87, 12), 1406 => to_unsigned(1887, 12), 1407 => to_unsigned(3755, 12), 1408 => to_unsigned(2514, 12), 1409 => to_unsigned(566, 12), 1410 => to_unsigned(268, 12), 1411 => to_unsigned(240, 12), 1412 => to_unsigned(3839, 12), 1413 => to_unsigned(2051, 12), 1414 => to_unsigned(3944, 12), 1415 => to_unsigned(1617, 12), 1416 => to_unsigned(3851, 12), 1417 => to_unsigned(3430, 12), 1418 => to_unsigned(3583, 12), 1419 => to_unsigned(866, 12), 1420 => to_unsigned(2364, 12), 1421 => to_unsigned(2336, 12), 1422 => to_unsigned(2433, 12), 1423 => to_unsigned(2111, 12), 1424 => to_unsigned(3883, 12), 1425 => to_unsigned(1047, 12), 1426 => to_unsigned(513, 12), 1427 => to_unsigned(2878, 12), 1428 => to_unsigned(248, 12), 1429 => to_unsigned(3639, 12), 1430 => to_unsigned(2354, 12), 1431 => to_unsigned(418, 12), 1432 => to_unsigned(35, 12), 1433 => to_unsigned(2880, 12), 1434 => to_unsigned(2843, 12), 1435 => to_unsigned(1244, 12), 1436 => to_unsigned(3726, 12), 1437 => to_unsigned(2142, 12), 1438 => to_unsigned(1673, 12), 1439 => to_unsigned(907, 12), 1440 => to_unsigned(985, 12), 1441 => to_unsigned(87, 12), 1442 => to_unsigned(1908, 12), 1443 => to_unsigned(3419, 12), 1444 => to_unsigned(2334, 12), 1445 => to_unsigned(2687, 12), 1446 => to_unsigned(607, 12), 1447 => to_unsigned(2893, 12), 1448 => to_unsigned(4040, 12), 1449 => to_unsigned(1682, 12), 1450 => to_unsigned(1680, 12), 1451 => to_unsigned(3140, 12), 1452 => to_unsigned(398, 12), 1453 => to_unsigned(3063, 12), 1454 => to_unsigned(2699, 12), 1455 => to_unsigned(4055, 12), 1456 => to_unsigned(257, 12), 1457 => to_unsigned(3052, 12), 1458 => to_unsigned(3643, 12), 1459 => to_unsigned(2514, 12), 1460 => to_unsigned(1863, 12), 1461 => to_unsigned(922, 12), 1462 => to_unsigned(1397, 12), 1463 => to_unsigned(3788, 12), 1464 => to_unsigned(1833, 12), 1465 => to_unsigned(3369, 12), 1466 => to_unsigned(688, 12), 1467 => to_unsigned(2258, 12), 1468 => to_unsigned(580, 12), 1469 => to_unsigned(835, 12), 1470 => to_unsigned(1897, 12), 1471 => to_unsigned(2434, 12), 1472 => to_unsigned(534, 12), 1473 => to_unsigned(2557, 12), 1474 => to_unsigned(2058, 12), 1475 => to_unsigned(1708, 12), 1476 => to_unsigned(2152, 12), 1477 => to_unsigned(2182, 12), 1478 => to_unsigned(3189, 12), 1479 => to_unsigned(101, 12), 1480 => to_unsigned(2725, 12), 1481 => to_unsigned(2703, 12), 1482 => to_unsigned(849, 12), 1483 => to_unsigned(3174, 12), 1484 => to_unsigned(2023, 12), 1485 => to_unsigned(1601, 12), 1486 => to_unsigned(3047, 12), 1487 => to_unsigned(3333, 12), 1488 => to_unsigned(2374, 12), 1489 => to_unsigned(3662, 12), 1490 => to_unsigned(3226, 12), 1491 => to_unsigned(2952, 12), 1492 => to_unsigned(3528, 12), 1493 => to_unsigned(2125, 12), 1494 => to_unsigned(3864, 12), 1495 => to_unsigned(1887, 12), 1496 => to_unsigned(3376, 12), 1497 => to_unsigned(3925, 12), 1498 => to_unsigned(3189, 12), 1499 => to_unsigned(3179, 12), 1500 => to_unsigned(1600, 12), 1501 => to_unsigned(1102, 12), 1502 => to_unsigned(1756, 12), 1503 => to_unsigned(1312, 12), 1504 => to_unsigned(254, 12), 1505 => to_unsigned(315, 12), 1506 => to_unsigned(3521, 12), 1507 => to_unsigned(2551, 12), 1508 => to_unsigned(1782, 12), 1509 => to_unsigned(671, 12), 1510 => to_unsigned(597, 12), 1511 => to_unsigned(1738, 12), 1512 => to_unsigned(3903, 12), 1513 => to_unsigned(1432, 12), 1514 => to_unsigned(1679, 12), 1515 => to_unsigned(2112, 12), 1516 => to_unsigned(2681, 12), 1517 => to_unsigned(407, 12), 1518 => to_unsigned(3386, 12), 1519 => to_unsigned(2375, 12), 1520 => to_unsigned(2406, 12), 1521 => to_unsigned(2395, 12), 1522 => to_unsigned(1107, 12), 1523 => to_unsigned(2728, 12), 1524 => to_unsigned(681, 12), 1525 => to_unsigned(1787, 12), 1526 => to_unsigned(1490, 12), 1527 => to_unsigned(824, 12), 1528 => to_unsigned(2045, 12), 1529 => to_unsigned(3478, 12), 1530 => to_unsigned(2091, 12), 1531 => to_unsigned(444, 12), 1532 => to_unsigned(3854, 12), 1533 => to_unsigned(165, 12), 1534 => to_unsigned(3792, 12), 1535 => to_unsigned(96, 12), 1536 => to_unsigned(1255, 12), 1537 => to_unsigned(680, 12), 1538 => to_unsigned(3489, 12), 1539 => to_unsigned(800, 12), 1540 => to_unsigned(443, 12), 1541 => to_unsigned(1887, 12), 1542 => to_unsigned(4076, 12), 1543 => to_unsigned(1119, 12), 1544 => to_unsigned(1245, 12), 1545 => to_unsigned(284, 12), 1546 => to_unsigned(687, 12), 1547 => to_unsigned(3785, 12), 1548 => to_unsigned(1726, 12), 1549 => to_unsigned(243, 12), 1550 => to_unsigned(1049, 12), 1551 => to_unsigned(3159, 12), 1552 => to_unsigned(1697, 12), 1553 => to_unsigned(2544, 12), 1554 => to_unsigned(1186, 12), 1555 => to_unsigned(2213, 12), 1556 => to_unsigned(4057, 12), 1557 => to_unsigned(401, 12), 1558 => to_unsigned(2295, 12), 1559 => to_unsigned(3692, 12), 1560 => to_unsigned(3186, 12), 1561 => to_unsigned(3303, 12), 1562 => to_unsigned(3994, 12), 1563 => to_unsigned(2380, 12), 1564 => to_unsigned(973, 12), 1565 => to_unsigned(2278, 12), 1566 => to_unsigned(1372, 12), 1567 => to_unsigned(2409, 12), 1568 => to_unsigned(3378, 12), 1569 => to_unsigned(2993, 12), 1570 => to_unsigned(3736, 12), 1571 => to_unsigned(963, 12), 1572 => to_unsigned(3736, 12), 1573 => to_unsigned(3357, 12), 1574 => to_unsigned(3524, 12), 1575 => to_unsigned(4041, 12), 1576 => to_unsigned(2372, 12), 1577 => to_unsigned(1840, 12), 1578 => to_unsigned(1384, 12), 1579 => to_unsigned(1317, 12), 1580 => to_unsigned(762, 12), 1581 => to_unsigned(1730, 12), 1582 => to_unsigned(2134, 12), 1583 => to_unsigned(3127, 12), 1584 => to_unsigned(200, 12), 1585 => to_unsigned(3117, 12), 1586 => to_unsigned(2368, 12), 1587 => to_unsigned(59, 12), 1588 => to_unsigned(2501, 12), 1589 => to_unsigned(268, 12), 1590 => to_unsigned(955, 12), 1591 => to_unsigned(3602, 12), 1592 => to_unsigned(3914, 12), 1593 => to_unsigned(1819, 12), 1594 => to_unsigned(386, 12), 1595 => to_unsigned(3699, 12), 1596 => to_unsigned(1294, 12), 1597 => to_unsigned(879, 12), 1598 => to_unsigned(2417, 12), 1599 => to_unsigned(2016, 12), 1600 => to_unsigned(1414, 12), 1601 => to_unsigned(3644, 12), 1602 => to_unsigned(4092, 12), 1603 => to_unsigned(3204, 12), 1604 => to_unsigned(194, 12), 1605 => to_unsigned(2754, 12), 1606 => to_unsigned(2605, 12), 1607 => to_unsigned(3289, 12), 1608 => to_unsigned(1097, 12), 1609 => to_unsigned(2554, 12), 1610 => to_unsigned(2015, 12), 1611 => to_unsigned(2686, 12), 1612 => to_unsigned(2840, 12), 1613 => to_unsigned(2383, 12), 1614 => to_unsigned(530, 12), 1615 => to_unsigned(270, 12), 1616 => to_unsigned(2123, 12), 1617 => to_unsigned(3242, 12), 1618 => to_unsigned(751, 12), 1619 => to_unsigned(2464, 12), 1620 => to_unsigned(1101, 12), 1621 => to_unsigned(1934, 12), 1622 => to_unsigned(490, 12), 1623 => to_unsigned(2066, 12), 1624 => to_unsigned(1310, 12), 1625 => to_unsigned(1866, 12), 1626 => to_unsigned(951, 12), 1627 => to_unsigned(633, 12), 1628 => to_unsigned(738, 12), 1629 => to_unsigned(1709, 12), 1630 => to_unsigned(227, 12), 1631 => to_unsigned(2859, 12), 1632 => to_unsigned(878, 12), 1633 => to_unsigned(1109, 12), 1634 => to_unsigned(1620, 12), 1635 => to_unsigned(3606, 12), 1636 => to_unsigned(3535, 12), 1637 => to_unsigned(417, 12), 1638 => to_unsigned(1208, 12), 1639 => to_unsigned(4059, 12), 1640 => to_unsigned(2913, 12), 1641 => to_unsigned(2016, 12), 1642 => to_unsigned(859, 12), 1643 => to_unsigned(1632, 12), 1644 => to_unsigned(497, 12), 1645 => to_unsigned(2524, 12), 1646 => to_unsigned(3453, 12), 1647 => to_unsigned(773, 12), 1648 => to_unsigned(1556, 12), 1649 => to_unsigned(3453, 12), 1650 => to_unsigned(3721, 12), 1651 => to_unsigned(2661, 12), 1652 => to_unsigned(550, 12), 1653 => to_unsigned(3857, 12), 1654 => to_unsigned(262, 12), 1655 => to_unsigned(3524, 12), 1656 => to_unsigned(3274, 12), 1657 => to_unsigned(1118, 12), 1658 => to_unsigned(3074, 12), 1659 => to_unsigned(2926, 12), 1660 => to_unsigned(402, 12), 1661 => to_unsigned(3128, 12), 1662 => to_unsigned(3882, 12), 1663 => to_unsigned(3615, 12), 1664 => to_unsigned(3357, 12), 1665 => to_unsigned(1588, 12), 1666 => to_unsigned(2098, 12), 1667 => to_unsigned(1979, 12), 1668 => to_unsigned(3420, 12), 1669 => to_unsigned(356, 12), 1670 => to_unsigned(3890, 12), 1671 => to_unsigned(341, 12), 1672 => to_unsigned(1084, 12), 1673 => to_unsigned(3747, 12), 1674 => to_unsigned(3408, 12), 1675 => to_unsigned(3817, 12), 1676 => to_unsigned(273, 12), 1677 => to_unsigned(1819, 12), 1678 => to_unsigned(1747, 12), 1679 => to_unsigned(1101, 12), 1680 => to_unsigned(1697, 12), 1681 => to_unsigned(1753, 12), 1682 => to_unsigned(3725, 12), 1683 => to_unsigned(2940, 12), 1684 => to_unsigned(5, 12), 1685 => to_unsigned(2729, 12), 1686 => to_unsigned(565, 12), 1687 => to_unsigned(3672, 12), 1688 => to_unsigned(1132, 12), 1689 => to_unsigned(1282, 12), 1690 => to_unsigned(2761, 12), 1691 => to_unsigned(975, 12), 1692 => to_unsigned(2879, 12), 1693 => to_unsigned(2819, 12), 1694 => to_unsigned(61, 12), 1695 => to_unsigned(1216, 12), 1696 => to_unsigned(1068, 12), 1697 => to_unsigned(3920, 12), 1698 => to_unsigned(3682, 12), 1699 => to_unsigned(670, 12), 1700 => to_unsigned(1364, 12), 1701 => to_unsigned(614, 12), 1702 => to_unsigned(177, 12), 1703 => to_unsigned(3290, 12), 1704 => to_unsigned(3678, 12), 1705 => to_unsigned(1622, 12), 1706 => to_unsigned(2254, 12), 1707 => to_unsigned(2999, 12), 1708 => to_unsigned(1571, 12), 1709 => to_unsigned(3648, 12), 1710 => to_unsigned(2944, 12), 1711 => to_unsigned(3021, 12), 1712 => to_unsigned(1014, 12), 1713 => to_unsigned(1216, 12), 1714 => to_unsigned(1774, 12), 1715 => to_unsigned(60, 12), 1716 => to_unsigned(2888, 12), 1717 => to_unsigned(3790, 12), 1718 => to_unsigned(1800, 12), 1719 => to_unsigned(2801, 12), 1720 => to_unsigned(3945, 12), 1721 => to_unsigned(4089, 12), 1722 => to_unsigned(2945, 12), 1723 => to_unsigned(1473, 12), 1724 => to_unsigned(3458, 12), 1725 => to_unsigned(3343, 12), 1726 => to_unsigned(149, 12), 1727 => to_unsigned(942, 12), 1728 => to_unsigned(3330, 12), 1729 => to_unsigned(1872, 12), 1730 => to_unsigned(993, 12), 1731 => to_unsigned(720, 12), 1732 => to_unsigned(3226, 12), 1733 => to_unsigned(1095, 12), 1734 => to_unsigned(1776, 12), 1735 => to_unsigned(3981, 12), 1736 => to_unsigned(739, 12), 1737 => to_unsigned(1156, 12), 1738 => to_unsigned(1450, 12), 1739 => to_unsigned(2758, 12), 1740 => to_unsigned(2730, 12), 1741 => to_unsigned(2811, 12), 1742 => to_unsigned(1740, 12), 1743 => to_unsigned(2401, 12), 1744 => to_unsigned(204, 12), 1745 => to_unsigned(2110, 12), 1746 => to_unsigned(1395, 12), 1747 => to_unsigned(3756, 12), 1748 => to_unsigned(3299, 12), 1749 => to_unsigned(3533, 12), 1750 => to_unsigned(726, 12), 1751 => to_unsigned(1079, 12), 1752 => to_unsigned(1559, 12), 1753 => to_unsigned(3659, 12), 1754 => to_unsigned(609, 12), 1755 => to_unsigned(2985, 12), 1756 => to_unsigned(1788, 12), 1757 => to_unsigned(2830, 12), 1758 => to_unsigned(3353, 12), 1759 => to_unsigned(746, 12), 1760 => to_unsigned(1038, 12), 1761 => to_unsigned(3180, 12), 1762 => to_unsigned(1656, 12), 1763 => to_unsigned(671, 12), 1764 => to_unsigned(1628, 12), 1765 => to_unsigned(1774, 12), 1766 => to_unsigned(2510, 12), 1767 => to_unsigned(114, 12), 1768 => to_unsigned(3208, 12), 1769 => to_unsigned(1814, 12), 1770 => to_unsigned(124, 12), 1771 => to_unsigned(110, 12), 1772 => to_unsigned(2947, 12), 1773 => to_unsigned(1539, 12), 1774 => to_unsigned(3117, 12), 1775 => to_unsigned(1144, 12), 1776 => to_unsigned(213, 12), 1777 => to_unsigned(2815, 12), 1778 => to_unsigned(2519, 12), 1779 => to_unsigned(3751, 12), 1780 => to_unsigned(2408, 12), 1781 => to_unsigned(129, 12), 1782 => to_unsigned(964, 12), 1783 => to_unsigned(1322, 12), 1784 => to_unsigned(1424, 12), 1785 => to_unsigned(784, 12), 1786 => to_unsigned(2286, 12), 1787 => to_unsigned(4001, 12), 1788 => to_unsigned(1236, 12), 1789 => to_unsigned(1625, 12), 1790 => to_unsigned(1408, 12), 1791 => to_unsigned(2499, 12), 1792 => to_unsigned(256, 12), 1793 => to_unsigned(773, 12), 1794 => to_unsigned(713, 12), 1795 => to_unsigned(2493, 12), 1796 => to_unsigned(3189, 12), 1797 => to_unsigned(3010, 12), 1798 => to_unsigned(1108, 12), 1799 => to_unsigned(1111, 12), 1800 => to_unsigned(3821, 12), 1801 => to_unsigned(3633, 12), 1802 => to_unsigned(2186, 12), 1803 => to_unsigned(155, 12), 1804 => to_unsigned(3898, 12), 1805 => to_unsigned(42, 12), 1806 => to_unsigned(1580, 12), 1807 => to_unsigned(3325, 12), 1808 => to_unsigned(253, 12), 1809 => to_unsigned(550, 12), 1810 => to_unsigned(3724, 12), 1811 => to_unsigned(138, 12), 1812 => to_unsigned(1121, 12), 1813 => to_unsigned(3360, 12), 1814 => to_unsigned(3471, 12), 1815 => to_unsigned(1328, 12), 1816 => to_unsigned(1071, 12), 1817 => to_unsigned(4057, 12), 1818 => to_unsigned(1182, 12), 1819 => to_unsigned(1558, 12), 1820 => to_unsigned(3763, 12), 1821 => to_unsigned(1329, 12), 1822 => to_unsigned(936, 12), 1823 => to_unsigned(1932, 12), 1824 => to_unsigned(460, 12), 1825 => to_unsigned(2228, 12), 1826 => to_unsigned(3191, 12), 1827 => to_unsigned(524, 12), 1828 => to_unsigned(2588, 12), 1829 => to_unsigned(749, 12), 1830 => to_unsigned(2130, 12), 1831 => to_unsigned(1715, 12), 1832 => to_unsigned(2268, 12), 1833 => to_unsigned(171, 12), 1834 => to_unsigned(3883, 12), 1835 => to_unsigned(1066, 12), 1836 => to_unsigned(2171, 12), 1837 => to_unsigned(1478, 12), 1838 => to_unsigned(2870, 12), 1839 => to_unsigned(2009, 12), 1840 => to_unsigned(1560, 12), 1841 => to_unsigned(1796, 12), 1842 => to_unsigned(1886, 12), 1843 => to_unsigned(1596, 12), 1844 => to_unsigned(972, 12), 1845 => to_unsigned(1806, 12), 1846 => to_unsigned(3254, 12), 1847 => to_unsigned(562, 12), 1848 => to_unsigned(655, 12), 1849 => to_unsigned(103, 12), 1850 => to_unsigned(688, 12), 1851 => to_unsigned(1164, 12), 1852 => to_unsigned(3992, 12), 1853 => to_unsigned(479, 12), 1854 => to_unsigned(3537, 12), 1855 => to_unsigned(582, 12), 1856 => to_unsigned(2439, 12), 1857 => to_unsigned(3977, 12), 1858 => to_unsigned(332, 12), 1859 => to_unsigned(1588, 12), 1860 => to_unsigned(785, 12), 1861 => to_unsigned(3493, 12), 1862 => to_unsigned(2999, 12), 1863 => to_unsigned(729, 12), 1864 => to_unsigned(2120, 12), 1865 => to_unsigned(3966, 12), 1866 => to_unsigned(2581, 12), 1867 => to_unsigned(1297, 12), 1868 => to_unsigned(2116, 12), 1869 => to_unsigned(925, 12), 1870 => to_unsigned(421, 12), 1871 => to_unsigned(1177, 12), 1872 => to_unsigned(3272, 12), 1873 => to_unsigned(999, 12), 1874 => to_unsigned(11, 12), 1875 => to_unsigned(2647, 12), 1876 => to_unsigned(3163, 12), 1877 => to_unsigned(3984, 12), 1878 => to_unsigned(3016, 12), 1879 => to_unsigned(1044, 12), 1880 => to_unsigned(1313, 12), 1881 => to_unsigned(537, 12), 1882 => to_unsigned(2382, 12), 1883 => to_unsigned(1161, 12), 1884 => to_unsigned(2969, 12), 1885 => to_unsigned(2756, 12), 1886 => to_unsigned(3430, 12), 1887 => to_unsigned(3169, 12), 1888 => to_unsigned(2292, 12), 1889 => to_unsigned(2304, 12), 1890 => to_unsigned(296, 12), 1891 => to_unsigned(3789, 12), 1892 => to_unsigned(2766, 12), 1893 => to_unsigned(715, 12), 1894 => to_unsigned(5, 12), 1895 => to_unsigned(3096, 12), 1896 => to_unsigned(3323, 12), 1897 => to_unsigned(3853, 12), 1898 => to_unsigned(2426, 12), 1899 => to_unsigned(3818, 12), 1900 => to_unsigned(1730, 12), 1901 => to_unsigned(2946, 12), 1902 => to_unsigned(1929, 12), 1903 => to_unsigned(4064, 12), 1904 => to_unsigned(1729, 12), 1905 => to_unsigned(237, 12), 1906 => to_unsigned(750, 12), 1907 => to_unsigned(4092, 12), 1908 => to_unsigned(2087, 12), 1909 => to_unsigned(3137, 12), 1910 => to_unsigned(1874, 12), 1911 => to_unsigned(2039, 12), 1912 => to_unsigned(922, 12), 1913 => to_unsigned(681, 12), 1914 => to_unsigned(3151, 12), 1915 => to_unsigned(2695, 12), 1916 => to_unsigned(771, 12), 1917 => to_unsigned(1903, 12), 1918 => to_unsigned(2169, 12), 1919 => to_unsigned(2984, 12), 1920 => to_unsigned(164, 12), 1921 => to_unsigned(2861, 12), 1922 => to_unsigned(2080, 12), 1923 => to_unsigned(3662, 12), 1924 => to_unsigned(3885, 12), 1925 => to_unsigned(1326, 12), 1926 => to_unsigned(1189, 12), 1927 => to_unsigned(2036, 12), 1928 => to_unsigned(2020, 12), 1929 => to_unsigned(414, 12), 1930 => to_unsigned(1675, 12), 1931 => to_unsigned(1364, 12), 1932 => to_unsigned(3446, 12), 1933 => to_unsigned(1961, 12), 1934 => to_unsigned(2788, 12), 1935 => to_unsigned(3831, 12), 1936 => to_unsigned(1944, 12), 1937 => to_unsigned(1008, 12), 1938 => to_unsigned(3370, 12), 1939 => to_unsigned(3880, 12), 1940 => to_unsigned(2059, 12), 1941 => to_unsigned(2593, 12), 1942 => to_unsigned(2856, 12), 1943 => to_unsigned(1709, 12), 1944 => to_unsigned(819, 12), 1945 => to_unsigned(1526, 12), 1946 => to_unsigned(1044, 12), 1947 => to_unsigned(1940, 12), 1948 => to_unsigned(3042, 12), 1949 => to_unsigned(332, 12), 1950 => to_unsigned(2705, 12), 1951 => to_unsigned(7, 12), 1952 => to_unsigned(1093, 12), 1953 => to_unsigned(840, 12), 1954 => to_unsigned(1711, 12), 1955 => to_unsigned(3875, 12), 1956 => to_unsigned(3506, 12), 1957 => to_unsigned(1911, 12), 1958 => to_unsigned(3964, 12), 1959 => to_unsigned(1981, 12), 1960 => to_unsigned(622, 12), 1961 => to_unsigned(683, 12), 1962 => to_unsigned(3620, 12), 1963 => to_unsigned(926, 12), 1964 => to_unsigned(2432, 12), 1965 => to_unsigned(3226, 12), 1966 => to_unsigned(370, 12), 1967 => to_unsigned(2911, 12), 1968 => to_unsigned(2053, 12), 1969 => to_unsigned(1964, 12), 1970 => to_unsigned(3747, 12), 1971 => to_unsigned(2165, 12), 1972 => to_unsigned(1862, 12), 1973 => to_unsigned(722, 12), 1974 => to_unsigned(2712, 12), 1975 => to_unsigned(532, 12), 1976 => to_unsigned(1483, 12), 1977 => to_unsigned(3562, 12), 1978 => to_unsigned(4075, 12), 1979 => to_unsigned(2836, 12), 1980 => to_unsigned(812, 12), 1981 => to_unsigned(276, 12), 1982 => to_unsigned(3677, 12), 1983 => to_unsigned(117, 12), 1984 => to_unsigned(2744, 12), 1985 => to_unsigned(1998, 12), 1986 => to_unsigned(2112, 12), 1987 => to_unsigned(3759, 12), 1988 => to_unsigned(2634, 12), 1989 => to_unsigned(1406, 12), 1990 => to_unsigned(2677, 12), 1991 => to_unsigned(1270, 12), 1992 => to_unsigned(1458, 12), 1993 => to_unsigned(2331, 12), 1994 => to_unsigned(1750, 12), 1995 => to_unsigned(2345, 12), 1996 => to_unsigned(1202, 12), 1997 => to_unsigned(1799, 12), 1998 => to_unsigned(200, 12), 1999 => to_unsigned(1773, 12), 2000 => to_unsigned(3104, 12), 2001 => to_unsigned(545, 12), 2002 => to_unsigned(825, 12), 2003 => to_unsigned(1238, 12), 2004 => to_unsigned(3097, 12), 2005 => to_unsigned(3672, 12), 2006 => to_unsigned(2174, 12), 2007 => to_unsigned(2643, 12), 2008 => to_unsigned(2584, 12), 2009 => to_unsigned(127, 12), 2010 => to_unsigned(2411, 12), 2011 => to_unsigned(3002, 12), 2012 => to_unsigned(1055, 12), 2013 => to_unsigned(2880, 12), 2014 => to_unsigned(2238, 12), 2015 => to_unsigned(617, 12), 2016 => to_unsigned(3395, 12), 2017 => to_unsigned(3953, 12), 2018 => to_unsigned(3493, 12), 2019 => to_unsigned(3581, 12), 2020 => to_unsigned(425, 12), 2021 => to_unsigned(1654, 12), 2022 => to_unsigned(1712, 12), 2023 => to_unsigned(3180, 12), 2024 => to_unsigned(3337, 12), 2025 => to_unsigned(3005, 12), 2026 => to_unsigned(1663, 12), 2027 => to_unsigned(2101, 12), 2028 => to_unsigned(1876, 12), 2029 => to_unsigned(1709, 12), 2030 => to_unsigned(792, 12), 2031 => to_unsigned(3366, 12), 2032 => to_unsigned(247, 12), 2033 => to_unsigned(2595, 12), 2034 => to_unsigned(1404, 12), 2035 => to_unsigned(1605, 12), 2036 => to_unsigned(934, 12), 2037 => to_unsigned(227, 12), 2038 => to_unsigned(2916, 12), 2039 => to_unsigned(581, 12), 2040 => to_unsigned(1305, 12), 2041 => to_unsigned(2404, 12), 2042 => to_unsigned(1400, 12), 2043 => to_unsigned(3087, 12), 2044 => to_unsigned(2305, 12), 2045 => to_unsigned(3326, 12), 2046 => to_unsigned(1206, 12), 2047 => to_unsigned(2849, 12)),
            9 => (0 => to_unsigned(1735, 12), 1 => to_unsigned(558, 12), 2 => to_unsigned(477, 12), 3 => to_unsigned(1114, 12), 4 => to_unsigned(2232, 12), 5 => to_unsigned(2138, 12), 6 => to_unsigned(3467, 12), 7 => to_unsigned(1701, 12), 8 => to_unsigned(1475, 12), 9 => to_unsigned(153, 12), 10 => to_unsigned(3296, 12), 11 => to_unsigned(3716, 12), 12 => to_unsigned(3136, 12), 13 => to_unsigned(3608, 12), 14 => to_unsigned(3590, 12), 15 => to_unsigned(132, 12), 16 => to_unsigned(2464, 12), 17 => to_unsigned(2667, 12), 18 => to_unsigned(3416, 12), 19 => to_unsigned(1531, 12), 20 => to_unsigned(627, 12), 21 => to_unsigned(3924, 12), 22 => to_unsigned(3761, 12), 23 => to_unsigned(2875, 12), 24 => to_unsigned(3978, 12), 25 => to_unsigned(3412, 12), 26 => to_unsigned(609, 12), 27 => to_unsigned(2627, 12), 28 => to_unsigned(1678, 12), 29 => to_unsigned(3178, 12), 30 => to_unsigned(964, 12), 31 => to_unsigned(1616, 12), 32 => to_unsigned(1027, 12), 33 => to_unsigned(1782, 12), 34 => to_unsigned(3653, 12), 35 => to_unsigned(1464, 12), 36 => to_unsigned(3076, 12), 37 => to_unsigned(627, 12), 38 => to_unsigned(3542, 12), 39 => to_unsigned(540, 12), 40 => to_unsigned(1, 12), 41 => to_unsigned(3976, 12), 42 => to_unsigned(1254, 12), 43 => to_unsigned(2664, 12), 44 => to_unsigned(3530, 12), 45 => to_unsigned(1252, 12), 46 => to_unsigned(847, 12), 47 => to_unsigned(831, 12), 48 => to_unsigned(188, 12), 49 => to_unsigned(1929, 12), 50 => to_unsigned(2630, 12), 51 => to_unsigned(599, 12), 52 => to_unsigned(3962, 12), 53 => to_unsigned(2804, 12), 54 => to_unsigned(2140, 12), 55 => to_unsigned(107, 12), 56 => to_unsigned(3091, 12), 57 => to_unsigned(1428, 12), 58 => to_unsigned(2391, 12), 59 => to_unsigned(4074, 12), 60 => to_unsigned(2024, 12), 61 => to_unsigned(3368, 12), 62 => to_unsigned(3533, 12), 63 => to_unsigned(947, 12), 64 => to_unsigned(1402, 12), 65 => to_unsigned(947, 12), 66 => to_unsigned(3044, 12), 67 => to_unsigned(987, 12), 68 => to_unsigned(2151, 12), 69 => to_unsigned(1382, 12), 70 => to_unsigned(2008, 12), 71 => to_unsigned(2546, 12), 72 => to_unsigned(2294, 12), 73 => to_unsigned(4080, 12), 74 => to_unsigned(1387, 12), 75 => to_unsigned(1626, 12), 76 => to_unsigned(3310, 12), 77 => to_unsigned(789, 12), 78 => to_unsigned(3150, 12), 79 => to_unsigned(1779, 12), 80 => to_unsigned(2167, 12), 81 => to_unsigned(2553, 12), 82 => to_unsigned(652, 12), 83 => to_unsigned(204, 12), 84 => to_unsigned(156, 12), 85 => to_unsigned(3118, 12), 86 => to_unsigned(2722, 12), 87 => to_unsigned(1739, 12), 88 => to_unsigned(2410, 12), 89 => to_unsigned(784, 12), 90 => to_unsigned(3369, 12), 91 => to_unsigned(973, 12), 92 => to_unsigned(2599, 12), 93 => to_unsigned(3157, 12), 94 => to_unsigned(3311, 12), 95 => to_unsigned(3976, 12), 96 => to_unsigned(2617, 12), 97 => to_unsigned(2189, 12), 98 => to_unsigned(3357, 12), 99 => to_unsigned(676, 12), 100 => to_unsigned(1502, 12), 101 => to_unsigned(3063, 12), 102 => to_unsigned(3501, 12), 103 => to_unsigned(1049, 12), 104 => to_unsigned(3854, 12), 105 => to_unsigned(1383, 12), 106 => to_unsigned(6, 12), 107 => to_unsigned(1508, 12), 108 => to_unsigned(3679, 12), 109 => to_unsigned(3966, 12), 110 => to_unsigned(1320, 12), 111 => to_unsigned(729, 12), 112 => to_unsigned(1901, 12), 113 => to_unsigned(1135, 12), 114 => to_unsigned(3616, 12), 115 => to_unsigned(3032, 12), 116 => to_unsigned(161, 12), 117 => to_unsigned(2543, 12), 118 => to_unsigned(2474, 12), 119 => to_unsigned(281, 12), 120 => to_unsigned(3484, 12), 121 => to_unsigned(2637, 12), 122 => to_unsigned(931, 12), 123 => to_unsigned(419, 12), 124 => to_unsigned(2250, 12), 125 => to_unsigned(2034, 12), 126 => to_unsigned(2072, 12), 127 => to_unsigned(1186, 12), 128 => to_unsigned(3815, 12), 129 => to_unsigned(695, 12), 130 => to_unsigned(1873, 12), 131 => to_unsigned(3836, 12), 132 => to_unsigned(2334, 12), 133 => to_unsigned(1780, 12), 134 => to_unsigned(2798, 12), 135 => to_unsigned(2788, 12), 136 => to_unsigned(1211, 12), 137 => to_unsigned(1374, 12), 138 => to_unsigned(1152, 12), 139 => to_unsigned(2704, 12), 140 => to_unsigned(3654, 12), 141 => to_unsigned(1560, 12), 142 => to_unsigned(350, 12), 143 => to_unsigned(3512, 12), 144 => to_unsigned(2395, 12), 145 => to_unsigned(2659, 12), 146 => to_unsigned(287, 12), 147 => to_unsigned(2259, 12), 148 => to_unsigned(2658, 12), 149 => to_unsigned(3655, 12), 150 => to_unsigned(3480, 12), 151 => to_unsigned(2903, 12), 152 => to_unsigned(1154, 12), 153 => to_unsigned(4018, 12), 154 => to_unsigned(925, 12), 155 => to_unsigned(805, 12), 156 => to_unsigned(100, 12), 157 => to_unsigned(1856, 12), 158 => to_unsigned(3409, 12), 159 => to_unsigned(2450, 12), 160 => to_unsigned(1608, 12), 161 => to_unsigned(3974, 12), 162 => to_unsigned(630, 12), 163 => to_unsigned(1744, 12), 164 => to_unsigned(1440, 12), 165 => to_unsigned(2210, 12), 166 => to_unsigned(3850, 12), 167 => to_unsigned(2880, 12), 168 => to_unsigned(3667, 12), 169 => to_unsigned(300, 12), 170 => to_unsigned(2490, 12), 171 => to_unsigned(2206, 12), 172 => to_unsigned(482, 12), 173 => to_unsigned(1095, 12), 174 => to_unsigned(3587, 12), 175 => to_unsigned(1736, 12), 176 => to_unsigned(907, 12), 177 => to_unsigned(1027, 12), 178 => to_unsigned(2934, 12), 179 => to_unsigned(3024, 12), 180 => to_unsigned(341, 12), 181 => to_unsigned(3706, 12), 182 => to_unsigned(2015, 12), 183 => to_unsigned(3042, 12), 184 => to_unsigned(1048, 12), 185 => to_unsigned(3428, 12), 186 => to_unsigned(1215, 12), 187 => to_unsigned(2847, 12), 188 => to_unsigned(505, 12), 189 => to_unsigned(3707, 12), 190 => to_unsigned(392, 12), 191 => to_unsigned(849, 12), 192 => to_unsigned(3614, 12), 193 => to_unsigned(1062, 12), 194 => to_unsigned(3836, 12), 195 => to_unsigned(1699, 12), 196 => to_unsigned(2616, 12), 197 => to_unsigned(3741, 12), 198 => to_unsigned(1680, 12), 199 => to_unsigned(755, 12), 200 => to_unsigned(2483, 12), 201 => to_unsigned(554, 12), 202 => to_unsigned(1510, 12), 203 => to_unsigned(1695, 12), 204 => to_unsigned(3491, 12), 205 => to_unsigned(1532, 12), 206 => to_unsigned(1486, 12), 207 => to_unsigned(3650, 12), 208 => to_unsigned(3778, 12), 209 => to_unsigned(1346, 12), 210 => to_unsigned(1396, 12), 211 => to_unsigned(1467, 12), 212 => to_unsigned(2152, 12), 213 => to_unsigned(688, 12), 214 => to_unsigned(3413, 12), 215 => to_unsigned(2466, 12), 216 => to_unsigned(360, 12), 217 => to_unsigned(3930, 12), 218 => to_unsigned(2907, 12), 219 => to_unsigned(1419, 12), 220 => to_unsigned(1683, 12), 221 => to_unsigned(2994, 12), 222 => to_unsigned(804, 12), 223 => to_unsigned(1899, 12), 224 => to_unsigned(367, 12), 225 => to_unsigned(1236, 12), 226 => to_unsigned(1396, 12), 227 => to_unsigned(3872, 12), 228 => to_unsigned(3363, 12), 229 => to_unsigned(1771, 12), 230 => to_unsigned(3957, 12), 231 => to_unsigned(3100, 12), 232 => to_unsigned(1465, 12), 233 => to_unsigned(433, 12), 234 => to_unsigned(2426, 12), 235 => to_unsigned(1201, 12), 236 => to_unsigned(2858, 12), 237 => to_unsigned(3029, 12), 238 => to_unsigned(2983, 12), 239 => to_unsigned(2740, 12), 240 => to_unsigned(3663, 12), 241 => to_unsigned(1563, 12), 242 => to_unsigned(2850, 12), 243 => to_unsigned(959, 12), 244 => to_unsigned(1098, 12), 245 => to_unsigned(2639, 12), 246 => to_unsigned(3344, 12), 247 => to_unsigned(867, 12), 248 => to_unsigned(543, 12), 249 => to_unsigned(2862, 12), 250 => to_unsigned(171, 12), 251 => to_unsigned(2117, 12), 252 => to_unsigned(322, 12), 253 => to_unsigned(258, 12), 254 => to_unsigned(3987, 12), 255 => to_unsigned(2462, 12), 256 => to_unsigned(2681, 12), 257 => to_unsigned(805, 12), 258 => to_unsigned(1960, 12), 259 => to_unsigned(257, 12), 260 => to_unsigned(2151, 12), 261 => to_unsigned(1461, 12), 262 => to_unsigned(2820, 12), 263 => to_unsigned(2594, 12), 264 => to_unsigned(277, 12), 265 => to_unsigned(3562, 12), 266 => to_unsigned(179, 12), 267 => to_unsigned(1740, 12), 268 => to_unsigned(1761, 12), 269 => to_unsigned(2038, 12), 270 => to_unsigned(2996, 12), 271 => to_unsigned(3849, 12), 272 => to_unsigned(229, 12), 273 => to_unsigned(3859, 12), 274 => to_unsigned(3697, 12), 275 => to_unsigned(3167, 12), 276 => to_unsigned(3053, 12), 277 => to_unsigned(2116, 12), 278 => to_unsigned(5, 12), 279 => to_unsigned(1115, 12), 280 => to_unsigned(2150, 12), 281 => to_unsigned(2485, 12), 282 => to_unsigned(977, 12), 283 => to_unsigned(3918, 12), 284 => to_unsigned(2409, 12), 285 => to_unsigned(1864, 12), 286 => to_unsigned(2257, 12), 287 => to_unsigned(1232, 12), 288 => to_unsigned(1988, 12), 289 => to_unsigned(237, 12), 290 => to_unsigned(1065, 12), 291 => to_unsigned(1437, 12), 292 => to_unsigned(2224, 12), 293 => to_unsigned(667, 12), 294 => to_unsigned(3650, 12), 295 => to_unsigned(3428, 12), 296 => to_unsigned(603, 12), 297 => to_unsigned(4021, 12), 298 => to_unsigned(687, 12), 299 => to_unsigned(1147, 12), 300 => to_unsigned(581, 12), 301 => to_unsigned(1774, 12), 302 => to_unsigned(1788, 12), 303 => to_unsigned(3547, 12), 304 => to_unsigned(3573, 12), 305 => to_unsigned(2171, 12), 306 => to_unsigned(912, 12), 307 => to_unsigned(1202, 12), 308 => to_unsigned(2787, 12), 309 => to_unsigned(682, 12), 310 => to_unsigned(2688, 12), 311 => to_unsigned(332, 12), 312 => to_unsigned(2311, 12), 313 => to_unsigned(3674, 12), 314 => to_unsigned(656, 12), 315 => to_unsigned(1720, 12), 316 => to_unsigned(1120, 12), 317 => to_unsigned(3031, 12), 318 => to_unsigned(1850, 12), 319 => to_unsigned(15, 12), 320 => to_unsigned(185, 12), 321 => to_unsigned(3499, 12), 322 => to_unsigned(1405, 12), 323 => to_unsigned(1368, 12), 324 => to_unsigned(3558, 12), 325 => to_unsigned(1292, 12), 326 => to_unsigned(2409, 12), 327 => to_unsigned(2273, 12), 328 => to_unsigned(2696, 12), 329 => to_unsigned(2716, 12), 330 => to_unsigned(139, 12), 331 => to_unsigned(3744, 12), 332 => to_unsigned(2637, 12), 333 => to_unsigned(1362, 12), 334 => to_unsigned(3661, 12), 335 => to_unsigned(1542, 12), 336 => to_unsigned(2770, 12), 337 => to_unsigned(4075, 12), 338 => to_unsigned(2764, 12), 339 => to_unsigned(1871, 12), 340 => to_unsigned(890, 12), 341 => to_unsigned(661, 12), 342 => to_unsigned(1961, 12), 343 => to_unsigned(3604, 12), 344 => to_unsigned(3802, 12), 345 => to_unsigned(145, 12), 346 => to_unsigned(2117, 12), 347 => to_unsigned(3036, 12), 348 => to_unsigned(32, 12), 349 => to_unsigned(1431, 12), 350 => to_unsigned(3118, 12), 351 => to_unsigned(3098, 12), 352 => to_unsigned(1164, 12), 353 => to_unsigned(2444, 12), 354 => to_unsigned(2819, 12), 355 => to_unsigned(3278, 12), 356 => to_unsigned(462, 12), 357 => to_unsigned(32, 12), 358 => to_unsigned(1548, 12), 359 => to_unsigned(545, 12), 360 => to_unsigned(3356, 12), 361 => to_unsigned(2701, 12), 362 => to_unsigned(2684, 12), 363 => to_unsigned(1612, 12), 364 => to_unsigned(287, 12), 365 => to_unsigned(975, 12), 366 => to_unsigned(3180, 12), 367 => to_unsigned(703, 12), 368 => to_unsigned(1623, 12), 369 => to_unsigned(92, 12), 370 => to_unsigned(2777, 12), 371 => to_unsigned(1322, 12), 372 => to_unsigned(2050, 12), 373 => to_unsigned(3290, 12), 374 => to_unsigned(3545, 12), 375 => to_unsigned(871, 12), 376 => to_unsigned(760, 12), 377 => to_unsigned(1902, 12), 378 => to_unsigned(2728, 12), 379 => to_unsigned(1004, 12), 380 => to_unsigned(1729, 12), 381 => to_unsigned(2995, 12), 382 => to_unsigned(3901, 12), 383 => to_unsigned(1637, 12), 384 => to_unsigned(2743, 12), 385 => to_unsigned(1622, 12), 386 => to_unsigned(3791, 12), 387 => to_unsigned(2247, 12), 388 => to_unsigned(3964, 12), 389 => to_unsigned(3814, 12), 390 => to_unsigned(1723, 12), 391 => to_unsigned(676, 12), 392 => to_unsigned(2870, 12), 393 => to_unsigned(3671, 12), 394 => to_unsigned(3456, 12), 395 => to_unsigned(535, 12), 396 => to_unsigned(2755, 12), 397 => to_unsigned(3463, 12), 398 => to_unsigned(3732, 12), 399 => to_unsigned(2808, 12), 400 => to_unsigned(1650, 12), 401 => to_unsigned(2966, 12), 402 => to_unsigned(1138, 12), 403 => to_unsigned(358, 12), 404 => to_unsigned(2910, 12), 405 => to_unsigned(3611, 12), 406 => to_unsigned(1451, 12), 407 => to_unsigned(3195, 12), 408 => to_unsigned(1089, 12), 409 => to_unsigned(2075, 12), 410 => to_unsigned(2271, 12), 411 => to_unsigned(1862, 12), 412 => to_unsigned(935, 12), 413 => to_unsigned(501, 12), 414 => to_unsigned(52, 12), 415 => to_unsigned(2437, 12), 416 => to_unsigned(82, 12), 417 => to_unsigned(3656, 12), 418 => to_unsigned(870, 12), 419 => to_unsigned(1428, 12), 420 => to_unsigned(89, 12), 421 => to_unsigned(3170, 12), 422 => to_unsigned(3471, 12), 423 => to_unsigned(2560, 12), 424 => to_unsigned(3538, 12), 425 => to_unsigned(32, 12), 426 => to_unsigned(3252, 12), 427 => to_unsigned(2755, 12), 428 => to_unsigned(1789, 12), 429 => to_unsigned(3283, 12), 430 => to_unsigned(118, 12), 431 => to_unsigned(3375, 12), 432 => to_unsigned(1661, 12), 433 => to_unsigned(2836, 12), 434 => to_unsigned(987, 12), 435 => to_unsigned(1708, 12), 436 => to_unsigned(2288, 12), 437 => to_unsigned(743, 12), 438 => to_unsigned(3598, 12), 439 => to_unsigned(1636, 12), 440 => to_unsigned(421, 12), 441 => to_unsigned(3999, 12), 442 => to_unsigned(1671, 12), 443 => to_unsigned(2649, 12), 444 => to_unsigned(2754, 12), 445 => to_unsigned(248, 12), 446 => to_unsigned(3483, 12), 447 => to_unsigned(244, 12), 448 => to_unsigned(3912, 12), 449 => to_unsigned(1309, 12), 450 => to_unsigned(2954, 12), 451 => to_unsigned(3969, 12), 452 => to_unsigned(1867, 12), 453 => to_unsigned(1600, 12), 454 => to_unsigned(1319, 12), 455 => to_unsigned(2523, 12), 456 => to_unsigned(3919, 12), 457 => to_unsigned(526, 12), 458 => to_unsigned(245, 12), 459 => to_unsigned(4072, 12), 460 => to_unsigned(2398, 12), 461 => to_unsigned(9, 12), 462 => to_unsigned(256, 12), 463 => to_unsigned(2218, 12), 464 => to_unsigned(3191, 12), 465 => to_unsigned(3261, 12), 466 => to_unsigned(1931, 12), 467 => to_unsigned(1940, 12), 468 => to_unsigned(4006, 12), 469 => to_unsigned(1567, 12), 470 => to_unsigned(3471, 12), 471 => to_unsigned(1024, 12), 472 => to_unsigned(1256, 12), 473 => to_unsigned(930, 12), 474 => to_unsigned(1840, 12), 475 => to_unsigned(1175, 12), 476 => to_unsigned(1991, 12), 477 => to_unsigned(446, 12), 478 => to_unsigned(446, 12), 479 => to_unsigned(1770, 12), 480 => to_unsigned(2085, 12), 481 => to_unsigned(856, 12), 482 => to_unsigned(2204, 12), 483 => to_unsigned(208, 12), 484 => to_unsigned(3762, 12), 485 => to_unsigned(1023, 12), 486 => to_unsigned(2890, 12), 487 => to_unsigned(366, 12), 488 => to_unsigned(4053, 12), 489 => to_unsigned(1357, 12), 490 => to_unsigned(92, 12), 491 => to_unsigned(1012, 12), 492 => to_unsigned(1318, 12), 493 => to_unsigned(1508, 12), 494 => to_unsigned(3334, 12), 495 => to_unsigned(1224, 12), 496 => to_unsigned(934, 12), 497 => to_unsigned(3451, 12), 498 => to_unsigned(1255, 12), 499 => to_unsigned(1060, 12), 500 => to_unsigned(1821, 12), 501 => to_unsigned(2747, 12), 502 => to_unsigned(2428, 12), 503 => to_unsigned(2700, 12), 504 => to_unsigned(2639, 12), 505 => to_unsigned(3977, 12), 506 => to_unsigned(2033, 12), 507 => to_unsigned(2980, 12), 508 => to_unsigned(153, 12), 509 => to_unsigned(2829, 12), 510 => to_unsigned(3761, 12), 511 => to_unsigned(582, 12), 512 => to_unsigned(2418, 12), 513 => to_unsigned(613, 12), 514 => to_unsigned(2974, 12), 515 => to_unsigned(433, 12), 516 => to_unsigned(3091, 12), 517 => to_unsigned(1564, 12), 518 => to_unsigned(972, 12), 519 => to_unsigned(1659, 12), 520 => to_unsigned(1064, 12), 521 => to_unsigned(3060, 12), 522 => to_unsigned(608, 12), 523 => to_unsigned(2297, 12), 524 => to_unsigned(865, 12), 525 => to_unsigned(2508, 12), 526 => to_unsigned(3895, 12), 527 => to_unsigned(2853, 12), 528 => to_unsigned(2064, 12), 529 => to_unsigned(722, 12), 530 => to_unsigned(3869, 12), 531 => to_unsigned(151, 12), 532 => to_unsigned(4020, 12), 533 => to_unsigned(3732, 12), 534 => to_unsigned(2303, 12), 535 => to_unsigned(855, 12), 536 => to_unsigned(1281, 12), 537 => to_unsigned(1779, 12), 538 => to_unsigned(2731, 12), 539 => to_unsigned(3352, 12), 540 => to_unsigned(1527, 12), 541 => to_unsigned(2205, 12), 542 => to_unsigned(1954, 12), 543 => to_unsigned(2157, 12), 544 => to_unsigned(4073, 12), 545 => to_unsigned(3954, 12), 546 => to_unsigned(2502, 12), 547 => to_unsigned(98, 12), 548 => to_unsigned(3275, 12), 549 => to_unsigned(3680, 12), 550 => to_unsigned(3459, 12), 551 => to_unsigned(2674, 12), 552 => to_unsigned(1105, 12), 553 => to_unsigned(3784, 12), 554 => to_unsigned(3884, 12), 555 => to_unsigned(1242, 12), 556 => to_unsigned(1082, 12), 557 => to_unsigned(3274, 12), 558 => to_unsigned(848, 12), 559 => to_unsigned(1626, 12), 560 => to_unsigned(2863, 12), 561 => to_unsigned(3087, 12), 562 => to_unsigned(2690, 12), 563 => to_unsigned(2714, 12), 564 => to_unsigned(1978, 12), 565 => to_unsigned(3350, 12), 566 => to_unsigned(1356, 12), 567 => to_unsigned(1168, 12), 568 => to_unsigned(1429, 12), 569 => to_unsigned(3475, 12), 570 => to_unsigned(133, 12), 571 => to_unsigned(1713, 12), 572 => to_unsigned(504, 12), 573 => to_unsigned(1299, 12), 574 => to_unsigned(2083, 12), 575 => to_unsigned(1207, 12), 576 => to_unsigned(531, 12), 577 => to_unsigned(1542, 12), 578 => to_unsigned(2550, 12), 579 => to_unsigned(1363, 12), 580 => to_unsigned(2846, 12), 581 => to_unsigned(1649, 12), 582 => to_unsigned(491, 12), 583 => to_unsigned(92, 12), 584 => to_unsigned(383, 12), 585 => to_unsigned(2951, 12), 586 => to_unsigned(265, 12), 587 => to_unsigned(733, 12), 588 => to_unsigned(2877, 12), 589 => to_unsigned(1630, 12), 590 => to_unsigned(2938, 12), 591 => to_unsigned(634, 12), 592 => to_unsigned(3985, 12), 593 => to_unsigned(903, 12), 594 => to_unsigned(2355, 12), 595 => to_unsigned(689, 12), 596 => to_unsigned(64, 12), 597 => to_unsigned(3926, 12), 598 => to_unsigned(3869, 12), 599 => to_unsigned(823, 12), 600 => to_unsigned(483, 12), 601 => to_unsigned(2932, 12), 602 => to_unsigned(2993, 12), 603 => to_unsigned(693, 12), 604 => to_unsigned(2717, 12), 605 => to_unsigned(1292, 12), 606 => to_unsigned(2648, 12), 607 => to_unsigned(3300, 12), 608 => to_unsigned(2734, 12), 609 => to_unsigned(304, 12), 610 => to_unsigned(942, 12), 611 => to_unsigned(457, 12), 612 => to_unsigned(2270, 12), 613 => to_unsigned(144, 12), 614 => to_unsigned(2170, 12), 615 => to_unsigned(1656, 12), 616 => to_unsigned(3977, 12), 617 => to_unsigned(3064, 12), 618 => to_unsigned(348, 12), 619 => to_unsigned(478, 12), 620 => to_unsigned(1556, 12), 621 => to_unsigned(3168, 12), 622 => to_unsigned(1551, 12), 623 => to_unsigned(2034, 12), 624 => to_unsigned(4006, 12), 625 => to_unsigned(1644, 12), 626 => to_unsigned(1804, 12), 627 => to_unsigned(1138, 12), 628 => to_unsigned(1615, 12), 629 => to_unsigned(3723, 12), 630 => to_unsigned(1867, 12), 631 => to_unsigned(3229, 12), 632 => to_unsigned(1683, 12), 633 => to_unsigned(3175, 12), 634 => to_unsigned(2394, 12), 635 => to_unsigned(2058, 12), 636 => to_unsigned(572, 12), 637 => to_unsigned(3050, 12), 638 => to_unsigned(2290, 12), 639 => to_unsigned(2785, 12), 640 => to_unsigned(2279, 12), 641 => to_unsigned(2524, 12), 642 => to_unsigned(1728, 12), 643 => to_unsigned(3917, 12), 644 => to_unsigned(458, 12), 645 => to_unsigned(307, 12), 646 => to_unsigned(279, 12), 647 => to_unsigned(3811, 12), 648 => to_unsigned(1749, 12), 649 => to_unsigned(1130, 12), 650 => to_unsigned(3962, 12), 651 => to_unsigned(509, 12), 652 => to_unsigned(3456, 12), 653 => to_unsigned(2440, 12), 654 => to_unsigned(3622, 12), 655 => to_unsigned(3195, 12), 656 => to_unsigned(1887, 12), 657 => to_unsigned(3739, 12), 658 => to_unsigned(2272, 12), 659 => to_unsigned(2141, 12), 660 => to_unsigned(3245, 12), 661 => to_unsigned(2163, 12), 662 => to_unsigned(2061, 12), 663 => to_unsigned(3287, 12), 664 => to_unsigned(3737, 12), 665 => to_unsigned(3205, 12), 666 => to_unsigned(2184, 12), 667 => to_unsigned(1554, 12), 668 => to_unsigned(2761, 12), 669 => to_unsigned(1062, 12), 670 => to_unsigned(3570, 12), 671 => to_unsigned(2863, 12), 672 => to_unsigned(1597, 12), 673 => to_unsigned(315, 12), 674 => to_unsigned(1442, 12), 675 => to_unsigned(2219, 12), 676 => to_unsigned(20, 12), 677 => to_unsigned(755, 12), 678 => to_unsigned(2083, 12), 679 => to_unsigned(42, 12), 680 => to_unsigned(30, 12), 681 => to_unsigned(3299, 12), 682 => to_unsigned(1749, 12), 683 => to_unsigned(3183, 12), 684 => to_unsigned(2492, 12), 685 => to_unsigned(3323, 12), 686 => to_unsigned(293, 12), 687 => to_unsigned(563, 12), 688 => to_unsigned(279, 12), 689 => to_unsigned(2101, 12), 690 => to_unsigned(224, 12), 691 => to_unsigned(2977, 12), 692 => to_unsigned(3510, 12), 693 => to_unsigned(3520, 12), 694 => to_unsigned(3188, 12), 695 => to_unsigned(57, 12), 696 => to_unsigned(3732, 12), 697 => to_unsigned(3027, 12), 698 => to_unsigned(3023, 12), 699 => to_unsigned(1233, 12), 700 => to_unsigned(3258, 12), 701 => to_unsigned(2165, 12), 702 => to_unsigned(3315, 12), 703 => to_unsigned(2393, 12), 704 => to_unsigned(79, 12), 705 => to_unsigned(2756, 12), 706 => to_unsigned(1160, 12), 707 => to_unsigned(1589, 12), 708 => to_unsigned(3543, 12), 709 => to_unsigned(642, 12), 710 => to_unsigned(3749, 12), 711 => to_unsigned(2606, 12), 712 => to_unsigned(3929, 12), 713 => to_unsigned(172, 12), 714 => to_unsigned(50, 12), 715 => to_unsigned(1189, 12), 716 => to_unsigned(191, 12), 717 => to_unsigned(726, 12), 718 => to_unsigned(1750, 12), 719 => to_unsigned(181, 12), 720 => to_unsigned(1179, 12), 721 => to_unsigned(1667, 12), 722 => to_unsigned(2503, 12), 723 => to_unsigned(3210, 12), 724 => to_unsigned(2385, 12), 725 => to_unsigned(485, 12), 726 => to_unsigned(262, 12), 727 => to_unsigned(2599, 12), 728 => to_unsigned(1589, 12), 729 => to_unsigned(3968, 12), 730 => to_unsigned(3971, 12), 731 => to_unsigned(3699, 12), 732 => to_unsigned(655, 12), 733 => to_unsigned(3966, 12), 734 => to_unsigned(492, 12), 735 => to_unsigned(592, 12), 736 => to_unsigned(1743, 12), 737 => to_unsigned(3200, 12), 738 => to_unsigned(288, 12), 739 => to_unsigned(3584, 12), 740 => to_unsigned(2699, 12), 741 => to_unsigned(187, 12), 742 => to_unsigned(1496, 12), 743 => to_unsigned(2843, 12), 744 => to_unsigned(2353, 12), 745 => to_unsigned(435, 12), 746 => to_unsigned(17, 12), 747 => to_unsigned(3294, 12), 748 => to_unsigned(1875, 12), 749 => to_unsigned(1708, 12), 750 => to_unsigned(987, 12), 751 => to_unsigned(2421, 12), 752 => to_unsigned(844, 12), 753 => to_unsigned(1738, 12), 754 => to_unsigned(3017, 12), 755 => to_unsigned(1161, 12), 756 => to_unsigned(1261, 12), 757 => to_unsigned(3196, 12), 758 => to_unsigned(3812, 12), 759 => to_unsigned(375, 12), 760 => to_unsigned(2427, 12), 761 => to_unsigned(2713, 12), 762 => to_unsigned(3484, 12), 763 => to_unsigned(2259, 12), 764 => to_unsigned(963, 12), 765 => to_unsigned(2655, 12), 766 => to_unsigned(2646, 12), 767 => to_unsigned(1005, 12), 768 => to_unsigned(861, 12), 769 => to_unsigned(3040, 12), 770 => to_unsigned(864, 12), 771 => to_unsigned(3110, 12), 772 => to_unsigned(541, 12), 773 => to_unsigned(1074, 12), 774 => to_unsigned(1135, 12), 775 => to_unsigned(3742, 12), 776 => to_unsigned(2665, 12), 777 => to_unsigned(526, 12), 778 => to_unsigned(2407, 12), 779 => to_unsigned(2085, 12), 780 => to_unsigned(132, 12), 781 => to_unsigned(3689, 12), 782 => to_unsigned(3643, 12), 783 => to_unsigned(2068, 12), 784 => to_unsigned(1175, 12), 785 => to_unsigned(2832, 12), 786 => to_unsigned(1332, 12), 787 => to_unsigned(1558, 12), 788 => to_unsigned(518, 12), 789 => to_unsigned(1560, 12), 790 => to_unsigned(3355, 12), 791 => to_unsigned(2391, 12), 792 => to_unsigned(4087, 12), 793 => to_unsigned(2858, 12), 794 => to_unsigned(1414, 12), 795 => to_unsigned(669, 12), 796 => to_unsigned(3717, 12), 797 => to_unsigned(3536, 12), 798 => to_unsigned(1133, 12), 799 => to_unsigned(3399, 12), 800 => to_unsigned(1024, 12), 801 => to_unsigned(698, 12), 802 => to_unsigned(3402, 12), 803 => to_unsigned(3884, 12), 804 => to_unsigned(2942, 12), 805 => to_unsigned(71, 12), 806 => to_unsigned(1453, 12), 807 => to_unsigned(1443, 12), 808 => to_unsigned(3841, 12), 809 => to_unsigned(392, 12), 810 => to_unsigned(2331, 12), 811 => to_unsigned(3947, 12), 812 => to_unsigned(1565, 12), 813 => to_unsigned(3557, 12), 814 => to_unsigned(3878, 12), 815 => to_unsigned(1039, 12), 816 => to_unsigned(1067, 12), 817 => to_unsigned(811, 12), 818 => to_unsigned(571, 12), 819 => to_unsigned(2572, 12), 820 => to_unsigned(268, 12), 821 => to_unsigned(1962, 12), 822 => to_unsigned(1812, 12), 823 => to_unsigned(1238, 12), 824 => to_unsigned(423, 12), 825 => to_unsigned(2528, 12), 826 => to_unsigned(3248, 12), 827 => to_unsigned(804, 12), 828 => to_unsigned(1575, 12), 829 => to_unsigned(1731, 12), 830 => to_unsigned(54, 12), 831 => to_unsigned(3202, 12), 832 => to_unsigned(1930, 12), 833 => to_unsigned(2197, 12), 834 => to_unsigned(2004, 12), 835 => to_unsigned(3543, 12), 836 => to_unsigned(2853, 12), 837 => to_unsigned(761, 12), 838 => to_unsigned(1436, 12), 839 => to_unsigned(1694, 12), 840 => to_unsigned(2339, 12), 841 => to_unsigned(2803, 12), 842 => to_unsigned(532, 12), 843 => to_unsigned(753, 12), 844 => to_unsigned(614, 12), 845 => to_unsigned(1775, 12), 846 => to_unsigned(1203, 12), 847 => to_unsigned(1872, 12), 848 => to_unsigned(728, 12), 849 => to_unsigned(287, 12), 850 => to_unsigned(2816, 12), 851 => to_unsigned(1040, 12), 852 => to_unsigned(790, 12), 853 => to_unsigned(43, 12), 854 => to_unsigned(990, 12), 855 => to_unsigned(3154, 12), 856 => to_unsigned(4091, 12), 857 => to_unsigned(3442, 12), 858 => to_unsigned(3966, 12), 859 => to_unsigned(3870, 12), 860 => to_unsigned(633, 12), 861 => to_unsigned(3905, 12), 862 => to_unsigned(2086, 12), 863 => to_unsigned(1830, 12), 864 => to_unsigned(1107, 12), 865 => to_unsigned(2410, 12), 866 => to_unsigned(1333, 12), 867 => to_unsigned(1691, 12), 868 => to_unsigned(443, 12), 869 => to_unsigned(1294, 12), 870 => to_unsigned(1234, 12), 871 => to_unsigned(3821, 12), 872 => to_unsigned(1326, 12), 873 => to_unsigned(2804, 12), 874 => to_unsigned(3441, 12), 875 => to_unsigned(3637, 12), 876 => to_unsigned(3197, 12), 877 => to_unsigned(1713, 12), 878 => to_unsigned(465, 12), 879 => to_unsigned(17, 12), 880 => to_unsigned(917, 12), 881 => to_unsigned(709, 12), 882 => to_unsigned(17, 12), 883 => to_unsigned(1923, 12), 884 => to_unsigned(1827, 12), 885 => to_unsigned(4023, 12), 886 => to_unsigned(910, 12), 887 => to_unsigned(371, 12), 888 => to_unsigned(2604, 12), 889 => to_unsigned(804, 12), 890 => to_unsigned(1028, 12), 891 => to_unsigned(834, 12), 892 => to_unsigned(3192, 12), 893 => to_unsigned(1131, 12), 894 => to_unsigned(2603, 12), 895 => to_unsigned(2557, 12), 896 => to_unsigned(70, 12), 897 => to_unsigned(1570, 12), 898 => to_unsigned(1501, 12), 899 => to_unsigned(3615, 12), 900 => to_unsigned(2370, 12), 901 => to_unsigned(2773, 12), 902 => to_unsigned(1385, 12), 903 => to_unsigned(2042, 12), 904 => to_unsigned(2146, 12), 905 => to_unsigned(169, 12), 906 => to_unsigned(3364, 12), 907 => to_unsigned(417, 12), 908 => to_unsigned(57, 12), 909 => to_unsigned(3777, 12), 910 => to_unsigned(2098, 12), 911 => to_unsigned(3096, 12), 912 => to_unsigned(2810, 12), 913 => to_unsigned(2875, 12), 914 => to_unsigned(1892, 12), 915 => to_unsigned(1792, 12), 916 => to_unsigned(3523, 12), 917 => to_unsigned(1634, 12), 918 => to_unsigned(1344, 12), 919 => to_unsigned(646, 12), 920 => to_unsigned(1860, 12), 921 => to_unsigned(153, 12), 922 => to_unsigned(1054, 12), 923 => to_unsigned(2327, 12), 924 => to_unsigned(2541, 12), 925 => to_unsigned(337, 12), 926 => to_unsigned(1374, 12), 927 => to_unsigned(4003, 12), 928 => to_unsigned(826, 12), 929 => to_unsigned(1994, 12), 930 => to_unsigned(1319, 12), 931 => to_unsigned(1150, 12), 932 => to_unsigned(1246, 12), 933 => to_unsigned(999, 12), 934 => to_unsigned(150, 12), 935 => to_unsigned(2324, 12), 936 => to_unsigned(3510, 12), 937 => to_unsigned(4082, 12), 938 => to_unsigned(1692, 12), 939 => to_unsigned(429, 12), 940 => to_unsigned(2747, 12), 941 => to_unsigned(1598, 12), 942 => to_unsigned(3045, 12), 943 => to_unsigned(3248, 12), 944 => to_unsigned(1509, 12), 945 => to_unsigned(2883, 12), 946 => to_unsigned(2419, 12), 947 => to_unsigned(3193, 12), 948 => to_unsigned(1002, 12), 949 => to_unsigned(3829, 12), 950 => to_unsigned(2831, 12), 951 => to_unsigned(3156, 12), 952 => to_unsigned(1031, 12), 953 => to_unsigned(1137, 12), 954 => to_unsigned(474, 12), 955 => to_unsigned(4046, 12), 956 => to_unsigned(1513, 12), 957 => to_unsigned(1176, 12), 958 => to_unsigned(242, 12), 959 => to_unsigned(2120, 12), 960 => to_unsigned(2166, 12), 961 => to_unsigned(949, 12), 962 => to_unsigned(2064, 12), 963 => to_unsigned(186, 12), 964 => to_unsigned(639, 12), 965 => to_unsigned(1224, 12), 966 => to_unsigned(2236, 12), 967 => to_unsigned(2764, 12), 968 => to_unsigned(35, 12), 969 => to_unsigned(2981, 12), 970 => to_unsigned(1609, 12), 971 => to_unsigned(1435, 12), 972 => to_unsigned(2753, 12), 973 => to_unsigned(3388, 12), 974 => to_unsigned(2701, 12), 975 => to_unsigned(2334, 12), 976 => to_unsigned(669, 12), 977 => to_unsigned(2236, 12), 978 => to_unsigned(1814, 12), 979 => to_unsigned(118, 12), 980 => to_unsigned(1726, 12), 981 => to_unsigned(831, 12), 982 => to_unsigned(940, 12), 983 => to_unsigned(576, 12), 984 => to_unsigned(1768, 12), 985 => to_unsigned(2677, 12), 986 => to_unsigned(3352, 12), 987 => to_unsigned(2855, 12), 988 => to_unsigned(2858, 12), 989 => to_unsigned(2992, 12), 990 => to_unsigned(3306, 12), 991 => to_unsigned(2992, 12), 992 => to_unsigned(2542, 12), 993 => to_unsigned(1634, 12), 994 => to_unsigned(2983, 12), 995 => to_unsigned(274, 12), 996 => to_unsigned(3550, 12), 997 => to_unsigned(2317, 12), 998 => to_unsigned(885, 12), 999 => to_unsigned(3709, 12), 1000 => to_unsigned(3099, 12), 1001 => to_unsigned(2227, 12), 1002 => to_unsigned(2712, 12), 1003 => to_unsigned(2915, 12), 1004 => to_unsigned(2583, 12), 1005 => to_unsigned(2418, 12), 1006 => to_unsigned(3384, 12), 1007 => to_unsigned(471, 12), 1008 => to_unsigned(3302, 12), 1009 => to_unsigned(2194, 12), 1010 => to_unsigned(3749, 12), 1011 => to_unsigned(785, 12), 1012 => to_unsigned(3512, 12), 1013 => to_unsigned(1452, 12), 1014 => to_unsigned(1529, 12), 1015 => to_unsigned(1678, 12), 1016 => to_unsigned(2930, 12), 1017 => to_unsigned(3707, 12), 1018 => to_unsigned(1336, 12), 1019 => to_unsigned(2872, 12), 1020 => to_unsigned(3816, 12), 1021 => to_unsigned(2621, 12), 1022 => to_unsigned(3271, 12), 1023 => to_unsigned(2915, 12), 1024 => to_unsigned(3528, 12), 1025 => to_unsigned(3462, 12), 1026 => to_unsigned(1062, 12), 1027 => to_unsigned(1591, 12), 1028 => to_unsigned(3721, 12), 1029 => to_unsigned(683, 12), 1030 => to_unsigned(2822, 12), 1031 => to_unsigned(3999, 12), 1032 => to_unsigned(2878, 12), 1033 => to_unsigned(1734, 12), 1034 => to_unsigned(915, 12), 1035 => to_unsigned(1068, 12), 1036 => to_unsigned(1579, 12), 1037 => to_unsigned(311, 12), 1038 => to_unsigned(3486, 12), 1039 => to_unsigned(1775, 12), 1040 => to_unsigned(3710, 12), 1041 => to_unsigned(518, 12), 1042 => to_unsigned(241, 12), 1043 => to_unsigned(1670, 12), 1044 => to_unsigned(400, 12), 1045 => to_unsigned(3430, 12), 1046 => to_unsigned(2494, 12), 1047 => to_unsigned(1203, 12), 1048 => to_unsigned(1227, 12), 1049 => to_unsigned(2880, 12), 1050 => to_unsigned(1277, 12), 1051 => to_unsigned(3459, 12), 1052 => to_unsigned(1754, 12), 1053 => to_unsigned(1549, 12), 1054 => to_unsigned(79, 12), 1055 => to_unsigned(510, 12), 1056 => to_unsigned(1054, 12), 1057 => to_unsigned(3919, 12), 1058 => to_unsigned(3569, 12), 1059 => to_unsigned(3596, 12), 1060 => to_unsigned(2687, 12), 1061 => to_unsigned(2397, 12), 1062 => to_unsigned(2602, 12), 1063 => to_unsigned(2737, 12), 1064 => to_unsigned(2318, 12), 1065 => to_unsigned(387, 12), 1066 => to_unsigned(3130, 12), 1067 => to_unsigned(2353, 12), 1068 => to_unsigned(138, 12), 1069 => to_unsigned(2617, 12), 1070 => to_unsigned(1208, 12), 1071 => to_unsigned(1786, 12), 1072 => to_unsigned(3024, 12), 1073 => to_unsigned(1091, 12), 1074 => to_unsigned(1037, 12), 1075 => to_unsigned(3207, 12), 1076 => to_unsigned(755, 12), 1077 => to_unsigned(2002, 12), 1078 => to_unsigned(3951, 12), 1079 => to_unsigned(3815, 12), 1080 => to_unsigned(1552, 12), 1081 => to_unsigned(3613, 12), 1082 => to_unsigned(1094, 12), 1083 => to_unsigned(2529, 12), 1084 => to_unsigned(1589, 12), 1085 => to_unsigned(862, 12), 1086 => to_unsigned(3115, 12), 1087 => to_unsigned(2177, 12), 1088 => to_unsigned(2440, 12), 1089 => to_unsigned(3993, 12), 1090 => to_unsigned(3518, 12), 1091 => to_unsigned(1511, 12), 1092 => to_unsigned(3299, 12), 1093 => to_unsigned(59, 12), 1094 => to_unsigned(645, 12), 1095 => to_unsigned(2710, 12), 1096 => to_unsigned(3323, 12), 1097 => to_unsigned(1843, 12), 1098 => to_unsigned(2812, 12), 1099 => to_unsigned(1413, 12), 1100 => to_unsigned(882, 12), 1101 => to_unsigned(1742, 12), 1102 => to_unsigned(2916, 12), 1103 => to_unsigned(917, 12), 1104 => to_unsigned(3348, 12), 1105 => to_unsigned(2949, 12), 1106 => to_unsigned(3454, 12), 1107 => to_unsigned(1875, 12), 1108 => to_unsigned(2830, 12), 1109 => to_unsigned(2606, 12), 1110 => to_unsigned(2123, 12), 1111 => to_unsigned(46, 12), 1112 => to_unsigned(135, 12), 1113 => to_unsigned(1669, 12), 1114 => to_unsigned(3986, 12), 1115 => to_unsigned(2836, 12), 1116 => to_unsigned(3464, 12), 1117 => to_unsigned(1297, 12), 1118 => to_unsigned(825, 12), 1119 => to_unsigned(291, 12), 1120 => to_unsigned(437, 12), 1121 => to_unsigned(1020, 12), 1122 => to_unsigned(863, 12), 1123 => to_unsigned(864, 12), 1124 => to_unsigned(3090, 12), 1125 => to_unsigned(1120, 12), 1126 => to_unsigned(2497, 12), 1127 => to_unsigned(3812, 12), 1128 => to_unsigned(3711, 12), 1129 => to_unsigned(2612, 12), 1130 => to_unsigned(187, 12), 1131 => to_unsigned(2872, 12), 1132 => to_unsigned(3729, 12), 1133 => to_unsigned(2343, 12), 1134 => to_unsigned(979, 12), 1135 => to_unsigned(3871, 12), 1136 => to_unsigned(682, 12), 1137 => to_unsigned(2951, 12), 1138 => to_unsigned(862, 12), 1139 => to_unsigned(1348, 12), 1140 => to_unsigned(2114, 12), 1141 => to_unsigned(3899, 12), 1142 => to_unsigned(4033, 12), 1143 => to_unsigned(38, 12), 1144 => to_unsigned(128, 12), 1145 => to_unsigned(3574, 12), 1146 => to_unsigned(3596, 12), 1147 => to_unsigned(1403, 12), 1148 => to_unsigned(1717, 12), 1149 => to_unsigned(942, 12), 1150 => to_unsigned(1313, 12), 1151 => to_unsigned(729, 12), 1152 => to_unsigned(1703, 12), 1153 => to_unsigned(2794, 12), 1154 => to_unsigned(1494, 12), 1155 => to_unsigned(3180, 12), 1156 => to_unsigned(269, 12), 1157 => to_unsigned(3847, 12), 1158 => to_unsigned(3713, 12), 1159 => to_unsigned(3490, 12), 1160 => to_unsigned(2579, 12), 1161 => to_unsigned(2631, 12), 1162 => to_unsigned(2710, 12), 1163 => to_unsigned(2591, 12), 1164 => to_unsigned(3234, 12), 1165 => to_unsigned(3111, 12), 1166 => to_unsigned(2780, 12), 1167 => to_unsigned(649, 12), 1168 => to_unsigned(3166, 12), 1169 => to_unsigned(3975, 12), 1170 => to_unsigned(2327, 12), 1171 => to_unsigned(615, 12), 1172 => to_unsigned(2683, 12), 1173 => to_unsigned(1570, 12), 1174 => to_unsigned(2598, 12), 1175 => to_unsigned(329, 12), 1176 => to_unsigned(1735, 12), 1177 => to_unsigned(100, 12), 1178 => to_unsigned(3863, 12), 1179 => to_unsigned(100, 12), 1180 => to_unsigned(1408, 12), 1181 => to_unsigned(2219, 12), 1182 => to_unsigned(1960, 12), 1183 => to_unsigned(1510, 12), 1184 => to_unsigned(4028, 12), 1185 => to_unsigned(1574, 12), 1186 => to_unsigned(3406, 12), 1187 => to_unsigned(3305, 12), 1188 => to_unsigned(2797, 12), 1189 => to_unsigned(1189, 12), 1190 => to_unsigned(1331, 12), 1191 => to_unsigned(586, 12), 1192 => to_unsigned(2240, 12), 1193 => to_unsigned(2782, 12), 1194 => to_unsigned(1969, 12), 1195 => to_unsigned(3991, 12), 1196 => to_unsigned(1750, 12), 1197 => to_unsigned(3149, 12), 1198 => to_unsigned(2077, 12), 1199 => to_unsigned(3741, 12), 1200 => to_unsigned(1693, 12), 1201 => to_unsigned(626, 12), 1202 => to_unsigned(2885, 12), 1203 => to_unsigned(1595, 12), 1204 => to_unsigned(403, 12), 1205 => to_unsigned(384, 12), 1206 => to_unsigned(2025, 12), 1207 => to_unsigned(897, 12), 1208 => to_unsigned(2799, 12), 1209 => to_unsigned(3285, 12), 1210 => to_unsigned(3619, 12), 1211 => to_unsigned(1879, 12), 1212 => to_unsigned(1260, 12), 1213 => to_unsigned(3438, 12), 1214 => to_unsigned(729, 12), 1215 => to_unsigned(3774, 12), 1216 => to_unsigned(1820, 12), 1217 => to_unsigned(1494, 12), 1218 => to_unsigned(1421, 12), 1219 => to_unsigned(1796, 12), 1220 => to_unsigned(813, 12), 1221 => to_unsigned(1626, 12), 1222 => to_unsigned(872, 12), 1223 => to_unsigned(3615, 12), 1224 => to_unsigned(603, 12), 1225 => to_unsigned(3115, 12), 1226 => to_unsigned(2098, 12), 1227 => to_unsigned(1021, 12), 1228 => to_unsigned(3212, 12), 1229 => to_unsigned(4009, 12), 1230 => to_unsigned(986, 12), 1231 => to_unsigned(206, 12), 1232 => to_unsigned(1978, 12), 1233 => to_unsigned(3516, 12), 1234 => to_unsigned(3327, 12), 1235 => to_unsigned(54, 12), 1236 => to_unsigned(337, 12), 1237 => to_unsigned(1618, 12), 1238 => to_unsigned(3415, 12), 1239 => to_unsigned(774, 12), 1240 => to_unsigned(1340, 12), 1241 => to_unsigned(2333, 12), 1242 => to_unsigned(2364, 12), 1243 => to_unsigned(868, 12), 1244 => to_unsigned(2604, 12), 1245 => to_unsigned(2862, 12), 1246 => to_unsigned(3090, 12), 1247 => to_unsigned(1883, 12), 1248 => to_unsigned(1826, 12), 1249 => to_unsigned(615, 12), 1250 => to_unsigned(1468, 12), 1251 => to_unsigned(2977, 12), 1252 => to_unsigned(2434, 12), 1253 => to_unsigned(327, 12), 1254 => to_unsigned(1241, 12), 1255 => to_unsigned(3776, 12), 1256 => to_unsigned(3550, 12), 1257 => to_unsigned(2204, 12), 1258 => to_unsigned(1810, 12), 1259 => to_unsigned(2012, 12), 1260 => to_unsigned(911, 12), 1261 => to_unsigned(89, 12), 1262 => to_unsigned(3483, 12), 1263 => to_unsigned(349, 12), 1264 => to_unsigned(2715, 12), 1265 => to_unsigned(110, 12), 1266 => to_unsigned(4071, 12), 1267 => to_unsigned(3837, 12), 1268 => to_unsigned(3079, 12), 1269 => to_unsigned(361, 12), 1270 => to_unsigned(2730, 12), 1271 => to_unsigned(804, 12), 1272 => to_unsigned(594, 12), 1273 => to_unsigned(801, 12), 1274 => to_unsigned(1093, 12), 1275 => to_unsigned(1852, 12), 1276 => to_unsigned(3037, 12), 1277 => to_unsigned(2511, 12), 1278 => to_unsigned(2526, 12), 1279 => to_unsigned(718, 12), 1280 => to_unsigned(3143, 12), 1281 => to_unsigned(2385, 12), 1282 => to_unsigned(1158, 12), 1283 => to_unsigned(1768, 12), 1284 => to_unsigned(4062, 12), 1285 => to_unsigned(2048, 12), 1286 => to_unsigned(253, 12), 1287 => to_unsigned(234, 12), 1288 => to_unsigned(2807, 12), 1289 => to_unsigned(1498, 12), 1290 => to_unsigned(2827, 12), 1291 => to_unsigned(1848, 12), 1292 => to_unsigned(1544, 12), 1293 => to_unsigned(732, 12), 1294 => to_unsigned(2686, 12), 1295 => to_unsigned(2867, 12), 1296 => to_unsigned(1271, 12), 1297 => to_unsigned(1617, 12), 1298 => to_unsigned(165, 12), 1299 => to_unsigned(36, 12), 1300 => to_unsigned(4091, 12), 1301 => to_unsigned(3366, 12), 1302 => to_unsigned(1764, 12), 1303 => to_unsigned(2627, 12), 1304 => to_unsigned(3264, 12), 1305 => to_unsigned(1285, 12), 1306 => to_unsigned(917, 12), 1307 => to_unsigned(3380, 12), 1308 => to_unsigned(954, 12), 1309 => to_unsigned(1868, 12), 1310 => to_unsigned(3795, 12), 1311 => to_unsigned(2218, 12), 1312 => to_unsigned(2438, 12), 1313 => to_unsigned(2048, 12), 1314 => to_unsigned(2136, 12), 1315 => to_unsigned(3084, 12), 1316 => to_unsigned(55, 12), 1317 => to_unsigned(4058, 12), 1318 => to_unsigned(319, 12), 1319 => to_unsigned(1595, 12), 1320 => to_unsigned(3444, 12), 1321 => to_unsigned(1738, 12), 1322 => to_unsigned(2594, 12), 1323 => to_unsigned(86, 12), 1324 => to_unsigned(3762, 12), 1325 => to_unsigned(313, 12), 1326 => to_unsigned(1614, 12), 1327 => to_unsigned(3872, 12), 1328 => to_unsigned(3291, 12), 1329 => to_unsigned(3007, 12), 1330 => to_unsigned(2840, 12), 1331 => to_unsigned(3871, 12), 1332 => to_unsigned(1100, 12), 1333 => to_unsigned(323, 12), 1334 => to_unsigned(858, 12), 1335 => to_unsigned(2096, 12), 1336 => to_unsigned(2391, 12), 1337 => to_unsigned(826, 12), 1338 => to_unsigned(3520, 12), 1339 => to_unsigned(2826, 12), 1340 => to_unsigned(1309, 12), 1341 => to_unsigned(673, 12), 1342 => to_unsigned(1511, 12), 1343 => to_unsigned(923, 12), 1344 => to_unsigned(533, 12), 1345 => to_unsigned(3422, 12), 1346 => to_unsigned(1871, 12), 1347 => to_unsigned(3961, 12), 1348 => to_unsigned(497, 12), 1349 => to_unsigned(4073, 12), 1350 => to_unsigned(1224, 12), 1351 => to_unsigned(1511, 12), 1352 => to_unsigned(2199, 12), 1353 => to_unsigned(3491, 12), 1354 => to_unsigned(2358, 12), 1355 => to_unsigned(247, 12), 1356 => to_unsigned(435, 12), 1357 => to_unsigned(946, 12), 1358 => to_unsigned(1304, 12), 1359 => to_unsigned(3354, 12), 1360 => to_unsigned(3612, 12), 1361 => to_unsigned(78, 12), 1362 => to_unsigned(4046, 12), 1363 => to_unsigned(123, 12), 1364 => to_unsigned(1492, 12), 1365 => to_unsigned(942, 12), 1366 => to_unsigned(3878, 12), 1367 => to_unsigned(1475, 12), 1368 => to_unsigned(911, 12), 1369 => to_unsigned(2327, 12), 1370 => to_unsigned(484, 12), 1371 => to_unsigned(2302, 12), 1372 => to_unsigned(1213, 12), 1373 => to_unsigned(1240, 12), 1374 => to_unsigned(977, 12), 1375 => to_unsigned(2910, 12), 1376 => to_unsigned(4049, 12), 1377 => to_unsigned(1169, 12), 1378 => to_unsigned(2362, 12), 1379 => to_unsigned(2726, 12), 1380 => to_unsigned(1459, 12), 1381 => to_unsigned(80, 12), 1382 => to_unsigned(47, 12), 1383 => to_unsigned(1802, 12), 1384 => to_unsigned(3461, 12), 1385 => to_unsigned(1218, 12), 1386 => to_unsigned(782, 12), 1387 => to_unsigned(2789, 12), 1388 => to_unsigned(1332, 12), 1389 => to_unsigned(1472, 12), 1390 => to_unsigned(1565, 12), 1391 => to_unsigned(1940, 12), 1392 => to_unsigned(3013, 12), 1393 => to_unsigned(2307, 12), 1394 => to_unsigned(1012, 12), 1395 => to_unsigned(4042, 12), 1396 => to_unsigned(462, 12), 1397 => to_unsigned(1285, 12), 1398 => to_unsigned(2454, 12), 1399 => to_unsigned(1091, 12), 1400 => to_unsigned(2828, 12), 1401 => to_unsigned(876, 12), 1402 => to_unsigned(1536, 12), 1403 => to_unsigned(2208, 12), 1404 => to_unsigned(2086, 12), 1405 => to_unsigned(1660, 12), 1406 => to_unsigned(2244, 12), 1407 => to_unsigned(3032, 12), 1408 => to_unsigned(3806, 12), 1409 => to_unsigned(2932, 12), 1410 => to_unsigned(2344, 12), 1411 => to_unsigned(126, 12), 1412 => to_unsigned(2116, 12), 1413 => to_unsigned(906, 12), 1414 => to_unsigned(3804, 12), 1415 => to_unsigned(2845, 12), 1416 => to_unsigned(656, 12), 1417 => to_unsigned(468, 12), 1418 => to_unsigned(3088, 12), 1419 => to_unsigned(459, 12), 1420 => to_unsigned(3924, 12), 1421 => to_unsigned(1161, 12), 1422 => to_unsigned(1685, 12), 1423 => to_unsigned(2686, 12), 1424 => to_unsigned(3154, 12), 1425 => to_unsigned(2126, 12), 1426 => to_unsigned(3447, 12), 1427 => to_unsigned(4023, 12), 1428 => to_unsigned(3099, 12), 1429 => to_unsigned(639, 12), 1430 => to_unsigned(1449, 12), 1431 => to_unsigned(3571, 12), 1432 => to_unsigned(1481, 12), 1433 => to_unsigned(1315, 12), 1434 => to_unsigned(4031, 12), 1435 => to_unsigned(1527, 12), 1436 => to_unsigned(2131, 12), 1437 => to_unsigned(1850, 12), 1438 => to_unsigned(10, 12), 1439 => to_unsigned(1589, 12), 1440 => to_unsigned(3776, 12), 1441 => to_unsigned(2710, 12), 1442 => to_unsigned(2022, 12), 1443 => to_unsigned(2475, 12), 1444 => to_unsigned(3966, 12), 1445 => to_unsigned(3016, 12), 1446 => to_unsigned(203, 12), 1447 => to_unsigned(1117, 12), 1448 => to_unsigned(3740, 12), 1449 => to_unsigned(3764, 12), 1450 => to_unsigned(128, 12), 1451 => to_unsigned(4033, 12), 1452 => to_unsigned(81, 12), 1453 => to_unsigned(3084, 12), 1454 => to_unsigned(1068, 12), 1455 => to_unsigned(4063, 12), 1456 => to_unsigned(3763, 12), 1457 => to_unsigned(739, 12), 1458 => to_unsigned(3945, 12), 1459 => to_unsigned(266, 12), 1460 => to_unsigned(3833, 12), 1461 => to_unsigned(3772, 12), 1462 => to_unsigned(1641, 12), 1463 => to_unsigned(1196, 12), 1464 => to_unsigned(1683, 12), 1465 => to_unsigned(1085, 12), 1466 => to_unsigned(1458, 12), 1467 => to_unsigned(3514, 12), 1468 => to_unsigned(3701, 12), 1469 => to_unsigned(1852, 12), 1470 => to_unsigned(2938, 12), 1471 => to_unsigned(3180, 12), 1472 => to_unsigned(2451, 12), 1473 => to_unsigned(1766, 12), 1474 => to_unsigned(2249, 12), 1475 => to_unsigned(3853, 12), 1476 => to_unsigned(2638, 12), 1477 => to_unsigned(2885, 12), 1478 => to_unsigned(1267, 12), 1479 => to_unsigned(1517, 12), 1480 => to_unsigned(2291, 12), 1481 => to_unsigned(1265, 12), 1482 => to_unsigned(2234, 12), 1483 => to_unsigned(3700, 12), 1484 => to_unsigned(3795, 12), 1485 => to_unsigned(2731, 12), 1486 => to_unsigned(1148, 12), 1487 => to_unsigned(3169, 12), 1488 => to_unsigned(804, 12), 1489 => to_unsigned(1388, 12), 1490 => to_unsigned(3811, 12), 1491 => to_unsigned(2932, 12), 1492 => to_unsigned(670, 12), 1493 => to_unsigned(3256, 12), 1494 => to_unsigned(3320, 12), 1495 => to_unsigned(1536, 12), 1496 => to_unsigned(2973, 12), 1497 => to_unsigned(2811, 12), 1498 => to_unsigned(3443, 12), 1499 => to_unsigned(3689, 12), 1500 => to_unsigned(353, 12), 1501 => to_unsigned(2571, 12), 1502 => to_unsigned(2865, 12), 1503 => to_unsigned(3626, 12), 1504 => to_unsigned(3333, 12), 1505 => to_unsigned(393, 12), 1506 => to_unsigned(2459, 12), 1507 => to_unsigned(3758, 12), 1508 => to_unsigned(2219, 12), 1509 => to_unsigned(1551, 12), 1510 => to_unsigned(3519, 12), 1511 => to_unsigned(1955, 12), 1512 => to_unsigned(1034, 12), 1513 => to_unsigned(3975, 12), 1514 => to_unsigned(3598, 12), 1515 => to_unsigned(2640, 12), 1516 => to_unsigned(2211, 12), 1517 => to_unsigned(1162, 12), 1518 => to_unsigned(492, 12), 1519 => to_unsigned(3206, 12), 1520 => to_unsigned(2587, 12), 1521 => to_unsigned(2801, 12), 1522 => to_unsigned(2287, 12), 1523 => to_unsigned(2806, 12), 1524 => to_unsigned(1942, 12), 1525 => to_unsigned(1247, 12), 1526 => to_unsigned(1074, 12), 1527 => to_unsigned(140, 12), 1528 => to_unsigned(1151, 12), 1529 => to_unsigned(3513, 12), 1530 => to_unsigned(3362, 12), 1531 => to_unsigned(3928, 12), 1532 => to_unsigned(2033, 12), 1533 => to_unsigned(298, 12), 1534 => to_unsigned(3534, 12), 1535 => to_unsigned(3568, 12), 1536 => to_unsigned(1744, 12), 1537 => to_unsigned(1646, 12), 1538 => to_unsigned(689, 12), 1539 => to_unsigned(1684, 12), 1540 => to_unsigned(665, 12), 1541 => to_unsigned(784, 12), 1542 => to_unsigned(242, 12), 1543 => to_unsigned(4070, 12), 1544 => to_unsigned(2222, 12), 1545 => to_unsigned(704, 12), 1546 => to_unsigned(497, 12), 1547 => to_unsigned(2901, 12), 1548 => to_unsigned(3432, 12), 1549 => to_unsigned(1436, 12), 1550 => to_unsigned(453, 12), 1551 => to_unsigned(3424, 12), 1552 => to_unsigned(844, 12), 1553 => to_unsigned(2524, 12), 1554 => to_unsigned(1226, 12), 1555 => to_unsigned(1272, 12), 1556 => to_unsigned(4042, 12), 1557 => to_unsigned(1275, 12), 1558 => to_unsigned(1338, 12), 1559 => to_unsigned(3994, 12), 1560 => to_unsigned(1463, 12), 1561 => to_unsigned(132, 12), 1562 => to_unsigned(4084, 12), 1563 => to_unsigned(2811, 12), 1564 => to_unsigned(3781, 12), 1565 => to_unsigned(3156, 12), 1566 => to_unsigned(1220, 12), 1567 => to_unsigned(530, 12), 1568 => to_unsigned(3484, 12), 1569 => to_unsigned(3176, 12), 1570 => to_unsigned(955, 12), 1571 => to_unsigned(3932, 12), 1572 => to_unsigned(1345, 12), 1573 => to_unsigned(1538, 12), 1574 => to_unsigned(2653, 12), 1575 => to_unsigned(175, 12), 1576 => to_unsigned(1386, 12), 1577 => to_unsigned(3392, 12), 1578 => to_unsigned(2375, 12), 1579 => to_unsigned(1393, 12), 1580 => to_unsigned(1221, 12), 1581 => to_unsigned(411, 12), 1582 => to_unsigned(962, 12), 1583 => to_unsigned(3008, 12), 1584 => to_unsigned(1412, 12), 1585 => to_unsigned(843, 12), 1586 => to_unsigned(1706, 12), 1587 => to_unsigned(1439, 12), 1588 => to_unsigned(1500, 12), 1589 => to_unsigned(1108, 12), 1590 => to_unsigned(3240, 12), 1591 => to_unsigned(773, 12), 1592 => to_unsigned(3172, 12), 1593 => to_unsigned(2499, 12), 1594 => to_unsigned(535, 12), 1595 => to_unsigned(157, 12), 1596 => to_unsigned(1908, 12), 1597 => to_unsigned(3933, 12), 1598 => to_unsigned(290, 12), 1599 => to_unsigned(1751, 12), 1600 => to_unsigned(2237, 12), 1601 => to_unsigned(38, 12), 1602 => to_unsigned(3507, 12), 1603 => to_unsigned(3563, 12), 1604 => to_unsigned(1591, 12), 1605 => to_unsigned(1632, 12), 1606 => to_unsigned(3399, 12), 1607 => to_unsigned(3152, 12), 1608 => to_unsigned(3432, 12), 1609 => to_unsigned(793, 12), 1610 => to_unsigned(1454, 12), 1611 => to_unsigned(2353, 12), 1612 => to_unsigned(176, 12), 1613 => to_unsigned(3982, 12), 1614 => to_unsigned(68, 12), 1615 => to_unsigned(3006, 12), 1616 => to_unsigned(2180, 12), 1617 => to_unsigned(3227, 12), 1618 => to_unsigned(2301, 12), 1619 => to_unsigned(2988, 12), 1620 => to_unsigned(3140, 12), 1621 => to_unsigned(1158, 12), 1622 => to_unsigned(938, 12), 1623 => to_unsigned(1531, 12), 1624 => to_unsigned(152, 12), 1625 => to_unsigned(3384, 12), 1626 => to_unsigned(1332, 12), 1627 => to_unsigned(2607, 12), 1628 => to_unsigned(1840, 12), 1629 => to_unsigned(887, 12), 1630 => to_unsigned(3231, 12), 1631 => to_unsigned(3608, 12), 1632 => to_unsigned(2260, 12), 1633 => to_unsigned(1775, 12), 1634 => to_unsigned(1517, 12), 1635 => to_unsigned(3174, 12), 1636 => to_unsigned(438, 12), 1637 => to_unsigned(2180, 12), 1638 => to_unsigned(2470, 12), 1639 => to_unsigned(3048, 12), 1640 => to_unsigned(3514, 12), 1641 => to_unsigned(315, 12), 1642 => to_unsigned(1437, 12), 1643 => to_unsigned(1146, 12), 1644 => to_unsigned(3134, 12), 1645 => to_unsigned(3684, 12), 1646 => to_unsigned(1411, 12), 1647 => to_unsigned(1922, 12), 1648 => to_unsigned(2945, 12), 1649 => to_unsigned(178, 12), 1650 => to_unsigned(1422, 12), 1651 => to_unsigned(3063, 12), 1652 => to_unsigned(1254, 12), 1653 => to_unsigned(2205, 12), 1654 => to_unsigned(4069, 12), 1655 => to_unsigned(741, 12), 1656 => to_unsigned(3517, 12), 1657 => to_unsigned(1688, 12), 1658 => to_unsigned(1687, 12), 1659 => to_unsigned(472, 12), 1660 => to_unsigned(3880, 12), 1661 => to_unsigned(1924, 12), 1662 => to_unsigned(3982, 12), 1663 => to_unsigned(2368, 12), 1664 => to_unsigned(3867, 12), 1665 => to_unsigned(3202, 12), 1666 => to_unsigned(2986, 12), 1667 => to_unsigned(3700, 12), 1668 => to_unsigned(1499, 12), 1669 => to_unsigned(1359, 12), 1670 => to_unsigned(2519, 12), 1671 => to_unsigned(915, 12), 1672 => to_unsigned(3267, 12), 1673 => to_unsigned(1897, 12), 1674 => to_unsigned(2456, 12), 1675 => to_unsigned(3433, 12), 1676 => to_unsigned(3190, 12), 1677 => to_unsigned(4050, 12), 1678 => to_unsigned(38, 12), 1679 => to_unsigned(1388, 12), 1680 => to_unsigned(2443, 12), 1681 => to_unsigned(128, 12), 1682 => to_unsigned(2097, 12), 1683 => to_unsigned(2413, 12), 1684 => to_unsigned(3185, 12), 1685 => to_unsigned(1824, 12), 1686 => to_unsigned(478, 12), 1687 => to_unsigned(901, 12), 1688 => to_unsigned(3197, 12), 1689 => to_unsigned(1266, 12), 1690 => to_unsigned(3581, 12), 1691 => to_unsigned(1206, 12), 1692 => to_unsigned(2048, 12), 1693 => to_unsigned(186, 12), 1694 => to_unsigned(27, 12), 1695 => to_unsigned(3635, 12), 1696 => to_unsigned(3562, 12), 1697 => to_unsigned(2938, 12), 1698 => to_unsigned(1982, 12), 1699 => to_unsigned(1646, 12), 1700 => to_unsigned(1853, 12), 1701 => to_unsigned(1387, 12), 1702 => to_unsigned(3678, 12), 1703 => to_unsigned(2636, 12), 1704 => to_unsigned(4027, 12), 1705 => to_unsigned(3622, 12), 1706 => to_unsigned(1454, 12), 1707 => to_unsigned(287, 12), 1708 => to_unsigned(758, 12), 1709 => to_unsigned(178, 12), 1710 => to_unsigned(2597, 12), 1711 => to_unsigned(1831, 12), 1712 => to_unsigned(2156, 12), 1713 => to_unsigned(3187, 12), 1714 => to_unsigned(3550, 12), 1715 => to_unsigned(1393, 12), 1716 => to_unsigned(896, 12), 1717 => to_unsigned(3761, 12), 1718 => to_unsigned(1664, 12), 1719 => to_unsigned(2405, 12), 1720 => to_unsigned(497, 12), 1721 => to_unsigned(1015, 12), 1722 => to_unsigned(3260, 12), 1723 => to_unsigned(1131, 12), 1724 => to_unsigned(3610, 12), 1725 => to_unsigned(3812, 12), 1726 => to_unsigned(2153, 12), 1727 => to_unsigned(960, 12), 1728 => to_unsigned(3631, 12), 1729 => to_unsigned(564, 12), 1730 => to_unsigned(36, 12), 1731 => to_unsigned(215, 12), 1732 => to_unsigned(2281, 12), 1733 => to_unsigned(1081, 12), 1734 => to_unsigned(1123, 12), 1735 => to_unsigned(2458, 12), 1736 => to_unsigned(1079, 12), 1737 => to_unsigned(2873, 12), 1738 => to_unsigned(466, 12), 1739 => to_unsigned(661, 12), 1740 => to_unsigned(3950, 12), 1741 => to_unsigned(1020, 12), 1742 => to_unsigned(1789, 12), 1743 => to_unsigned(3454, 12), 1744 => to_unsigned(1477, 12), 1745 => to_unsigned(2659, 12), 1746 => to_unsigned(2102, 12), 1747 => to_unsigned(3156, 12), 1748 => to_unsigned(1173, 12), 1749 => to_unsigned(2044, 12), 1750 => to_unsigned(1620, 12), 1751 => to_unsigned(2028, 12), 1752 => to_unsigned(3699, 12), 1753 => to_unsigned(3496, 12), 1754 => to_unsigned(2423, 12), 1755 => to_unsigned(2574, 12), 1756 => to_unsigned(2117, 12), 1757 => to_unsigned(2792, 12), 1758 => to_unsigned(3730, 12), 1759 => to_unsigned(1698, 12), 1760 => to_unsigned(1560, 12), 1761 => to_unsigned(3018, 12), 1762 => to_unsigned(2830, 12), 1763 => to_unsigned(1226, 12), 1764 => to_unsigned(271, 12), 1765 => to_unsigned(3735, 12), 1766 => to_unsigned(3945, 12), 1767 => to_unsigned(833, 12), 1768 => to_unsigned(702, 12), 1769 => to_unsigned(3615, 12), 1770 => to_unsigned(1920, 12), 1771 => to_unsigned(1580, 12), 1772 => to_unsigned(3766, 12), 1773 => to_unsigned(1091, 12), 1774 => to_unsigned(3393, 12), 1775 => to_unsigned(3318, 12), 1776 => to_unsigned(360, 12), 1777 => to_unsigned(2557, 12), 1778 => to_unsigned(1320, 12), 1779 => to_unsigned(635, 12), 1780 => to_unsigned(3608, 12), 1781 => to_unsigned(2143, 12), 1782 => to_unsigned(3099, 12), 1783 => to_unsigned(2598, 12), 1784 => to_unsigned(1329, 12), 1785 => to_unsigned(1747, 12), 1786 => to_unsigned(2970, 12), 1787 => to_unsigned(1164, 12), 1788 => to_unsigned(2389, 12), 1789 => to_unsigned(2873, 12), 1790 => to_unsigned(3991, 12), 1791 => to_unsigned(2473, 12), 1792 => to_unsigned(1697, 12), 1793 => to_unsigned(3228, 12), 1794 => to_unsigned(1964, 12), 1795 => to_unsigned(2774, 12), 1796 => to_unsigned(75, 12), 1797 => to_unsigned(3075, 12), 1798 => to_unsigned(1774, 12), 1799 => to_unsigned(1410, 12), 1800 => to_unsigned(691, 12), 1801 => to_unsigned(3931, 12), 1802 => to_unsigned(2790, 12), 1803 => to_unsigned(490, 12), 1804 => to_unsigned(3322, 12), 1805 => to_unsigned(1763, 12), 1806 => to_unsigned(1879, 12), 1807 => to_unsigned(1602, 12), 1808 => to_unsigned(3137, 12), 1809 => to_unsigned(3520, 12), 1810 => to_unsigned(3062, 12), 1811 => to_unsigned(3320, 12), 1812 => to_unsigned(950, 12), 1813 => to_unsigned(620, 12), 1814 => to_unsigned(703, 12), 1815 => to_unsigned(1764, 12), 1816 => to_unsigned(281, 12), 1817 => to_unsigned(1949, 12), 1818 => to_unsigned(3937, 12), 1819 => to_unsigned(2266, 12), 1820 => to_unsigned(2103, 12), 1821 => to_unsigned(202, 12), 1822 => to_unsigned(1942, 12), 1823 => to_unsigned(1269, 12), 1824 => to_unsigned(195, 12), 1825 => to_unsigned(484, 12), 1826 => to_unsigned(3571, 12), 1827 => to_unsigned(3496, 12), 1828 => to_unsigned(2792, 12), 1829 => to_unsigned(751, 12), 1830 => to_unsigned(1342, 12), 1831 => to_unsigned(3610, 12), 1832 => to_unsigned(3766, 12), 1833 => to_unsigned(3764, 12), 1834 => to_unsigned(2175, 12), 1835 => to_unsigned(81, 12), 1836 => to_unsigned(2940, 12), 1837 => to_unsigned(1769, 12), 1838 => to_unsigned(2727, 12), 1839 => to_unsigned(3515, 12), 1840 => to_unsigned(2985, 12), 1841 => to_unsigned(525, 12), 1842 => to_unsigned(698, 12), 1843 => to_unsigned(188, 12), 1844 => to_unsigned(4041, 12), 1845 => to_unsigned(3893, 12), 1846 => to_unsigned(1925, 12), 1847 => to_unsigned(3931, 12), 1848 => to_unsigned(1118, 12), 1849 => to_unsigned(3673, 12), 1850 => to_unsigned(99, 12), 1851 => to_unsigned(447, 12), 1852 => to_unsigned(1209, 12), 1853 => to_unsigned(3696, 12), 1854 => to_unsigned(1698, 12), 1855 => to_unsigned(967, 12), 1856 => to_unsigned(3439, 12), 1857 => to_unsigned(3997, 12), 1858 => to_unsigned(815, 12), 1859 => to_unsigned(684, 12), 1860 => to_unsigned(2538, 12), 1861 => to_unsigned(2460, 12), 1862 => to_unsigned(2561, 12), 1863 => to_unsigned(762, 12), 1864 => to_unsigned(2176, 12), 1865 => to_unsigned(1969, 12), 1866 => to_unsigned(776, 12), 1867 => to_unsigned(1481, 12), 1868 => to_unsigned(3371, 12), 1869 => to_unsigned(932, 12), 1870 => to_unsigned(732, 12), 1871 => to_unsigned(1245, 12), 1872 => to_unsigned(288, 12), 1873 => to_unsigned(3440, 12), 1874 => to_unsigned(1655, 12), 1875 => to_unsigned(640, 12), 1876 => to_unsigned(3131, 12), 1877 => to_unsigned(969, 12), 1878 => to_unsigned(42, 12), 1879 => to_unsigned(1024, 12), 1880 => to_unsigned(2039, 12), 1881 => to_unsigned(1326, 12), 1882 => to_unsigned(3360, 12), 1883 => to_unsigned(253, 12), 1884 => to_unsigned(987, 12), 1885 => to_unsigned(1189, 12), 1886 => to_unsigned(1642, 12), 1887 => to_unsigned(3196, 12), 1888 => to_unsigned(869, 12), 1889 => to_unsigned(1943, 12), 1890 => to_unsigned(2536, 12), 1891 => to_unsigned(276, 12), 1892 => to_unsigned(1160, 12), 1893 => to_unsigned(3753, 12), 1894 => to_unsigned(1422, 12), 1895 => to_unsigned(1472, 12), 1896 => to_unsigned(2640, 12), 1897 => to_unsigned(4085, 12), 1898 => to_unsigned(3024, 12), 1899 => to_unsigned(2483, 12), 1900 => to_unsigned(3343, 12), 1901 => to_unsigned(2443, 12), 1902 => to_unsigned(432, 12), 1903 => to_unsigned(2955, 12), 1904 => to_unsigned(2883, 12), 1905 => to_unsigned(3426, 12), 1906 => to_unsigned(1592, 12), 1907 => to_unsigned(3702, 12), 1908 => to_unsigned(3523, 12), 1909 => to_unsigned(2380, 12), 1910 => to_unsigned(1876, 12), 1911 => to_unsigned(3490, 12), 1912 => to_unsigned(2861, 12), 1913 => to_unsigned(1679, 12), 1914 => to_unsigned(4087, 12), 1915 => to_unsigned(17, 12), 1916 => to_unsigned(972, 12), 1917 => to_unsigned(2362, 12), 1918 => to_unsigned(1047, 12), 1919 => to_unsigned(3149, 12), 1920 => to_unsigned(355, 12), 1921 => to_unsigned(1487, 12), 1922 => to_unsigned(2337, 12), 1923 => to_unsigned(1337, 12), 1924 => to_unsigned(3145, 12), 1925 => to_unsigned(3271, 12), 1926 => to_unsigned(2741, 12), 1927 => to_unsigned(500, 12), 1928 => to_unsigned(289, 12), 1929 => to_unsigned(2848, 12), 1930 => to_unsigned(15, 12), 1931 => to_unsigned(771, 12), 1932 => to_unsigned(1307, 12), 1933 => to_unsigned(2213, 12), 1934 => to_unsigned(878, 12), 1935 => to_unsigned(2009, 12), 1936 => to_unsigned(2353, 12), 1937 => to_unsigned(3119, 12), 1938 => to_unsigned(121, 12), 1939 => to_unsigned(3054, 12), 1940 => to_unsigned(219, 12), 1941 => to_unsigned(1521, 12), 1942 => to_unsigned(1753, 12), 1943 => to_unsigned(2283, 12), 1944 => to_unsigned(1282, 12), 1945 => to_unsigned(2998, 12), 1946 => to_unsigned(3595, 12), 1947 => to_unsigned(1906, 12), 1948 => to_unsigned(3308, 12), 1949 => to_unsigned(1804, 12), 1950 => to_unsigned(2250, 12), 1951 => to_unsigned(1131, 12), 1952 => to_unsigned(4078, 12), 1953 => to_unsigned(2255, 12), 1954 => to_unsigned(2880, 12), 1955 => to_unsigned(715, 12), 1956 => to_unsigned(1035, 12), 1957 => to_unsigned(2575, 12), 1958 => to_unsigned(1959, 12), 1959 => to_unsigned(82, 12), 1960 => to_unsigned(950, 12), 1961 => to_unsigned(573, 12), 1962 => to_unsigned(312, 12), 1963 => to_unsigned(112, 12), 1964 => to_unsigned(3436, 12), 1965 => to_unsigned(2287, 12), 1966 => to_unsigned(432, 12), 1967 => to_unsigned(2290, 12), 1968 => to_unsigned(1786, 12), 1969 => to_unsigned(1823, 12), 1970 => to_unsigned(3648, 12), 1971 => to_unsigned(3320, 12), 1972 => to_unsigned(3619, 12), 1973 => to_unsigned(3530, 12), 1974 => to_unsigned(3921, 12), 1975 => to_unsigned(734, 12), 1976 => to_unsigned(291, 12), 1977 => to_unsigned(46, 12), 1978 => to_unsigned(1114, 12), 1979 => to_unsigned(3943, 12), 1980 => to_unsigned(2394, 12), 1981 => to_unsigned(332, 12), 1982 => to_unsigned(421, 12), 1983 => to_unsigned(2899, 12), 1984 => to_unsigned(582, 12), 1985 => to_unsigned(2138, 12), 1986 => to_unsigned(2614, 12), 1987 => to_unsigned(67, 12), 1988 => to_unsigned(666, 12), 1989 => to_unsigned(3970, 12), 1990 => to_unsigned(3369, 12), 1991 => to_unsigned(580, 12), 1992 => to_unsigned(3819, 12), 1993 => to_unsigned(1866, 12), 1994 => to_unsigned(1651, 12), 1995 => to_unsigned(867, 12), 1996 => to_unsigned(543, 12), 1997 => to_unsigned(712, 12), 1998 => to_unsigned(294, 12), 1999 => to_unsigned(2835, 12), 2000 => to_unsigned(2704, 12), 2001 => to_unsigned(1363, 12), 2002 => to_unsigned(2147, 12), 2003 => to_unsigned(1807, 12), 2004 => to_unsigned(1344, 12), 2005 => to_unsigned(2799, 12), 2006 => to_unsigned(3516, 12), 2007 => to_unsigned(1606, 12), 2008 => to_unsigned(3342, 12), 2009 => to_unsigned(3067, 12), 2010 => to_unsigned(166, 12), 2011 => to_unsigned(786, 12), 2012 => to_unsigned(1332, 12), 2013 => to_unsigned(478, 12), 2014 => to_unsigned(3865, 12), 2015 => to_unsigned(347, 12), 2016 => to_unsigned(2217, 12), 2017 => to_unsigned(3948, 12), 2018 => to_unsigned(314, 12), 2019 => to_unsigned(1318, 12), 2020 => to_unsigned(3707, 12), 2021 => to_unsigned(1200, 12), 2022 => to_unsigned(3031, 12), 2023 => to_unsigned(2089, 12), 2024 => to_unsigned(1512, 12), 2025 => to_unsigned(3510, 12), 2026 => to_unsigned(3796, 12), 2027 => to_unsigned(2379, 12), 2028 => to_unsigned(3803, 12), 2029 => to_unsigned(1877, 12), 2030 => to_unsigned(3457, 12), 2031 => to_unsigned(2953, 12), 2032 => to_unsigned(1110, 12), 2033 => to_unsigned(2290, 12), 2034 => to_unsigned(2444, 12), 2035 => to_unsigned(225, 12), 2036 => to_unsigned(176, 12), 2037 => to_unsigned(693, 12), 2038 => to_unsigned(3822, 12), 2039 => to_unsigned(837, 12), 2040 => to_unsigned(3640, 12), 2041 => to_unsigned(955, 12), 2042 => to_unsigned(2652, 12), 2043 => to_unsigned(797, 12), 2044 => to_unsigned(3202, 12), 2045 => to_unsigned(1405, 12), 2046 => to_unsigned(3102, 12), 2047 => to_unsigned(2338, 12))
        ),
        1 => (
            0 => (0 => to_unsigned(1594, 12), 1 => to_unsigned(2289, 12), 2 => to_unsigned(332, 12), 3 => to_unsigned(1621, 12), 4 => to_unsigned(4044, 12), 5 => to_unsigned(80, 12), 6 => to_unsigned(2647, 12), 7 => to_unsigned(3786, 12), 8 => to_unsigned(3920, 12), 9 => to_unsigned(1109, 12), 10 => to_unsigned(2137, 12), 11 => to_unsigned(2067, 12), 12 => to_unsigned(2530, 12), 13 => to_unsigned(3991, 12), 14 => to_unsigned(1168, 12), 15 => to_unsigned(2412, 12), 16 => to_unsigned(2720, 12), 17 => to_unsigned(3649, 12), 18 => to_unsigned(2394, 12), 19 => to_unsigned(1549, 12), 20 => to_unsigned(286, 12), 21 => to_unsigned(163, 12), 22 => to_unsigned(3049, 12), 23 => to_unsigned(2348, 12), 24 => to_unsigned(2591, 12), 25 => to_unsigned(2217, 12), 26 => to_unsigned(4024, 12), 27 => to_unsigned(2518, 12), 28 => to_unsigned(3585, 12), 29 => to_unsigned(2558, 12), 30 => to_unsigned(767, 12), 31 => to_unsigned(399, 12), 32 => to_unsigned(415, 12), 33 => to_unsigned(2174, 12), 34 => to_unsigned(322, 12), 35 => to_unsigned(717, 12), 36 => to_unsigned(3584, 12), 37 => to_unsigned(3840, 12), 38 => to_unsigned(10, 12), 39 => to_unsigned(784, 12), 40 => to_unsigned(2808, 12), 41 => to_unsigned(1547, 12), 42 => to_unsigned(444, 12), 43 => to_unsigned(2009, 12), 44 => to_unsigned(2326, 12), 45 => to_unsigned(3327, 12), 46 => to_unsigned(2623, 12), 47 => to_unsigned(3909, 12), 48 => to_unsigned(1347, 12), 49 => to_unsigned(2670, 12), 50 => to_unsigned(1276, 12), 51 => to_unsigned(3347, 12), 52 => to_unsigned(2630, 12), 53 => to_unsigned(2355, 12), 54 => to_unsigned(2449, 12), 55 => to_unsigned(3383, 12), 56 => to_unsigned(400, 12), 57 => to_unsigned(1945, 12), 58 => to_unsigned(508, 12), 59 => to_unsigned(482, 12), 60 => to_unsigned(1206, 12), 61 => to_unsigned(3241, 12), 62 => to_unsigned(2001, 12), 63 => to_unsigned(3948, 12), 64 => to_unsigned(2456, 12), 65 => to_unsigned(2314, 12), 66 => to_unsigned(3698, 12), 67 => to_unsigned(3434, 12), 68 => to_unsigned(1306, 12), 69 => to_unsigned(4091, 12), 70 => to_unsigned(3127, 12), 71 => to_unsigned(2295, 12), 72 => to_unsigned(1636, 12), 73 => to_unsigned(3452, 12), 74 => to_unsigned(3294, 12), 75 => to_unsigned(3952, 12), 76 => to_unsigned(3794, 12), 77 => to_unsigned(3712, 12), 78 => to_unsigned(1027, 12), 79 => to_unsigned(1214, 12), 80 => to_unsigned(3170, 12), 81 => to_unsigned(3868, 12), 82 => to_unsigned(511, 12), 83 => to_unsigned(3839, 12), 84 => to_unsigned(3978, 12), 85 => to_unsigned(1617, 12), 86 => to_unsigned(3656, 12), 87 => to_unsigned(4029, 12), 88 => to_unsigned(2965, 12), 89 => to_unsigned(2479, 12), 90 => to_unsigned(1627, 12), 91 => to_unsigned(2126, 12), 92 => to_unsigned(2456, 12), 93 => to_unsigned(3922, 12), 94 => to_unsigned(802, 12), 95 => to_unsigned(3055, 12), 96 => to_unsigned(3066, 12), 97 => to_unsigned(3959, 12), 98 => to_unsigned(4051, 12), 99 => to_unsigned(1391, 12), 100 => to_unsigned(2652, 12), 101 => to_unsigned(4043, 12), 102 => to_unsigned(3794, 12), 103 => to_unsigned(2880, 12), 104 => to_unsigned(2470, 12), 105 => to_unsigned(3306, 12), 106 => to_unsigned(4079, 12), 107 => to_unsigned(2093, 12), 108 => to_unsigned(1316, 12), 109 => to_unsigned(1537, 12), 110 => to_unsigned(3112, 12), 111 => to_unsigned(2412, 12), 112 => to_unsigned(1119, 12), 113 => to_unsigned(1899, 12), 114 => to_unsigned(1649, 12), 115 => to_unsigned(352, 12), 116 => to_unsigned(1432, 12), 117 => to_unsigned(2240, 12), 118 => to_unsigned(1181, 12), 119 => to_unsigned(958, 12), 120 => to_unsigned(2551, 12), 121 => to_unsigned(1132, 12), 122 => to_unsigned(1250, 12), 123 => to_unsigned(1519, 12), 124 => to_unsigned(1010, 12), 125 => to_unsigned(4076, 12), 126 => to_unsigned(2732, 12), 127 => to_unsigned(3394, 12), 128 => to_unsigned(2578, 12), 129 => to_unsigned(2765, 12), 130 => to_unsigned(501, 12), 131 => to_unsigned(200, 12), 132 => to_unsigned(516, 12), 133 => to_unsigned(3347, 12), 134 => to_unsigned(2953, 12), 135 => to_unsigned(1117, 12), 136 => to_unsigned(576, 12), 137 => to_unsigned(2342, 12), 138 => to_unsigned(4081, 12), 139 => to_unsigned(534, 12), 140 => to_unsigned(921, 12), 141 => to_unsigned(539, 12), 142 => to_unsigned(2705, 12), 143 => to_unsigned(701, 12), 144 => to_unsigned(3770, 12), 145 => to_unsigned(2294, 12), 146 => to_unsigned(3417, 12), 147 => to_unsigned(118, 12), 148 => to_unsigned(3190, 12), 149 => to_unsigned(1131, 12), 150 => to_unsigned(3019, 12), 151 => to_unsigned(2502, 12), 152 => to_unsigned(1348, 12), 153 => to_unsigned(2718, 12), 154 => to_unsigned(2696, 12), 155 => to_unsigned(2876, 12), 156 => to_unsigned(3727, 12), 157 => to_unsigned(3603, 12), 158 => to_unsigned(144, 12), 159 => to_unsigned(1504, 12), 160 => to_unsigned(860, 12), 161 => to_unsigned(266, 12), 162 => to_unsigned(3770, 12), 163 => to_unsigned(2205, 12), 164 => to_unsigned(3789, 12), 165 => to_unsigned(3751, 12), 166 => to_unsigned(995, 12), 167 => to_unsigned(1393, 12), 168 => to_unsigned(2163, 12), 169 => to_unsigned(299, 12), 170 => to_unsigned(442, 12), 171 => to_unsigned(2027, 12), 172 => to_unsigned(2694, 12), 173 => to_unsigned(3178, 12), 174 => to_unsigned(518, 12), 175 => to_unsigned(1971, 12), 176 => to_unsigned(476, 12), 177 => to_unsigned(2089, 12), 178 => to_unsigned(1741, 12), 179 => to_unsigned(1764, 12), 180 => to_unsigned(2726, 12), 181 => to_unsigned(753, 12), 182 => to_unsigned(1684, 12), 183 => to_unsigned(113, 12), 184 => to_unsigned(3867, 12), 185 => to_unsigned(981, 12), 186 => to_unsigned(1123, 12), 187 => to_unsigned(782, 12), 188 => to_unsigned(2018, 12), 189 => to_unsigned(2930, 12), 190 => to_unsigned(3058, 12), 191 => to_unsigned(4072, 12), 192 => to_unsigned(2448, 12), 193 => to_unsigned(316, 12), 194 => to_unsigned(782, 12), 195 => to_unsigned(1185, 12), 196 => to_unsigned(2869, 12), 197 => to_unsigned(1428, 12), 198 => to_unsigned(2030, 12), 199 => to_unsigned(3408, 12), 200 => to_unsigned(2102, 12), 201 => to_unsigned(94, 12), 202 => to_unsigned(3882, 12), 203 => to_unsigned(1166, 12), 204 => to_unsigned(882, 12), 205 => to_unsigned(2965, 12), 206 => to_unsigned(3847, 12), 207 => to_unsigned(3257, 12), 208 => to_unsigned(3890, 12), 209 => to_unsigned(185, 12), 210 => to_unsigned(1697, 12), 211 => to_unsigned(3849, 12), 212 => to_unsigned(257, 12), 213 => to_unsigned(3016, 12), 214 => to_unsigned(3461, 12), 215 => to_unsigned(1134, 12), 216 => to_unsigned(1580, 12), 217 => to_unsigned(667, 12), 218 => to_unsigned(150, 12), 219 => to_unsigned(1795, 12), 220 => to_unsigned(827, 12), 221 => to_unsigned(2808, 12), 222 => to_unsigned(3027, 12), 223 => to_unsigned(3247, 12), 224 => to_unsigned(3896, 12), 225 => to_unsigned(2507, 12), 226 => to_unsigned(3123, 12), 227 => to_unsigned(1259, 12), 228 => to_unsigned(3140, 12), 229 => to_unsigned(1330, 12), 230 => to_unsigned(648, 12), 231 => to_unsigned(2148, 12), 232 => to_unsigned(163, 12), 233 => to_unsigned(565, 12), 234 => to_unsigned(1487, 12), 235 => to_unsigned(1041, 12), 236 => to_unsigned(1910, 12), 237 => to_unsigned(3541, 12), 238 => to_unsigned(571, 12), 239 => to_unsigned(322, 12), 240 => to_unsigned(4059, 12), 241 => to_unsigned(2631, 12), 242 => to_unsigned(1434, 12), 243 => to_unsigned(0, 12), 244 => to_unsigned(608, 12), 245 => to_unsigned(264, 12), 246 => to_unsigned(2367, 12), 247 => to_unsigned(4026, 12), 248 => to_unsigned(2119, 12), 249 => to_unsigned(442, 12), 250 => to_unsigned(92, 12), 251 => to_unsigned(879, 12), 252 => to_unsigned(2331, 12), 253 => to_unsigned(3405, 12), 254 => to_unsigned(1428, 12), 255 => to_unsigned(3775, 12), 256 => to_unsigned(2405, 12), 257 => to_unsigned(3217, 12), 258 => to_unsigned(2928, 12), 259 => to_unsigned(1112, 12), 260 => to_unsigned(2004, 12), 261 => to_unsigned(1092, 12), 262 => to_unsigned(3596, 12), 263 => to_unsigned(2059, 12), 264 => to_unsigned(1546, 12), 265 => to_unsigned(3640, 12), 266 => to_unsigned(1869, 12), 267 => to_unsigned(1082, 12), 268 => to_unsigned(523, 12), 269 => to_unsigned(3744, 12), 270 => to_unsigned(3292, 12), 271 => to_unsigned(2364, 12), 272 => to_unsigned(3019, 12), 273 => to_unsigned(423, 12), 274 => to_unsigned(965, 12), 275 => to_unsigned(2289, 12), 276 => to_unsigned(1651, 12), 277 => to_unsigned(2465, 12), 278 => to_unsigned(1764, 12), 279 => to_unsigned(3261, 12), 280 => to_unsigned(3425, 12), 281 => to_unsigned(3233, 12), 282 => to_unsigned(1542, 12), 283 => to_unsigned(2206, 12), 284 => to_unsigned(3558, 12), 285 => to_unsigned(859, 12), 286 => to_unsigned(2446, 12), 287 => to_unsigned(1121, 12), 288 => to_unsigned(2010, 12), 289 => to_unsigned(3043, 12), 290 => to_unsigned(3927, 12), 291 => to_unsigned(1492, 12), 292 => to_unsigned(2755, 12), 293 => to_unsigned(3030, 12), 294 => to_unsigned(325, 12), 295 => to_unsigned(1805, 12), 296 => to_unsigned(3231, 12), 297 => to_unsigned(755, 12), 298 => to_unsigned(719, 12), 299 => to_unsigned(2373, 12), 300 => to_unsigned(820, 12), 301 => to_unsigned(3153, 12), 302 => to_unsigned(870, 12), 303 => to_unsigned(2527, 12), 304 => to_unsigned(2163, 12), 305 => to_unsigned(344, 12), 306 => to_unsigned(3926, 12), 307 => to_unsigned(953, 12), 308 => to_unsigned(1809, 12), 309 => to_unsigned(2683, 12), 310 => to_unsigned(1214, 12), 311 => to_unsigned(836, 12), 312 => to_unsigned(1131, 12), 313 => to_unsigned(3025, 12), 314 => to_unsigned(3245, 12), 315 => to_unsigned(182, 12), 316 => to_unsigned(703, 12), 317 => to_unsigned(1513, 12), 318 => to_unsigned(1862, 12), 319 => to_unsigned(4076, 12), 320 => to_unsigned(2235, 12), 321 => to_unsigned(3797, 12), 322 => to_unsigned(3462, 12), 323 => to_unsigned(1836, 12), 324 => to_unsigned(2846, 12), 325 => to_unsigned(1588, 12), 326 => to_unsigned(2454, 12), 327 => to_unsigned(1520, 12), 328 => to_unsigned(1814, 12), 329 => to_unsigned(938, 12), 330 => to_unsigned(2101, 12), 331 => to_unsigned(305, 12), 332 => to_unsigned(2138, 12), 333 => to_unsigned(3496, 12), 334 => to_unsigned(2039, 12), 335 => to_unsigned(2893, 12), 336 => to_unsigned(3848, 12), 337 => to_unsigned(2351, 12), 338 => to_unsigned(2557, 12), 339 => to_unsigned(3980, 12), 340 => to_unsigned(3032, 12), 341 => to_unsigned(495, 12), 342 => to_unsigned(2047, 12), 343 => to_unsigned(3735, 12), 344 => to_unsigned(1650, 12), 345 => to_unsigned(805, 12), 346 => to_unsigned(2057, 12), 347 => to_unsigned(289, 12), 348 => to_unsigned(4088, 12), 349 => to_unsigned(604, 12), 350 => to_unsigned(2529, 12), 351 => to_unsigned(1674, 12), 352 => to_unsigned(898, 12), 353 => to_unsigned(2267, 12), 354 => to_unsigned(3214, 12), 355 => to_unsigned(1882, 12), 356 => to_unsigned(3843, 12), 357 => to_unsigned(1555, 12), 358 => to_unsigned(1471, 12), 359 => to_unsigned(3788, 12), 360 => to_unsigned(2615, 12), 361 => to_unsigned(3290, 12), 362 => to_unsigned(842, 12), 363 => to_unsigned(1842, 12), 364 => to_unsigned(920, 12), 365 => to_unsigned(996, 12), 366 => to_unsigned(2744, 12), 367 => to_unsigned(1907, 12), 368 => to_unsigned(4010, 12), 369 => to_unsigned(2046, 12), 370 => to_unsigned(4069, 12), 371 => to_unsigned(2436, 12), 372 => to_unsigned(515, 12), 373 => to_unsigned(964, 12), 374 => to_unsigned(3593, 12), 375 => to_unsigned(105, 12), 376 => to_unsigned(4047, 12), 377 => to_unsigned(2211, 12), 378 => to_unsigned(3690, 12), 379 => to_unsigned(3452, 12), 380 => to_unsigned(3715, 12), 381 => to_unsigned(966, 12), 382 => to_unsigned(2126, 12), 383 => to_unsigned(3864, 12), 384 => to_unsigned(1349, 12), 385 => to_unsigned(2856, 12), 386 => to_unsigned(1608, 12), 387 => to_unsigned(680, 12), 388 => to_unsigned(1166, 12), 389 => to_unsigned(3848, 12), 390 => to_unsigned(2792, 12), 391 => to_unsigned(1648, 12), 392 => to_unsigned(2083, 12), 393 => to_unsigned(1173, 12), 394 => to_unsigned(1667, 12), 395 => to_unsigned(678, 12), 396 => to_unsigned(2262, 12), 397 => to_unsigned(2245, 12), 398 => to_unsigned(2173, 12), 399 => to_unsigned(1536, 12), 400 => to_unsigned(1072, 12), 401 => to_unsigned(1173, 12), 402 => to_unsigned(3631, 12), 403 => to_unsigned(3680, 12), 404 => to_unsigned(816, 12), 405 => to_unsigned(4024, 12), 406 => to_unsigned(2951, 12), 407 => to_unsigned(3479, 12), 408 => to_unsigned(1412, 12), 409 => to_unsigned(2590, 12), 410 => to_unsigned(1393, 12), 411 => to_unsigned(397, 12), 412 => to_unsigned(3762, 12), 413 => to_unsigned(1777, 12), 414 => to_unsigned(2563, 12), 415 => to_unsigned(954, 12), 416 => to_unsigned(2244, 12), 417 => to_unsigned(1706, 12), 418 => to_unsigned(3737, 12), 419 => to_unsigned(3922, 12), 420 => to_unsigned(3100, 12), 421 => to_unsigned(3920, 12), 422 => to_unsigned(49, 12), 423 => to_unsigned(945, 12), 424 => to_unsigned(2446, 12), 425 => to_unsigned(2667, 12), 426 => to_unsigned(1892, 12), 427 => to_unsigned(3786, 12), 428 => to_unsigned(2919, 12), 429 => to_unsigned(3425, 12), 430 => to_unsigned(1598, 12), 431 => to_unsigned(1113, 12), 432 => to_unsigned(3510, 12), 433 => to_unsigned(3829, 12), 434 => to_unsigned(3035, 12), 435 => to_unsigned(1652, 12), 436 => to_unsigned(2383, 12), 437 => to_unsigned(1963, 12), 438 => to_unsigned(2801, 12), 439 => to_unsigned(2674, 12), 440 => to_unsigned(1272, 12), 441 => to_unsigned(1451, 12), 442 => to_unsigned(3881, 12), 443 => to_unsigned(414, 12), 444 => to_unsigned(3770, 12), 445 => to_unsigned(725, 12), 446 => to_unsigned(1349, 12), 447 => to_unsigned(3476, 12), 448 => to_unsigned(3997, 12), 449 => to_unsigned(3041, 12), 450 => to_unsigned(2873, 12), 451 => to_unsigned(1279, 12), 452 => to_unsigned(562, 12), 453 => to_unsigned(1484, 12), 454 => to_unsigned(3916, 12), 455 => to_unsigned(1126, 12), 456 => to_unsigned(1561, 12), 457 => to_unsigned(1542, 12), 458 => to_unsigned(1186, 12), 459 => to_unsigned(805, 12), 460 => to_unsigned(2986, 12), 461 => to_unsigned(753, 12), 462 => to_unsigned(2662, 12), 463 => to_unsigned(3888, 12), 464 => to_unsigned(1462, 12), 465 => to_unsigned(946, 12), 466 => to_unsigned(95, 12), 467 => to_unsigned(3782, 12), 468 => to_unsigned(2413, 12), 469 => to_unsigned(3848, 12), 470 => to_unsigned(4027, 12), 471 => to_unsigned(1149, 12), 472 => to_unsigned(670, 12), 473 => to_unsigned(678, 12), 474 => to_unsigned(990, 12), 475 => to_unsigned(1913, 12), 476 => to_unsigned(3997, 12), 477 => to_unsigned(1374, 12), 478 => to_unsigned(3586, 12), 479 => to_unsigned(1150, 12), 480 => to_unsigned(634, 12), 481 => to_unsigned(2260, 12), 482 => to_unsigned(1465, 12), 483 => to_unsigned(1106, 12), 484 => to_unsigned(2804, 12), 485 => to_unsigned(311, 12), 486 => to_unsigned(472, 12), 487 => to_unsigned(2779, 12), 488 => to_unsigned(3616, 12), 489 => to_unsigned(2900, 12), 490 => to_unsigned(3237, 12), 491 => to_unsigned(2549, 12), 492 => to_unsigned(1601, 12), 493 => to_unsigned(1790, 12), 494 => to_unsigned(1190, 12), 495 => to_unsigned(1485, 12), 496 => to_unsigned(2061, 12), 497 => to_unsigned(2518, 12), 498 => to_unsigned(3959, 12), 499 => to_unsigned(837, 12), 500 => to_unsigned(3553, 12), 501 => to_unsigned(899, 12), 502 => to_unsigned(1705, 12), 503 => to_unsigned(773, 12), 504 => to_unsigned(1438, 12), 505 => to_unsigned(1412, 12), 506 => to_unsigned(3831, 12), 507 => to_unsigned(3052, 12), 508 => to_unsigned(4080, 12), 509 => to_unsigned(2916, 12), 510 => to_unsigned(2938, 12), 511 => to_unsigned(1075, 12), 512 => to_unsigned(1638, 12), 513 => to_unsigned(897, 12), 514 => to_unsigned(2827, 12), 515 => to_unsigned(946, 12), 516 => to_unsigned(3704, 12), 517 => to_unsigned(3411, 12), 518 => to_unsigned(2516, 12), 519 => to_unsigned(847, 12), 520 => to_unsigned(2112, 12), 521 => to_unsigned(2047, 12), 522 => to_unsigned(237, 12), 523 => to_unsigned(3509, 12), 524 => to_unsigned(294, 12), 525 => to_unsigned(344, 12), 526 => to_unsigned(2969, 12), 527 => to_unsigned(1130, 12), 528 => to_unsigned(3187, 12), 529 => to_unsigned(1998, 12), 530 => to_unsigned(2704, 12), 531 => to_unsigned(2914, 12), 532 => to_unsigned(2973, 12), 533 => to_unsigned(1717, 12), 534 => to_unsigned(2033, 12), 535 => to_unsigned(1368, 12), 536 => to_unsigned(2232, 12), 537 => to_unsigned(3993, 12), 538 => to_unsigned(2302, 12), 539 => to_unsigned(3342, 12), 540 => to_unsigned(2140, 12), 541 => to_unsigned(3155, 12), 542 => to_unsigned(1983, 12), 543 => to_unsigned(2184, 12), 544 => to_unsigned(3198, 12), 545 => to_unsigned(2131, 12), 546 => to_unsigned(3836, 12), 547 => to_unsigned(1184, 12), 548 => to_unsigned(1174, 12), 549 => to_unsigned(1296, 12), 550 => to_unsigned(2089, 12), 551 => to_unsigned(2207, 12), 552 => to_unsigned(1732, 12), 553 => to_unsigned(1044, 12), 554 => to_unsigned(2670, 12), 555 => to_unsigned(77, 12), 556 => to_unsigned(62, 12), 557 => to_unsigned(272, 12), 558 => to_unsigned(3021, 12), 559 => to_unsigned(218, 12), 560 => to_unsigned(1016, 12), 561 => to_unsigned(3616, 12), 562 => to_unsigned(198, 12), 563 => to_unsigned(1405, 12), 564 => to_unsigned(3301, 12), 565 => to_unsigned(3800, 12), 566 => to_unsigned(2825, 12), 567 => to_unsigned(2036, 12), 568 => to_unsigned(1493, 12), 569 => to_unsigned(3348, 12), 570 => to_unsigned(1692, 12), 571 => to_unsigned(1871, 12), 572 => to_unsigned(3087, 12), 573 => to_unsigned(1388, 12), 574 => to_unsigned(2572, 12), 575 => to_unsigned(3423, 12), 576 => to_unsigned(1068, 12), 577 => to_unsigned(3886, 12), 578 => to_unsigned(119, 12), 579 => to_unsigned(823, 12), 580 => to_unsigned(589, 12), 581 => to_unsigned(338, 12), 582 => to_unsigned(2521, 12), 583 => to_unsigned(900, 12), 584 => to_unsigned(1349, 12), 585 => to_unsigned(2462, 12), 586 => to_unsigned(2312, 12), 587 => to_unsigned(1766, 12), 588 => to_unsigned(3714, 12), 589 => to_unsigned(1953, 12), 590 => to_unsigned(2338, 12), 591 => to_unsigned(847, 12), 592 => to_unsigned(546, 12), 593 => to_unsigned(2912, 12), 594 => to_unsigned(3587, 12), 595 => to_unsigned(2618, 12), 596 => to_unsigned(4020, 12), 597 => to_unsigned(2282, 12), 598 => to_unsigned(2105, 12), 599 => to_unsigned(1787, 12), 600 => to_unsigned(451, 12), 601 => to_unsigned(853, 12), 602 => to_unsigned(2871, 12), 603 => to_unsigned(3876, 12), 604 => to_unsigned(4029, 12), 605 => to_unsigned(186, 12), 606 => to_unsigned(2630, 12), 607 => to_unsigned(3157, 12), 608 => to_unsigned(3449, 12), 609 => to_unsigned(1806, 12), 610 => to_unsigned(373, 12), 611 => to_unsigned(14, 12), 612 => to_unsigned(3793, 12), 613 => to_unsigned(350, 12), 614 => to_unsigned(1083, 12), 615 => to_unsigned(2515, 12), 616 => to_unsigned(2924, 12), 617 => to_unsigned(2541, 12), 618 => to_unsigned(3682, 12), 619 => to_unsigned(1376, 12), 620 => to_unsigned(3680, 12), 621 => to_unsigned(477, 12), 622 => to_unsigned(3126, 12), 623 => to_unsigned(23, 12), 624 => to_unsigned(1350, 12), 625 => to_unsigned(1386, 12), 626 => to_unsigned(55, 12), 627 => to_unsigned(991, 12), 628 => to_unsigned(3120, 12), 629 => to_unsigned(3734, 12), 630 => to_unsigned(2134, 12), 631 => to_unsigned(4022, 12), 632 => to_unsigned(2027, 12), 633 => to_unsigned(3424, 12), 634 => to_unsigned(897, 12), 635 => to_unsigned(1533, 12), 636 => to_unsigned(852, 12), 637 => to_unsigned(1684, 12), 638 => to_unsigned(3725, 12), 639 => to_unsigned(3390, 12), 640 => to_unsigned(1990, 12), 641 => to_unsigned(2405, 12), 642 => to_unsigned(3646, 12), 643 => to_unsigned(2224, 12), 644 => to_unsigned(3874, 12), 645 => to_unsigned(229, 12), 646 => to_unsigned(3558, 12), 647 => to_unsigned(3028, 12), 648 => to_unsigned(1005, 12), 649 => to_unsigned(2594, 12), 650 => to_unsigned(3379, 12), 651 => to_unsigned(1162, 12), 652 => to_unsigned(3669, 12), 653 => to_unsigned(350, 12), 654 => to_unsigned(170, 12), 655 => to_unsigned(897, 12), 656 => to_unsigned(2566, 12), 657 => to_unsigned(2204, 12), 658 => to_unsigned(2892, 12), 659 => to_unsigned(1968, 12), 660 => to_unsigned(2363, 12), 661 => to_unsigned(2482, 12), 662 => to_unsigned(1215, 12), 663 => to_unsigned(1355, 12), 664 => to_unsigned(746, 12), 665 => to_unsigned(1716, 12), 666 => to_unsigned(1397, 12), 667 => to_unsigned(1100, 12), 668 => to_unsigned(3823, 12), 669 => to_unsigned(3120, 12), 670 => to_unsigned(2437, 12), 671 => to_unsigned(3374, 12), 672 => to_unsigned(759, 12), 673 => to_unsigned(852, 12), 674 => to_unsigned(2575, 12), 675 => to_unsigned(2064, 12), 676 => to_unsigned(3955, 12), 677 => to_unsigned(2540, 12), 678 => to_unsigned(320, 12), 679 => to_unsigned(3481, 12), 680 => to_unsigned(3431, 12), 681 => to_unsigned(2404, 12), 682 => to_unsigned(1384, 12), 683 => to_unsigned(2239, 12), 684 => to_unsigned(3109, 12), 685 => to_unsigned(3951, 12), 686 => to_unsigned(2845, 12), 687 => to_unsigned(2473, 12), 688 => to_unsigned(3403, 12), 689 => to_unsigned(4009, 12), 690 => to_unsigned(90, 12), 691 => to_unsigned(646, 12), 692 => to_unsigned(3798, 12), 693 => to_unsigned(2536, 12), 694 => to_unsigned(1249, 12), 695 => to_unsigned(364, 12), 696 => to_unsigned(2333, 12), 697 => to_unsigned(1874, 12), 698 => to_unsigned(3034, 12), 699 => to_unsigned(2635, 12), 700 => to_unsigned(4085, 12), 701 => to_unsigned(1457, 12), 702 => to_unsigned(4053, 12), 703 => to_unsigned(1160, 12), 704 => to_unsigned(3434, 12), 705 => to_unsigned(2477, 12), 706 => to_unsigned(2025, 12), 707 => to_unsigned(944, 12), 708 => to_unsigned(1184, 12), 709 => to_unsigned(410, 12), 710 => to_unsigned(2319, 12), 711 => to_unsigned(690, 12), 712 => to_unsigned(208, 12), 713 => to_unsigned(1664, 12), 714 => to_unsigned(2633, 12), 715 => to_unsigned(1640, 12), 716 => to_unsigned(1927, 12), 717 => to_unsigned(1245, 12), 718 => to_unsigned(1507, 12), 719 => to_unsigned(3456, 12), 720 => to_unsigned(1008, 12), 721 => to_unsigned(4000, 12), 722 => to_unsigned(3040, 12), 723 => to_unsigned(398, 12), 724 => to_unsigned(2610, 12), 725 => to_unsigned(3143, 12), 726 => to_unsigned(2658, 12), 727 => to_unsigned(1304, 12), 728 => to_unsigned(802, 12), 729 => to_unsigned(3728, 12), 730 => to_unsigned(778, 12), 731 => to_unsigned(3638, 12), 732 => to_unsigned(3826, 12), 733 => to_unsigned(9, 12), 734 => to_unsigned(1419, 12), 735 => to_unsigned(1004, 12), 736 => to_unsigned(3732, 12), 737 => to_unsigned(446, 12), 738 => to_unsigned(531, 12), 739 => to_unsigned(429, 12), 740 => to_unsigned(340, 12), 741 => to_unsigned(2016, 12), 742 => to_unsigned(2290, 12), 743 => to_unsigned(1302, 12), 744 => to_unsigned(3031, 12), 745 => to_unsigned(241, 12), 746 => to_unsigned(2909, 12), 747 => to_unsigned(3927, 12), 748 => to_unsigned(1087, 12), 749 => to_unsigned(1968, 12), 750 => to_unsigned(454, 12), 751 => to_unsigned(3701, 12), 752 => to_unsigned(434, 12), 753 => to_unsigned(2231, 12), 754 => to_unsigned(2373, 12), 755 => to_unsigned(3726, 12), 756 => to_unsigned(2123, 12), 757 => to_unsigned(2074, 12), 758 => to_unsigned(1740, 12), 759 => to_unsigned(3878, 12), 760 => to_unsigned(2979, 12), 761 => to_unsigned(3885, 12), 762 => to_unsigned(4005, 12), 763 => to_unsigned(3105, 12), 764 => to_unsigned(923, 12), 765 => to_unsigned(299, 12), 766 => to_unsigned(1342, 12), 767 => to_unsigned(2392, 12), 768 => to_unsigned(555, 12), 769 => to_unsigned(2852, 12), 770 => to_unsigned(104, 12), 771 => to_unsigned(1581, 12), 772 => to_unsigned(2720, 12), 773 => to_unsigned(3202, 12), 774 => to_unsigned(2306, 12), 775 => to_unsigned(2252, 12), 776 => to_unsigned(3863, 12), 777 => to_unsigned(2645, 12), 778 => to_unsigned(1520, 12), 779 => to_unsigned(1927, 12), 780 => to_unsigned(2658, 12), 781 => to_unsigned(1503, 12), 782 => to_unsigned(3395, 12), 783 => to_unsigned(954, 12), 784 => to_unsigned(2502, 12), 785 => to_unsigned(1948, 12), 786 => to_unsigned(296, 12), 787 => to_unsigned(1490, 12), 788 => to_unsigned(1968, 12), 789 => to_unsigned(564, 12), 790 => to_unsigned(3788, 12), 791 => to_unsigned(1217, 12), 792 => to_unsigned(2189, 12), 793 => to_unsigned(3528, 12), 794 => to_unsigned(30, 12), 795 => to_unsigned(2767, 12), 796 => to_unsigned(2104, 12), 797 => to_unsigned(49, 12), 798 => to_unsigned(3045, 12), 799 => to_unsigned(3932, 12), 800 => to_unsigned(3301, 12), 801 => to_unsigned(3680, 12), 802 => to_unsigned(3867, 12), 803 => to_unsigned(3805, 12), 804 => to_unsigned(857, 12), 805 => to_unsigned(1700, 12), 806 => to_unsigned(2187, 12), 807 => to_unsigned(3154, 12), 808 => to_unsigned(1849, 12), 809 => to_unsigned(716, 12), 810 => to_unsigned(2261, 12), 811 => to_unsigned(3910, 12), 812 => to_unsigned(1993, 12), 813 => to_unsigned(485, 12), 814 => to_unsigned(3493, 12), 815 => to_unsigned(1579, 12), 816 => to_unsigned(256, 12), 817 => to_unsigned(3177, 12), 818 => to_unsigned(1989, 12), 819 => to_unsigned(3418, 12), 820 => to_unsigned(1060, 12), 821 => to_unsigned(2445, 12), 822 => to_unsigned(1038, 12), 823 => to_unsigned(1587, 12), 824 => to_unsigned(551, 12), 825 => to_unsigned(3644, 12), 826 => to_unsigned(3730, 12), 827 => to_unsigned(2555, 12), 828 => to_unsigned(1401, 12), 829 => to_unsigned(1960, 12), 830 => to_unsigned(1413, 12), 831 => to_unsigned(3838, 12), 832 => to_unsigned(3286, 12), 833 => to_unsigned(2678, 12), 834 => to_unsigned(2824, 12), 835 => to_unsigned(3832, 12), 836 => to_unsigned(227, 12), 837 => to_unsigned(3854, 12), 838 => to_unsigned(363, 12), 839 => to_unsigned(2739, 12), 840 => to_unsigned(4041, 12), 841 => to_unsigned(3437, 12), 842 => to_unsigned(105, 12), 843 => to_unsigned(1980, 12), 844 => to_unsigned(656, 12), 845 => to_unsigned(3690, 12), 846 => to_unsigned(786, 12), 847 => to_unsigned(3374, 12), 848 => to_unsigned(2340, 12), 849 => to_unsigned(3421, 12), 850 => to_unsigned(4082, 12), 851 => to_unsigned(1473, 12), 852 => to_unsigned(4071, 12), 853 => to_unsigned(2517, 12), 854 => to_unsigned(2810, 12), 855 => to_unsigned(3889, 12), 856 => to_unsigned(2339, 12), 857 => to_unsigned(343, 12), 858 => to_unsigned(708, 12), 859 => to_unsigned(1533, 12), 860 => to_unsigned(1857, 12), 861 => to_unsigned(758, 12), 862 => to_unsigned(533, 12), 863 => to_unsigned(1971, 12), 864 => to_unsigned(1311, 12), 865 => to_unsigned(1379, 12), 866 => to_unsigned(1158, 12), 867 => to_unsigned(514, 12), 868 => to_unsigned(655, 12), 869 => to_unsigned(3771, 12), 870 => to_unsigned(2037, 12), 871 => to_unsigned(2746, 12), 872 => to_unsigned(250, 12), 873 => to_unsigned(551, 12), 874 => to_unsigned(2964, 12), 875 => to_unsigned(288, 12), 876 => to_unsigned(216, 12), 877 => to_unsigned(2978, 12), 878 => to_unsigned(2758, 12), 879 => to_unsigned(2875, 12), 880 => to_unsigned(1462, 12), 881 => to_unsigned(2804, 12), 882 => to_unsigned(1768, 12), 883 => to_unsigned(1161, 12), 884 => to_unsigned(2091, 12), 885 => to_unsigned(2573, 12), 886 => to_unsigned(2249, 12), 887 => to_unsigned(2168, 12), 888 => to_unsigned(2900, 12), 889 => to_unsigned(1869, 12), 890 => to_unsigned(1782, 12), 891 => to_unsigned(3213, 12), 892 => to_unsigned(3572, 12), 893 => to_unsigned(2764, 12), 894 => to_unsigned(1493, 12), 895 => to_unsigned(634, 12), 896 => to_unsigned(1317, 12), 897 => to_unsigned(3276, 12), 898 => to_unsigned(3150, 12), 899 => to_unsigned(3529, 12), 900 => to_unsigned(1895, 12), 901 => to_unsigned(3355, 12), 902 => to_unsigned(2533, 12), 903 => to_unsigned(2014, 12), 904 => to_unsigned(1811, 12), 905 => to_unsigned(356, 12), 906 => to_unsigned(277, 12), 907 => to_unsigned(6, 12), 908 => to_unsigned(611, 12), 909 => to_unsigned(2882, 12), 910 => to_unsigned(3829, 12), 911 => to_unsigned(2342, 12), 912 => to_unsigned(2579, 12), 913 => to_unsigned(1796, 12), 914 => to_unsigned(2768, 12), 915 => to_unsigned(3281, 12), 916 => to_unsigned(3750, 12), 917 => to_unsigned(2637, 12), 918 => to_unsigned(1406, 12), 919 => to_unsigned(1771, 12), 920 => to_unsigned(1966, 12), 921 => to_unsigned(1701, 12), 922 => to_unsigned(3353, 12), 923 => to_unsigned(1549, 12), 924 => to_unsigned(981, 12), 925 => to_unsigned(2492, 12), 926 => to_unsigned(293, 12), 927 => to_unsigned(2346, 12), 928 => to_unsigned(2409, 12), 929 => to_unsigned(1768, 12), 930 => to_unsigned(260, 12), 931 => to_unsigned(3674, 12), 932 => to_unsigned(1977, 12), 933 => to_unsigned(2006, 12), 934 => to_unsigned(334, 12), 935 => to_unsigned(3313, 12), 936 => to_unsigned(3918, 12), 937 => to_unsigned(42, 12), 938 => to_unsigned(2771, 12), 939 => to_unsigned(921, 12), 940 => to_unsigned(2910, 12), 941 => to_unsigned(2224, 12), 942 => to_unsigned(36, 12), 943 => to_unsigned(1931, 12), 944 => to_unsigned(2998, 12), 945 => to_unsigned(1758, 12), 946 => to_unsigned(570, 12), 947 => to_unsigned(1558, 12), 948 => to_unsigned(1601, 12), 949 => to_unsigned(1899, 12), 950 => to_unsigned(628, 12), 951 => to_unsigned(2458, 12), 952 => to_unsigned(976, 12), 953 => to_unsigned(656, 12), 954 => to_unsigned(3808, 12), 955 => to_unsigned(208, 12), 956 => to_unsigned(837, 12), 957 => to_unsigned(2186, 12), 958 => to_unsigned(4043, 12), 959 => to_unsigned(533, 12), 960 => to_unsigned(2276, 12), 961 => to_unsigned(3491, 12), 962 => to_unsigned(3824, 12), 963 => to_unsigned(3132, 12), 964 => to_unsigned(3798, 12), 965 => to_unsigned(1504, 12), 966 => to_unsigned(3513, 12), 967 => to_unsigned(2528, 12), 968 => to_unsigned(529, 12), 969 => to_unsigned(2125, 12), 970 => to_unsigned(2451, 12), 971 => to_unsigned(1877, 12), 972 => to_unsigned(759, 12), 973 => to_unsigned(2794, 12), 974 => to_unsigned(580, 12), 975 => to_unsigned(600, 12), 976 => to_unsigned(2391, 12), 977 => to_unsigned(2945, 12), 978 => to_unsigned(2951, 12), 979 => to_unsigned(1578, 12), 980 => to_unsigned(1098, 12), 981 => to_unsigned(3841, 12), 982 => to_unsigned(3862, 12), 983 => to_unsigned(2354, 12), 984 => to_unsigned(4039, 12), 985 => to_unsigned(649, 12), 986 => to_unsigned(220, 12), 987 => to_unsigned(3835, 12), 988 => to_unsigned(3884, 12), 989 => to_unsigned(3963, 12), 990 => to_unsigned(3305, 12), 991 => to_unsigned(1838, 12), 992 => to_unsigned(3987, 12), 993 => to_unsigned(2298, 12), 994 => to_unsigned(1127, 12), 995 => to_unsigned(453, 12), 996 => to_unsigned(2138, 12), 997 => to_unsigned(264, 12), 998 => to_unsigned(2617, 12), 999 => to_unsigned(1068, 12), 1000 => to_unsigned(3157, 12), 1001 => to_unsigned(1169, 12), 1002 => to_unsigned(2693, 12), 1003 => to_unsigned(1998, 12), 1004 => to_unsigned(352, 12), 1005 => to_unsigned(2341, 12), 1006 => to_unsigned(1691, 12), 1007 => to_unsigned(4062, 12), 1008 => to_unsigned(3133, 12), 1009 => to_unsigned(828, 12), 1010 => to_unsigned(3260, 12), 1011 => to_unsigned(2490, 12), 1012 => to_unsigned(2232, 12), 1013 => to_unsigned(3014, 12), 1014 => to_unsigned(3276, 12), 1015 => to_unsigned(1611, 12), 1016 => to_unsigned(3227, 12), 1017 => to_unsigned(628, 12), 1018 => to_unsigned(209, 12), 1019 => to_unsigned(2770, 12), 1020 => to_unsigned(1231, 12), 1021 => to_unsigned(2820, 12), 1022 => to_unsigned(2576, 12), 1023 => to_unsigned(891, 12), 1024 => to_unsigned(359, 12), 1025 => to_unsigned(3656, 12), 1026 => to_unsigned(139, 12), 1027 => to_unsigned(937, 12), 1028 => to_unsigned(3114, 12), 1029 => to_unsigned(4030, 12), 1030 => to_unsigned(3852, 12), 1031 => to_unsigned(2173, 12), 1032 => to_unsigned(1828, 12), 1033 => to_unsigned(534, 12), 1034 => to_unsigned(2938, 12), 1035 => to_unsigned(981, 12), 1036 => to_unsigned(1148, 12), 1037 => to_unsigned(683, 12), 1038 => to_unsigned(1660, 12), 1039 => to_unsigned(318, 12), 1040 => to_unsigned(639, 12), 1041 => to_unsigned(2377, 12), 1042 => to_unsigned(376, 12), 1043 => to_unsigned(2171, 12), 1044 => to_unsigned(1868, 12), 1045 => to_unsigned(3025, 12), 1046 => to_unsigned(3287, 12), 1047 => to_unsigned(2740, 12), 1048 => to_unsigned(3127, 12), 1049 => to_unsigned(1167, 12), 1050 => to_unsigned(387, 12), 1051 => to_unsigned(351, 12), 1052 => to_unsigned(1082, 12), 1053 => to_unsigned(1277, 12), 1054 => to_unsigned(2351, 12), 1055 => to_unsigned(189, 12), 1056 => to_unsigned(3211, 12), 1057 => to_unsigned(1440, 12), 1058 => to_unsigned(2666, 12), 1059 => to_unsigned(3535, 12), 1060 => to_unsigned(3993, 12), 1061 => to_unsigned(3215, 12), 1062 => to_unsigned(2881, 12), 1063 => to_unsigned(605, 12), 1064 => to_unsigned(3600, 12), 1065 => to_unsigned(29, 12), 1066 => to_unsigned(2360, 12), 1067 => to_unsigned(2404, 12), 1068 => to_unsigned(2653, 12), 1069 => to_unsigned(448, 12), 1070 => to_unsigned(3645, 12), 1071 => to_unsigned(1783, 12), 1072 => to_unsigned(2343, 12), 1073 => to_unsigned(2902, 12), 1074 => to_unsigned(1282, 12), 1075 => to_unsigned(2405, 12), 1076 => to_unsigned(3760, 12), 1077 => to_unsigned(1278, 12), 1078 => to_unsigned(2835, 12), 1079 => to_unsigned(1735, 12), 1080 => to_unsigned(910, 12), 1081 => to_unsigned(1506, 12), 1082 => to_unsigned(2974, 12), 1083 => to_unsigned(3459, 12), 1084 => to_unsigned(2634, 12), 1085 => to_unsigned(1656, 12), 1086 => to_unsigned(236, 12), 1087 => to_unsigned(1558, 12), 1088 => to_unsigned(2863, 12), 1089 => to_unsigned(3818, 12), 1090 => to_unsigned(3894, 12), 1091 => to_unsigned(238, 12), 1092 => to_unsigned(3031, 12), 1093 => to_unsigned(2992, 12), 1094 => to_unsigned(3199, 12), 1095 => to_unsigned(73, 12), 1096 => to_unsigned(545, 12), 1097 => to_unsigned(2929, 12), 1098 => to_unsigned(3290, 12), 1099 => to_unsigned(1160, 12), 1100 => to_unsigned(1181, 12), 1101 => to_unsigned(1372, 12), 1102 => to_unsigned(993, 12), 1103 => to_unsigned(3249, 12), 1104 => to_unsigned(1384, 12), 1105 => to_unsigned(3317, 12), 1106 => to_unsigned(182, 12), 1107 => to_unsigned(2988, 12), 1108 => to_unsigned(2940, 12), 1109 => to_unsigned(146, 12), 1110 => to_unsigned(2510, 12), 1111 => to_unsigned(1794, 12), 1112 => to_unsigned(1000, 12), 1113 => to_unsigned(650, 12), 1114 => to_unsigned(2265, 12), 1115 => to_unsigned(3398, 12), 1116 => to_unsigned(1180, 12), 1117 => to_unsigned(3125, 12), 1118 => to_unsigned(3548, 12), 1119 => to_unsigned(3472, 12), 1120 => to_unsigned(1767, 12), 1121 => to_unsigned(2133, 12), 1122 => to_unsigned(3158, 12), 1123 => to_unsigned(2109, 12), 1124 => to_unsigned(3576, 12), 1125 => to_unsigned(722, 12), 1126 => to_unsigned(128, 12), 1127 => to_unsigned(968, 12), 1128 => to_unsigned(2417, 12), 1129 => to_unsigned(3394, 12), 1130 => to_unsigned(3771, 12), 1131 => to_unsigned(4086, 12), 1132 => to_unsigned(3081, 12), 1133 => to_unsigned(3363, 12), 1134 => to_unsigned(3917, 12), 1135 => to_unsigned(1386, 12), 1136 => to_unsigned(2490, 12), 1137 => to_unsigned(1628, 12), 1138 => to_unsigned(2476, 12), 1139 => to_unsigned(1941, 12), 1140 => to_unsigned(3072, 12), 1141 => to_unsigned(1747, 12), 1142 => to_unsigned(456, 12), 1143 => to_unsigned(3362, 12), 1144 => to_unsigned(954, 12), 1145 => to_unsigned(2136, 12), 1146 => to_unsigned(1843, 12), 1147 => to_unsigned(3402, 12), 1148 => to_unsigned(1524, 12), 1149 => to_unsigned(2157, 12), 1150 => to_unsigned(908, 12), 1151 => to_unsigned(3845, 12), 1152 => to_unsigned(2020, 12), 1153 => to_unsigned(3753, 12), 1154 => to_unsigned(2932, 12), 1155 => to_unsigned(2632, 12), 1156 => to_unsigned(2242, 12), 1157 => to_unsigned(3703, 12), 1158 => to_unsigned(3314, 12), 1159 => to_unsigned(1752, 12), 1160 => to_unsigned(2793, 12), 1161 => to_unsigned(874, 12), 1162 => to_unsigned(666, 12), 1163 => to_unsigned(2642, 12), 1164 => to_unsigned(1061, 12), 1165 => to_unsigned(2090, 12), 1166 => to_unsigned(3838, 12), 1167 => to_unsigned(1231, 12), 1168 => to_unsigned(145, 12), 1169 => to_unsigned(360, 12), 1170 => to_unsigned(1167, 12), 1171 => to_unsigned(1265, 12), 1172 => to_unsigned(3056, 12), 1173 => to_unsigned(2176, 12), 1174 => to_unsigned(1641, 12), 1175 => to_unsigned(3040, 12), 1176 => to_unsigned(3438, 12), 1177 => to_unsigned(3959, 12), 1178 => to_unsigned(3798, 12), 1179 => to_unsigned(675, 12), 1180 => to_unsigned(398, 12), 1181 => to_unsigned(2173, 12), 1182 => to_unsigned(1568, 12), 1183 => to_unsigned(288, 12), 1184 => to_unsigned(2765, 12), 1185 => to_unsigned(2362, 12), 1186 => to_unsigned(3221, 12), 1187 => to_unsigned(1174, 12), 1188 => to_unsigned(2570, 12), 1189 => to_unsigned(2581, 12), 1190 => to_unsigned(1399, 12), 1191 => to_unsigned(979, 12), 1192 => to_unsigned(1665, 12), 1193 => to_unsigned(1961, 12), 1194 => to_unsigned(3811, 12), 1195 => to_unsigned(976, 12), 1196 => to_unsigned(3528, 12), 1197 => to_unsigned(3075, 12), 1198 => to_unsigned(1142, 12), 1199 => to_unsigned(2773, 12), 1200 => to_unsigned(3343, 12), 1201 => to_unsigned(2072, 12), 1202 => to_unsigned(3485, 12), 1203 => to_unsigned(983, 12), 1204 => to_unsigned(3520, 12), 1205 => to_unsigned(2796, 12), 1206 => to_unsigned(3968, 12), 1207 => to_unsigned(2999, 12), 1208 => to_unsigned(191, 12), 1209 => to_unsigned(33, 12), 1210 => to_unsigned(1671, 12), 1211 => to_unsigned(3227, 12), 1212 => to_unsigned(1494, 12), 1213 => to_unsigned(90, 12), 1214 => to_unsigned(1749, 12), 1215 => to_unsigned(1508, 12), 1216 => to_unsigned(1844, 12), 1217 => to_unsigned(3637, 12), 1218 => to_unsigned(3123, 12), 1219 => to_unsigned(89, 12), 1220 => to_unsigned(2267, 12), 1221 => to_unsigned(2825, 12), 1222 => to_unsigned(2617, 12), 1223 => to_unsigned(182, 12), 1224 => to_unsigned(688, 12), 1225 => to_unsigned(1437, 12), 1226 => to_unsigned(3418, 12), 1227 => to_unsigned(393, 12), 1228 => to_unsigned(3760, 12), 1229 => to_unsigned(925, 12), 1230 => to_unsigned(2932, 12), 1231 => to_unsigned(3755, 12), 1232 => to_unsigned(906, 12), 1233 => to_unsigned(3071, 12), 1234 => to_unsigned(2470, 12), 1235 => to_unsigned(3049, 12), 1236 => to_unsigned(2746, 12), 1237 => to_unsigned(1430, 12), 1238 => to_unsigned(1296, 12), 1239 => to_unsigned(3028, 12), 1240 => to_unsigned(3173, 12), 1241 => to_unsigned(2732, 12), 1242 => to_unsigned(2459, 12), 1243 => to_unsigned(266, 12), 1244 => to_unsigned(2413, 12), 1245 => to_unsigned(2215, 12), 1246 => to_unsigned(2093, 12), 1247 => to_unsigned(428, 12), 1248 => to_unsigned(4009, 12), 1249 => to_unsigned(3677, 12), 1250 => to_unsigned(635, 12), 1251 => to_unsigned(3069, 12), 1252 => to_unsigned(133, 12), 1253 => to_unsigned(2690, 12), 1254 => to_unsigned(304, 12), 1255 => to_unsigned(2578, 12), 1256 => to_unsigned(2020, 12), 1257 => to_unsigned(2150, 12), 1258 => to_unsigned(2655, 12), 1259 => to_unsigned(560, 12), 1260 => to_unsigned(823, 12), 1261 => to_unsigned(445, 12), 1262 => to_unsigned(2184, 12), 1263 => to_unsigned(3542, 12), 1264 => to_unsigned(934, 12), 1265 => to_unsigned(19, 12), 1266 => to_unsigned(762, 12), 1267 => to_unsigned(1111, 12), 1268 => to_unsigned(645, 12), 1269 => to_unsigned(3774, 12), 1270 => to_unsigned(1308, 12), 1271 => to_unsigned(1399, 12), 1272 => to_unsigned(801, 12), 1273 => to_unsigned(1729, 12), 1274 => to_unsigned(1082, 12), 1275 => to_unsigned(67, 12), 1276 => to_unsigned(1969, 12), 1277 => to_unsigned(3412, 12), 1278 => to_unsigned(2766, 12), 1279 => to_unsigned(134, 12), 1280 => to_unsigned(939, 12), 1281 => to_unsigned(2805, 12), 1282 => to_unsigned(2923, 12), 1283 => to_unsigned(828, 12), 1284 => to_unsigned(3739, 12), 1285 => to_unsigned(2194, 12), 1286 => to_unsigned(1629, 12), 1287 => to_unsigned(3249, 12), 1288 => to_unsigned(897, 12), 1289 => to_unsigned(3659, 12), 1290 => to_unsigned(2525, 12), 1291 => to_unsigned(438, 12), 1292 => to_unsigned(173, 12), 1293 => to_unsigned(1791, 12), 1294 => to_unsigned(375, 12), 1295 => to_unsigned(11, 12), 1296 => to_unsigned(3996, 12), 1297 => to_unsigned(3995, 12), 1298 => to_unsigned(2999, 12), 1299 => to_unsigned(534, 12), 1300 => to_unsigned(1178, 12), 1301 => to_unsigned(2933, 12), 1302 => to_unsigned(1699, 12), 1303 => to_unsigned(2414, 12), 1304 => to_unsigned(3158, 12), 1305 => to_unsigned(472, 12), 1306 => to_unsigned(2136, 12), 1307 => to_unsigned(1869, 12), 1308 => to_unsigned(3558, 12), 1309 => to_unsigned(3911, 12), 1310 => to_unsigned(1101, 12), 1311 => to_unsigned(2830, 12), 1312 => to_unsigned(2843, 12), 1313 => to_unsigned(1607, 12), 1314 => to_unsigned(341, 12), 1315 => to_unsigned(1396, 12), 1316 => to_unsigned(455, 12), 1317 => to_unsigned(1176, 12), 1318 => to_unsigned(303, 12), 1319 => to_unsigned(2517, 12), 1320 => to_unsigned(2170, 12), 1321 => to_unsigned(2521, 12), 1322 => to_unsigned(125, 12), 1323 => to_unsigned(115, 12), 1324 => to_unsigned(3877, 12), 1325 => to_unsigned(1968, 12), 1326 => to_unsigned(4041, 12), 1327 => to_unsigned(2874, 12), 1328 => to_unsigned(1588, 12), 1329 => to_unsigned(1415, 12), 1330 => to_unsigned(2561, 12), 1331 => to_unsigned(3755, 12), 1332 => to_unsigned(1913, 12), 1333 => to_unsigned(1155, 12), 1334 => to_unsigned(871, 12), 1335 => to_unsigned(31, 12), 1336 => to_unsigned(20, 12), 1337 => to_unsigned(469, 12), 1338 => to_unsigned(3600, 12), 1339 => to_unsigned(2380, 12), 1340 => to_unsigned(3387, 12), 1341 => to_unsigned(405, 12), 1342 => to_unsigned(2118, 12), 1343 => to_unsigned(375, 12), 1344 => to_unsigned(521, 12), 1345 => to_unsigned(1318, 12), 1346 => to_unsigned(3402, 12), 1347 => to_unsigned(3888, 12), 1348 => to_unsigned(798, 12), 1349 => to_unsigned(152, 12), 1350 => to_unsigned(169, 12), 1351 => to_unsigned(2098, 12), 1352 => to_unsigned(2120, 12), 1353 => to_unsigned(1519, 12), 1354 => to_unsigned(2855, 12), 1355 => to_unsigned(2170, 12), 1356 => to_unsigned(3265, 12), 1357 => to_unsigned(4043, 12), 1358 => to_unsigned(627, 12), 1359 => to_unsigned(1468, 12), 1360 => to_unsigned(3803, 12), 1361 => to_unsigned(744, 12), 1362 => to_unsigned(37, 12), 1363 => to_unsigned(3233, 12), 1364 => to_unsigned(2080, 12), 1365 => to_unsigned(2381, 12), 1366 => to_unsigned(2692, 12), 1367 => to_unsigned(2403, 12), 1368 => to_unsigned(817, 12), 1369 => to_unsigned(797, 12), 1370 => to_unsigned(129, 12), 1371 => to_unsigned(3262, 12), 1372 => to_unsigned(3637, 12), 1373 => to_unsigned(10, 12), 1374 => to_unsigned(1222, 12), 1375 => to_unsigned(2650, 12), 1376 => to_unsigned(41, 12), 1377 => to_unsigned(1531, 12), 1378 => to_unsigned(3870, 12), 1379 => to_unsigned(628, 12), 1380 => to_unsigned(1740, 12), 1381 => to_unsigned(2693, 12), 1382 => to_unsigned(3607, 12), 1383 => to_unsigned(3062, 12), 1384 => to_unsigned(2272, 12), 1385 => to_unsigned(2495, 12), 1386 => to_unsigned(928, 12), 1387 => to_unsigned(3653, 12), 1388 => to_unsigned(2274, 12), 1389 => to_unsigned(152, 12), 1390 => to_unsigned(1817, 12), 1391 => to_unsigned(3463, 12), 1392 => to_unsigned(2513, 12), 1393 => to_unsigned(984, 12), 1394 => to_unsigned(3534, 12), 1395 => to_unsigned(401, 12), 1396 => to_unsigned(820, 12), 1397 => to_unsigned(1669, 12), 1398 => to_unsigned(299, 12), 1399 => to_unsigned(929, 12), 1400 => to_unsigned(940, 12), 1401 => to_unsigned(3493, 12), 1402 => to_unsigned(660, 12), 1403 => to_unsigned(2789, 12), 1404 => to_unsigned(3457, 12), 1405 => to_unsigned(2572, 12), 1406 => to_unsigned(3365, 12), 1407 => to_unsigned(3947, 12), 1408 => to_unsigned(1232, 12), 1409 => to_unsigned(2222, 12), 1410 => to_unsigned(3690, 12), 1411 => to_unsigned(3300, 12), 1412 => to_unsigned(738, 12), 1413 => to_unsigned(1088, 12), 1414 => to_unsigned(419, 12), 1415 => to_unsigned(1202, 12), 1416 => to_unsigned(2446, 12), 1417 => to_unsigned(601, 12), 1418 => to_unsigned(3372, 12), 1419 => to_unsigned(46, 12), 1420 => to_unsigned(3717, 12), 1421 => to_unsigned(2877, 12), 1422 => to_unsigned(2076, 12), 1423 => to_unsigned(716, 12), 1424 => to_unsigned(176, 12), 1425 => to_unsigned(742, 12), 1426 => to_unsigned(2503, 12), 1427 => to_unsigned(1747, 12), 1428 => to_unsigned(1065, 12), 1429 => to_unsigned(469, 12), 1430 => to_unsigned(2216, 12), 1431 => to_unsigned(2303, 12), 1432 => to_unsigned(1049, 12), 1433 => to_unsigned(2880, 12), 1434 => to_unsigned(598, 12), 1435 => to_unsigned(2347, 12), 1436 => to_unsigned(3110, 12), 1437 => to_unsigned(1269, 12), 1438 => to_unsigned(3609, 12), 1439 => to_unsigned(383, 12), 1440 => to_unsigned(1592, 12), 1441 => to_unsigned(3500, 12), 1442 => to_unsigned(3548, 12), 1443 => to_unsigned(2817, 12), 1444 => to_unsigned(3266, 12), 1445 => to_unsigned(1462, 12), 1446 => to_unsigned(3210, 12), 1447 => to_unsigned(3821, 12), 1448 => to_unsigned(1901, 12), 1449 => to_unsigned(3254, 12), 1450 => to_unsigned(299, 12), 1451 => to_unsigned(3341, 12), 1452 => to_unsigned(988, 12), 1453 => to_unsigned(1773, 12), 1454 => to_unsigned(1025, 12), 1455 => to_unsigned(2815, 12), 1456 => to_unsigned(764, 12), 1457 => to_unsigned(2549, 12), 1458 => to_unsigned(3877, 12), 1459 => to_unsigned(2788, 12), 1460 => to_unsigned(2918, 12), 1461 => to_unsigned(1458, 12), 1462 => to_unsigned(633, 12), 1463 => to_unsigned(1506, 12), 1464 => to_unsigned(872, 12), 1465 => to_unsigned(296, 12), 1466 => to_unsigned(482, 12), 1467 => to_unsigned(1263, 12), 1468 => to_unsigned(1178, 12), 1469 => to_unsigned(3307, 12), 1470 => to_unsigned(2777, 12), 1471 => to_unsigned(601, 12), 1472 => to_unsigned(2617, 12), 1473 => to_unsigned(190, 12), 1474 => to_unsigned(2694, 12), 1475 => to_unsigned(2959, 12), 1476 => to_unsigned(1594, 12), 1477 => to_unsigned(1015, 12), 1478 => to_unsigned(1070, 12), 1479 => to_unsigned(3422, 12), 1480 => to_unsigned(3975, 12), 1481 => to_unsigned(3277, 12), 1482 => to_unsigned(3799, 12), 1483 => to_unsigned(3308, 12), 1484 => to_unsigned(2075, 12), 1485 => to_unsigned(842, 12), 1486 => to_unsigned(3002, 12), 1487 => to_unsigned(1444, 12), 1488 => to_unsigned(665, 12), 1489 => to_unsigned(2038, 12), 1490 => to_unsigned(334, 12), 1491 => to_unsigned(1761, 12), 1492 => to_unsigned(2936, 12), 1493 => to_unsigned(425, 12), 1494 => to_unsigned(3255, 12), 1495 => to_unsigned(999, 12), 1496 => to_unsigned(2918, 12), 1497 => to_unsigned(2847, 12), 1498 => to_unsigned(633, 12), 1499 => to_unsigned(1363, 12), 1500 => to_unsigned(3594, 12), 1501 => to_unsigned(3255, 12), 1502 => to_unsigned(1433, 12), 1503 => to_unsigned(4006, 12), 1504 => to_unsigned(2760, 12), 1505 => to_unsigned(2214, 12), 1506 => to_unsigned(1160, 12), 1507 => to_unsigned(2396, 12), 1508 => to_unsigned(1588, 12), 1509 => to_unsigned(2115, 12), 1510 => to_unsigned(1352, 12), 1511 => to_unsigned(3420, 12), 1512 => to_unsigned(938, 12), 1513 => to_unsigned(617, 12), 1514 => to_unsigned(3262, 12), 1515 => to_unsigned(910, 12), 1516 => to_unsigned(3345, 12), 1517 => to_unsigned(3049, 12), 1518 => to_unsigned(145, 12), 1519 => to_unsigned(650, 12), 1520 => to_unsigned(2756, 12), 1521 => to_unsigned(1919, 12), 1522 => to_unsigned(733, 12), 1523 => to_unsigned(1568, 12), 1524 => to_unsigned(1894, 12), 1525 => to_unsigned(3768, 12), 1526 => to_unsigned(483, 12), 1527 => to_unsigned(3149, 12), 1528 => to_unsigned(1693, 12), 1529 => to_unsigned(4030, 12), 1530 => to_unsigned(3283, 12), 1531 => to_unsigned(2284, 12), 1532 => to_unsigned(3083, 12), 1533 => to_unsigned(3749, 12), 1534 => to_unsigned(3427, 12), 1535 => to_unsigned(771, 12), 1536 => to_unsigned(1602, 12), 1537 => to_unsigned(122, 12), 1538 => to_unsigned(1297, 12), 1539 => to_unsigned(193, 12), 1540 => to_unsigned(2358, 12), 1541 => to_unsigned(1281, 12), 1542 => to_unsigned(4019, 12), 1543 => to_unsigned(1803, 12), 1544 => to_unsigned(925, 12), 1545 => to_unsigned(2178, 12), 1546 => to_unsigned(280, 12), 1547 => to_unsigned(3767, 12), 1548 => to_unsigned(2460, 12), 1549 => to_unsigned(285, 12), 1550 => to_unsigned(684, 12), 1551 => to_unsigned(3268, 12), 1552 => to_unsigned(2365, 12), 1553 => to_unsigned(1822, 12), 1554 => to_unsigned(1816, 12), 1555 => to_unsigned(2983, 12), 1556 => to_unsigned(3421, 12), 1557 => to_unsigned(3604, 12), 1558 => to_unsigned(3700, 12), 1559 => to_unsigned(854, 12), 1560 => to_unsigned(2967, 12), 1561 => to_unsigned(267, 12), 1562 => to_unsigned(4020, 12), 1563 => to_unsigned(3677, 12), 1564 => to_unsigned(396, 12), 1565 => to_unsigned(3822, 12), 1566 => to_unsigned(161, 12), 1567 => to_unsigned(3, 12), 1568 => to_unsigned(327, 12), 1569 => to_unsigned(1850, 12), 1570 => to_unsigned(171, 12), 1571 => to_unsigned(1381, 12), 1572 => to_unsigned(3980, 12), 1573 => to_unsigned(3096, 12), 1574 => to_unsigned(1265, 12), 1575 => to_unsigned(4058, 12), 1576 => to_unsigned(2805, 12), 1577 => to_unsigned(1039, 12), 1578 => to_unsigned(117, 12), 1579 => to_unsigned(3734, 12), 1580 => to_unsigned(483, 12), 1581 => to_unsigned(1377, 12), 1582 => to_unsigned(1914, 12), 1583 => to_unsigned(3664, 12), 1584 => to_unsigned(3692, 12), 1585 => to_unsigned(125, 12), 1586 => to_unsigned(1271, 12), 1587 => to_unsigned(3264, 12), 1588 => to_unsigned(2934, 12), 1589 => to_unsigned(196, 12), 1590 => to_unsigned(1542, 12), 1591 => to_unsigned(3506, 12), 1592 => to_unsigned(3449, 12), 1593 => to_unsigned(1950, 12), 1594 => to_unsigned(762, 12), 1595 => to_unsigned(1747, 12), 1596 => to_unsigned(528, 12), 1597 => to_unsigned(81, 12), 1598 => to_unsigned(3485, 12), 1599 => to_unsigned(365, 12), 1600 => to_unsigned(1612, 12), 1601 => to_unsigned(1354, 12), 1602 => to_unsigned(2449, 12), 1603 => to_unsigned(501, 12), 1604 => to_unsigned(1718, 12), 1605 => to_unsigned(994, 12), 1606 => to_unsigned(2856, 12), 1607 => to_unsigned(3544, 12), 1608 => to_unsigned(2075, 12), 1609 => to_unsigned(1570, 12), 1610 => to_unsigned(1466, 12), 1611 => to_unsigned(3854, 12), 1612 => to_unsigned(776, 12), 1613 => to_unsigned(2100, 12), 1614 => to_unsigned(3884, 12), 1615 => to_unsigned(2962, 12), 1616 => to_unsigned(475, 12), 1617 => to_unsigned(3290, 12), 1618 => to_unsigned(2034, 12), 1619 => to_unsigned(3799, 12), 1620 => to_unsigned(2503, 12), 1621 => to_unsigned(970, 12), 1622 => to_unsigned(1986, 12), 1623 => to_unsigned(1045, 12), 1624 => to_unsigned(2764, 12), 1625 => to_unsigned(3174, 12), 1626 => to_unsigned(395, 12), 1627 => to_unsigned(2710, 12), 1628 => to_unsigned(956, 12), 1629 => to_unsigned(3751, 12), 1630 => to_unsigned(3533, 12), 1631 => to_unsigned(4089, 12), 1632 => to_unsigned(289, 12), 1633 => to_unsigned(2025, 12), 1634 => to_unsigned(4056, 12), 1635 => to_unsigned(757, 12), 1636 => to_unsigned(251, 12), 1637 => to_unsigned(3767, 12), 1638 => to_unsigned(2519, 12), 1639 => to_unsigned(3671, 12), 1640 => to_unsigned(1244, 12), 1641 => to_unsigned(2318, 12), 1642 => to_unsigned(2013, 12), 1643 => to_unsigned(1213, 12), 1644 => to_unsigned(2475, 12), 1645 => to_unsigned(2215, 12), 1646 => to_unsigned(4033, 12), 1647 => to_unsigned(3420, 12), 1648 => to_unsigned(2805, 12), 1649 => to_unsigned(3504, 12), 1650 => to_unsigned(574, 12), 1651 => to_unsigned(3698, 12), 1652 => to_unsigned(1782, 12), 1653 => to_unsigned(3550, 12), 1654 => to_unsigned(1167, 12), 1655 => to_unsigned(3423, 12), 1656 => to_unsigned(2460, 12), 1657 => to_unsigned(264, 12), 1658 => to_unsigned(1380, 12), 1659 => to_unsigned(876, 12), 1660 => to_unsigned(467, 12), 1661 => to_unsigned(3599, 12), 1662 => to_unsigned(1014, 12), 1663 => to_unsigned(2130, 12), 1664 => to_unsigned(2921, 12), 1665 => to_unsigned(699, 12), 1666 => to_unsigned(2368, 12), 1667 => to_unsigned(2624, 12), 1668 => to_unsigned(567, 12), 1669 => to_unsigned(2737, 12), 1670 => to_unsigned(3389, 12), 1671 => to_unsigned(961, 12), 1672 => to_unsigned(1354, 12), 1673 => to_unsigned(222, 12), 1674 => to_unsigned(2954, 12), 1675 => to_unsigned(3491, 12), 1676 => to_unsigned(3586, 12), 1677 => to_unsigned(1793, 12), 1678 => to_unsigned(1481, 12), 1679 => to_unsigned(3062, 12), 1680 => to_unsigned(1962, 12), 1681 => to_unsigned(1136, 12), 1682 => to_unsigned(1908, 12), 1683 => to_unsigned(2499, 12), 1684 => to_unsigned(2542, 12), 1685 => to_unsigned(2411, 12), 1686 => to_unsigned(3108, 12), 1687 => to_unsigned(525, 12), 1688 => to_unsigned(2211, 12), 1689 => to_unsigned(245, 12), 1690 => to_unsigned(3855, 12), 1691 => to_unsigned(3762, 12), 1692 => to_unsigned(878, 12), 1693 => to_unsigned(3017, 12), 1694 => to_unsigned(871, 12), 1695 => to_unsigned(2002, 12), 1696 => to_unsigned(3010, 12), 1697 => to_unsigned(4013, 12), 1698 => to_unsigned(3625, 12), 1699 => to_unsigned(4, 12), 1700 => to_unsigned(2812, 12), 1701 => to_unsigned(2156, 12), 1702 => to_unsigned(3534, 12), 1703 => to_unsigned(1935, 12), 1704 => to_unsigned(1132, 12), 1705 => to_unsigned(2004, 12), 1706 => to_unsigned(1497, 12), 1707 => to_unsigned(3626, 12), 1708 => to_unsigned(3026, 12), 1709 => to_unsigned(3926, 12), 1710 => to_unsigned(2964, 12), 1711 => to_unsigned(3454, 12), 1712 => to_unsigned(1515, 12), 1713 => to_unsigned(2933, 12), 1714 => to_unsigned(2350, 12), 1715 => to_unsigned(2876, 12), 1716 => to_unsigned(1002, 12), 1717 => to_unsigned(818, 12), 1718 => to_unsigned(1474, 12), 1719 => to_unsigned(3015, 12), 1720 => to_unsigned(4016, 12), 1721 => to_unsigned(2962, 12), 1722 => to_unsigned(2125, 12), 1723 => to_unsigned(1345, 12), 1724 => to_unsigned(3379, 12), 1725 => to_unsigned(1396, 12), 1726 => to_unsigned(1632, 12), 1727 => to_unsigned(2499, 12), 1728 => to_unsigned(2038, 12), 1729 => to_unsigned(1892, 12), 1730 => to_unsigned(2224, 12), 1731 => to_unsigned(3056, 12), 1732 => to_unsigned(2589, 12), 1733 => to_unsigned(2115, 12), 1734 => to_unsigned(1605, 12), 1735 => to_unsigned(1691, 12), 1736 => to_unsigned(2442, 12), 1737 => to_unsigned(1076, 12), 1738 => to_unsigned(2286, 12), 1739 => to_unsigned(2822, 12), 1740 => to_unsigned(3852, 12), 1741 => to_unsigned(321, 12), 1742 => to_unsigned(1347, 12), 1743 => to_unsigned(703, 12), 1744 => to_unsigned(3080, 12), 1745 => to_unsigned(1380, 12), 1746 => to_unsigned(395, 12), 1747 => to_unsigned(465, 12), 1748 => to_unsigned(872, 12), 1749 => to_unsigned(34, 12), 1750 => to_unsigned(1283, 12), 1751 => to_unsigned(3745, 12), 1752 => to_unsigned(1683, 12), 1753 => to_unsigned(643, 12), 1754 => to_unsigned(1261, 12), 1755 => to_unsigned(2141, 12), 1756 => to_unsigned(1306, 12), 1757 => to_unsigned(731, 12), 1758 => to_unsigned(2407, 12), 1759 => to_unsigned(1523, 12), 1760 => to_unsigned(4080, 12), 1761 => to_unsigned(2885, 12), 1762 => to_unsigned(3734, 12), 1763 => to_unsigned(2516, 12), 1764 => to_unsigned(3661, 12), 1765 => to_unsigned(3290, 12), 1766 => to_unsigned(2975, 12), 1767 => to_unsigned(3314, 12), 1768 => to_unsigned(1062, 12), 1769 => to_unsigned(901, 12), 1770 => to_unsigned(689, 12), 1771 => to_unsigned(3814, 12), 1772 => to_unsigned(2185, 12), 1773 => to_unsigned(231, 12), 1774 => to_unsigned(3421, 12), 1775 => to_unsigned(1900, 12), 1776 => to_unsigned(3256, 12), 1777 => to_unsigned(3261, 12), 1778 => to_unsigned(2696, 12), 1779 => to_unsigned(3040, 12), 1780 => to_unsigned(946, 12), 1781 => to_unsigned(1680, 12), 1782 => to_unsigned(2453, 12), 1783 => to_unsigned(735, 12), 1784 => to_unsigned(3179, 12), 1785 => to_unsigned(504, 12), 1786 => to_unsigned(248, 12), 1787 => to_unsigned(2986, 12), 1788 => to_unsigned(3013, 12), 1789 => to_unsigned(2290, 12), 1790 => to_unsigned(131, 12), 1791 => to_unsigned(59, 12), 1792 => to_unsigned(3160, 12), 1793 => to_unsigned(3550, 12), 1794 => to_unsigned(11, 12), 1795 => to_unsigned(3705, 12), 1796 => to_unsigned(3820, 12), 1797 => to_unsigned(2473, 12), 1798 => to_unsigned(2595, 12), 1799 => to_unsigned(3319, 12), 1800 => to_unsigned(538, 12), 1801 => to_unsigned(3699, 12), 1802 => to_unsigned(3248, 12), 1803 => to_unsigned(130, 12), 1804 => to_unsigned(390, 12), 1805 => to_unsigned(3377, 12), 1806 => to_unsigned(2671, 12), 1807 => to_unsigned(1035, 12), 1808 => to_unsigned(1066, 12), 1809 => to_unsigned(2581, 12), 1810 => to_unsigned(126, 12), 1811 => to_unsigned(3861, 12), 1812 => to_unsigned(2128, 12), 1813 => to_unsigned(3848, 12), 1814 => to_unsigned(2263, 12), 1815 => to_unsigned(2919, 12), 1816 => to_unsigned(3056, 12), 1817 => to_unsigned(3797, 12), 1818 => to_unsigned(3008, 12), 1819 => to_unsigned(3557, 12), 1820 => to_unsigned(2287, 12), 1821 => to_unsigned(523, 12), 1822 => to_unsigned(675, 12), 1823 => to_unsigned(3810, 12), 1824 => to_unsigned(2394, 12), 1825 => to_unsigned(544, 12), 1826 => to_unsigned(2145, 12), 1827 => to_unsigned(2155, 12), 1828 => to_unsigned(2812, 12), 1829 => to_unsigned(1494, 12), 1830 => to_unsigned(2451, 12), 1831 => to_unsigned(1000, 12), 1832 => to_unsigned(3558, 12), 1833 => to_unsigned(3637, 12), 1834 => to_unsigned(2792, 12), 1835 => to_unsigned(56, 12), 1836 => to_unsigned(1533, 12), 1837 => to_unsigned(3773, 12), 1838 => to_unsigned(1465, 12), 1839 => to_unsigned(1090, 12), 1840 => to_unsigned(3676, 12), 1841 => to_unsigned(2592, 12), 1842 => to_unsigned(1287, 12), 1843 => to_unsigned(1277, 12), 1844 => to_unsigned(2703, 12), 1845 => to_unsigned(619, 12), 1846 => to_unsigned(3935, 12), 1847 => to_unsigned(3057, 12), 1848 => to_unsigned(3806, 12), 1849 => to_unsigned(3500, 12), 1850 => to_unsigned(2517, 12), 1851 => to_unsigned(2257, 12), 1852 => to_unsigned(205, 12), 1853 => to_unsigned(2530, 12), 1854 => to_unsigned(2864, 12), 1855 => to_unsigned(987, 12), 1856 => to_unsigned(2248, 12), 1857 => to_unsigned(3748, 12), 1858 => to_unsigned(468, 12), 1859 => to_unsigned(2660, 12), 1860 => to_unsigned(2714, 12), 1861 => to_unsigned(823, 12), 1862 => to_unsigned(3109, 12), 1863 => to_unsigned(3250, 12), 1864 => to_unsigned(3692, 12), 1865 => to_unsigned(2722, 12), 1866 => to_unsigned(2058, 12), 1867 => to_unsigned(1759, 12), 1868 => to_unsigned(1364, 12), 1869 => to_unsigned(1807, 12), 1870 => to_unsigned(2923, 12), 1871 => to_unsigned(1069, 12), 1872 => to_unsigned(889, 12), 1873 => to_unsigned(2730, 12), 1874 => to_unsigned(279, 12), 1875 => to_unsigned(1468, 12), 1876 => to_unsigned(4014, 12), 1877 => to_unsigned(779, 12), 1878 => to_unsigned(3989, 12), 1879 => to_unsigned(3594, 12), 1880 => to_unsigned(3009, 12), 1881 => to_unsigned(579, 12), 1882 => to_unsigned(307, 12), 1883 => to_unsigned(1913, 12), 1884 => to_unsigned(1316, 12), 1885 => to_unsigned(2353, 12), 1886 => to_unsigned(481, 12), 1887 => to_unsigned(1916, 12), 1888 => to_unsigned(3524, 12), 1889 => to_unsigned(2760, 12), 1890 => to_unsigned(323, 12), 1891 => to_unsigned(867, 12), 1892 => to_unsigned(847, 12), 1893 => to_unsigned(820, 12), 1894 => to_unsigned(1374, 12), 1895 => to_unsigned(168, 12), 1896 => to_unsigned(895, 12), 1897 => to_unsigned(1873, 12), 1898 => to_unsigned(801, 12), 1899 => to_unsigned(530, 12), 1900 => to_unsigned(639, 12), 1901 => to_unsigned(1347, 12), 1902 => to_unsigned(1017, 12), 1903 => to_unsigned(3605, 12), 1904 => to_unsigned(1720, 12), 1905 => to_unsigned(2611, 12), 1906 => to_unsigned(3572, 12), 1907 => to_unsigned(3309, 12), 1908 => to_unsigned(726, 12), 1909 => to_unsigned(464, 12), 1910 => to_unsigned(1742, 12), 1911 => to_unsigned(729, 12), 1912 => to_unsigned(525, 12), 1913 => to_unsigned(1411, 12), 1914 => to_unsigned(985, 12), 1915 => to_unsigned(1786, 12), 1916 => to_unsigned(3537, 12), 1917 => to_unsigned(1484, 12), 1918 => to_unsigned(2077, 12), 1919 => to_unsigned(2734, 12), 1920 => to_unsigned(2221, 12), 1921 => to_unsigned(217, 12), 1922 => to_unsigned(2373, 12), 1923 => to_unsigned(492, 12), 1924 => to_unsigned(2568, 12), 1925 => to_unsigned(2990, 12), 1926 => to_unsigned(249, 12), 1927 => to_unsigned(2224, 12), 1928 => to_unsigned(3322, 12), 1929 => to_unsigned(3776, 12), 1930 => to_unsigned(2114, 12), 1931 => to_unsigned(1085, 12), 1932 => to_unsigned(393, 12), 1933 => to_unsigned(11, 12), 1934 => to_unsigned(3391, 12), 1935 => to_unsigned(1823, 12), 1936 => to_unsigned(3990, 12), 1937 => to_unsigned(1825, 12), 1938 => to_unsigned(2495, 12), 1939 => to_unsigned(2991, 12), 1940 => to_unsigned(2132, 12), 1941 => to_unsigned(713, 12), 1942 => to_unsigned(3926, 12), 1943 => to_unsigned(3419, 12), 1944 => to_unsigned(1353, 12), 1945 => to_unsigned(147, 12), 1946 => to_unsigned(2007, 12), 1947 => to_unsigned(185, 12), 1948 => to_unsigned(2999, 12), 1949 => to_unsigned(1844, 12), 1950 => to_unsigned(1276, 12), 1951 => to_unsigned(3032, 12), 1952 => to_unsigned(372, 12), 1953 => to_unsigned(1241, 12), 1954 => to_unsigned(2674, 12), 1955 => to_unsigned(198, 12), 1956 => to_unsigned(819, 12), 1957 => to_unsigned(3363, 12), 1958 => to_unsigned(2640, 12), 1959 => to_unsigned(479, 12), 1960 => to_unsigned(1569, 12), 1961 => to_unsigned(3461, 12), 1962 => to_unsigned(700, 12), 1963 => to_unsigned(1933, 12), 1964 => to_unsigned(2315, 12), 1965 => to_unsigned(1387, 12), 1966 => to_unsigned(2731, 12), 1967 => to_unsigned(4037, 12), 1968 => to_unsigned(2506, 12), 1969 => to_unsigned(210, 12), 1970 => to_unsigned(3906, 12), 1971 => to_unsigned(3774, 12), 1972 => to_unsigned(119, 12), 1973 => to_unsigned(2704, 12), 1974 => to_unsigned(3328, 12), 1975 => to_unsigned(1293, 12), 1976 => to_unsigned(1072, 12), 1977 => to_unsigned(918, 12), 1978 => to_unsigned(2977, 12), 1979 => to_unsigned(3840, 12), 1980 => to_unsigned(3562, 12), 1981 => to_unsigned(585, 12), 1982 => to_unsigned(2713, 12), 1983 => to_unsigned(2152, 12), 1984 => to_unsigned(3385, 12), 1985 => to_unsigned(2618, 12), 1986 => to_unsigned(450, 12), 1987 => to_unsigned(3598, 12), 1988 => to_unsigned(3446, 12), 1989 => to_unsigned(3898, 12), 1990 => to_unsigned(3996, 12), 1991 => to_unsigned(2773, 12), 1992 => to_unsigned(1986, 12), 1993 => to_unsigned(2454, 12), 1994 => to_unsigned(509, 12), 1995 => to_unsigned(2248, 12), 1996 => to_unsigned(239, 12), 1997 => to_unsigned(464, 12), 1998 => to_unsigned(1315, 12), 1999 => to_unsigned(2541, 12), 2000 => to_unsigned(3995, 12), 2001 => to_unsigned(1890, 12), 2002 => to_unsigned(2361, 12), 2003 => to_unsigned(2695, 12), 2004 => to_unsigned(2973, 12), 2005 => to_unsigned(2442, 12), 2006 => to_unsigned(1629, 12), 2007 => to_unsigned(1095, 12), 2008 => to_unsigned(2544, 12), 2009 => to_unsigned(3207, 12), 2010 => to_unsigned(2881, 12), 2011 => to_unsigned(2457, 12), 2012 => to_unsigned(3981, 12), 2013 => to_unsigned(2253, 12), 2014 => to_unsigned(2240, 12), 2015 => to_unsigned(3881, 12), 2016 => to_unsigned(3756, 12), 2017 => to_unsigned(3219, 12), 2018 => to_unsigned(2371, 12), 2019 => to_unsigned(3961, 12), 2020 => to_unsigned(2215, 12), 2021 => to_unsigned(2165, 12), 2022 => to_unsigned(2369, 12), 2023 => to_unsigned(81, 12), 2024 => to_unsigned(3131, 12), 2025 => to_unsigned(1270, 12), 2026 => to_unsigned(1762, 12), 2027 => to_unsigned(2154, 12), 2028 => to_unsigned(1285, 12), 2029 => to_unsigned(2882, 12), 2030 => to_unsigned(2891, 12), 2031 => to_unsigned(1087, 12), 2032 => to_unsigned(2795, 12), 2033 => to_unsigned(3013, 12), 2034 => to_unsigned(458, 12), 2035 => to_unsigned(2036, 12), 2036 => to_unsigned(1668, 12), 2037 => to_unsigned(301, 12), 2038 => to_unsigned(2431, 12), 2039 => to_unsigned(3360, 12), 2040 => to_unsigned(3380, 12), 2041 => to_unsigned(4016, 12), 2042 => to_unsigned(3795, 12), 2043 => to_unsigned(342, 12), 2044 => to_unsigned(3140, 12), 2045 => to_unsigned(2453, 12), 2046 => to_unsigned(3043, 12), 2047 => to_unsigned(460, 12)),
            1 => (0 => to_unsigned(671, 12), 1 => to_unsigned(3424, 12), 2 => to_unsigned(2779, 12), 3 => to_unsigned(2621, 12), 4 => to_unsigned(2765, 12), 5 => to_unsigned(1694, 12), 6 => to_unsigned(1106, 12), 7 => to_unsigned(1355, 12), 8 => to_unsigned(3040, 12), 9 => to_unsigned(2742, 12), 10 => to_unsigned(1394, 12), 11 => to_unsigned(779, 12), 12 => to_unsigned(82, 12), 13 => to_unsigned(369, 12), 14 => to_unsigned(2160, 12), 15 => to_unsigned(732, 12), 16 => to_unsigned(1515, 12), 17 => to_unsigned(530, 12), 18 => to_unsigned(3285, 12), 19 => to_unsigned(3523, 12), 20 => to_unsigned(1949, 12), 21 => to_unsigned(3617, 12), 22 => to_unsigned(2989, 12), 23 => to_unsigned(3704, 12), 24 => to_unsigned(3114, 12), 25 => to_unsigned(3293, 12), 26 => to_unsigned(1739, 12), 27 => to_unsigned(2003, 12), 28 => to_unsigned(2035, 12), 29 => to_unsigned(2104, 12), 30 => to_unsigned(3026, 12), 31 => to_unsigned(35, 12), 32 => to_unsigned(2221, 12), 33 => to_unsigned(486, 12), 34 => to_unsigned(3759, 12), 35 => to_unsigned(770, 12), 36 => to_unsigned(2691, 12), 37 => to_unsigned(1082, 12), 38 => to_unsigned(2947, 12), 39 => to_unsigned(2004, 12), 40 => to_unsigned(166, 12), 41 => to_unsigned(3344, 12), 42 => to_unsigned(3679, 12), 43 => to_unsigned(2189, 12), 44 => to_unsigned(3567, 12), 45 => to_unsigned(2827, 12), 46 => to_unsigned(3553, 12), 47 => to_unsigned(2781, 12), 48 => to_unsigned(594, 12), 49 => to_unsigned(3914, 12), 50 => to_unsigned(109, 12), 51 => to_unsigned(2136, 12), 52 => to_unsigned(2416, 12), 53 => to_unsigned(3988, 12), 54 => to_unsigned(3778, 12), 55 => to_unsigned(1105, 12), 56 => to_unsigned(3402, 12), 57 => to_unsigned(3228, 12), 58 => to_unsigned(732, 12), 59 => to_unsigned(3827, 12), 60 => to_unsigned(1125, 12), 61 => to_unsigned(3017, 12), 62 => to_unsigned(132, 12), 63 => to_unsigned(975, 12), 64 => to_unsigned(3511, 12), 65 => to_unsigned(3804, 12), 66 => to_unsigned(684, 12), 67 => to_unsigned(2316, 12), 68 => to_unsigned(1218, 12), 69 => to_unsigned(3167, 12), 70 => to_unsigned(1704, 12), 71 => to_unsigned(2367, 12), 72 => to_unsigned(1140, 12), 73 => to_unsigned(1595, 12), 74 => to_unsigned(2530, 12), 75 => to_unsigned(401, 12), 76 => to_unsigned(3144, 12), 77 => to_unsigned(2402, 12), 78 => to_unsigned(1694, 12), 79 => to_unsigned(456, 12), 80 => to_unsigned(1422, 12), 81 => to_unsigned(25, 12), 82 => to_unsigned(1549, 12), 83 => to_unsigned(3497, 12), 84 => to_unsigned(278, 12), 85 => to_unsigned(356, 12), 86 => to_unsigned(740, 12), 87 => to_unsigned(2129, 12), 88 => to_unsigned(3780, 12), 89 => to_unsigned(1536, 12), 90 => to_unsigned(3606, 12), 91 => to_unsigned(1444, 12), 92 => to_unsigned(2913, 12), 93 => to_unsigned(1419, 12), 94 => to_unsigned(2940, 12), 95 => to_unsigned(3636, 12), 96 => to_unsigned(2166, 12), 97 => to_unsigned(1668, 12), 98 => to_unsigned(3570, 12), 99 => to_unsigned(3052, 12), 100 => to_unsigned(3399, 12), 101 => to_unsigned(1730, 12), 102 => to_unsigned(76, 12), 103 => to_unsigned(3839, 12), 104 => to_unsigned(2191, 12), 105 => to_unsigned(1816, 12), 106 => to_unsigned(1026, 12), 107 => to_unsigned(3169, 12), 108 => to_unsigned(2555, 12), 109 => to_unsigned(2769, 12), 110 => to_unsigned(112, 12), 111 => to_unsigned(1059, 12), 112 => to_unsigned(270, 12), 113 => to_unsigned(1275, 12), 114 => to_unsigned(458, 12), 115 => to_unsigned(2865, 12), 116 => to_unsigned(2997, 12), 117 => to_unsigned(4074, 12), 118 => to_unsigned(1647, 12), 119 => to_unsigned(1022, 12), 120 => to_unsigned(2224, 12), 121 => to_unsigned(3304, 12), 122 => to_unsigned(1095, 12), 123 => to_unsigned(3146, 12), 124 => to_unsigned(1021, 12), 125 => to_unsigned(2109, 12), 126 => to_unsigned(671, 12), 127 => to_unsigned(2255, 12), 128 => to_unsigned(4056, 12), 129 => to_unsigned(1809, 12), 130 => to_unsigned(758, 12), 131 => to_unsigned(2619, 12), 132 => to_unsigned(656, 12), 133 => to_unsigned(856, 12), 134 => to_unsigned(2390, 12), 135 => to_unsigned(2988, 12), 136 => to_unsigned(1866, 12), 137 => to_unsigned(2278, 12), 138 => to_unsigned(277, 12), 139 => to_unsigned(2809, 12), 140 => to_unsigned(823, 12), 141 => to_unsigned(1856, 12), 142 => to_unsigned(1222, 12), 143 => to_unsigned(1263, 12), 144 => to_unsigned(500, 12), 145 => to_unsigned(1082, 12), 146 => to_unsigned(3504, 12), 147 => to_unsigned(1459, 12), 148 => to_unsigned(3804, 12), 149 => to_unsigned(3664, 12), 150 => to_unsigned(1203, 12), 151 => to_unsigned(3261, 12), 152 => to_unsigned(1287, 12), 153 => to_unsigned(2030, 12), 154 => to_unsigned(3269, 12), 155 => to_unsigned(2689, 12), 156 => to_unsigned(1536, 12), 157 => to_unsigned(2787, 12), 158 => to_unsigned(1989, 12), 159 => to_unsigned(1035, 12), 160 => to_unsigned(3015, 12), 161 => to_unsigned(112, 12), 162 => to_unsigned(1858, 12), 163 => to_unsigned(563, 12), 164 => to_unsigned(1855, 12), 165 => to_unsigned(1873, 12), 166 => to_unsigned(609, 12), 167 => to_unsigned(2556, 12), 168 => to_unsigned(2479, 12), 169 => to_unsigned(715, 12), 170 => to_unsigned(567, 12), 171 => to_unsigned(236, 12), 172 => to_unsigned(2355, 12), 173 => to_unsigned(847, 12), 174 => to_unsigned(417, 12), 175 => to_unsigned(2268, 12), 176 => to_unsigned(3636, 12), 177 => to_unsigned(107, 12), 178 => to_unsigned(2582, 12), 179 => to_unsigned(2677, 12), 180 => to_unsigned(2958, 12), 181 => to_unsigned(2052, 12), 182 => to_unsigned(2399, 12), 183 => to_unsigned(3366, 12), 184 => to_unsigned(429, 12), 185 => to_unsigned(3425, 12), 186 => to_unsigned(839, 12), 187 => to_unsigned(3965, 12), 188 => to_unsigned(1764, 12), 189 => to_unsigned(2756, 12), 190 => to_unsigned(2292, 12), 191 => to_unsigned(2406, 12), 192 => to_unsigned(2169, 12), 193 => to_unsigned(2602, 12), 194 => to_unsigned(1181, 12), 195 => to_unsigned(3839, 12), 196 => to_unsigned(3572, 12), 197 => to_unsigned(59, 12), 198 => to_unsigned(3977, 12), 199 => to_unsigned(3295, 12), 200 => to_unsigned(3508, 12), 201 => to_unsigned(2101, 12), 202 => to_unsigned(1385, 12), 203 => to_unsigned(262, 12), 204 => to_unsigned(3688, 12), 205 => to_unsigned(1895, 12), 206 => to_unsigned(2710, 12), 207 => to_unsigned(3698, 12), 208 => to_unsigned(2832, 12), 209 => to_unsigned(1372, 12), 210 => to_unsigned(1551, 12), 211 => to_unsigned(2086, 12), 212 => to_unsigned(905, 12), 213 => to_unsigned(2716, 12), 214 => to_unsigned(1332, 12), 215 => to_unsigned(909, 12), 216 => to_unsigned(2375, 12), 217 => to_unsigned(55, 12), 218 => to_unsigned(2614, 12), 219 => to_unsigned(3115, 12), 220 => to_unsigned(1210, 12), 221 => to_unsigned(2007, 12), 222 => to_unsigned(1899, 12), 223 => to_unsigned(1206, 12), 224 => to_unsigned(1642, 12), 225 => to_unsigned(1905, 12), 226 => to_unsigned(1402, 12), 227 => to_unsigned(1490, 12), 228 => to_unsigned(1147, 12), 229 => to_unsigned(3702, 12), 230 => to_unsigned(2113, 12), 231 => to_unsigned(3551, 12), 232 => to_unsigned(3429, 12), 233 => to_unsigned(1330, 12), 234 => to_unsigned(3162, 12), 235 => to_unsigned(2864, 12), 236 => to_unsigned(234, 12), 237 => to_unsigned(3556, 12), 238 => to_unsigned(3500, 12), 239 => to_unsigned(157, 12), 240 => to_unsigned(3819, 12), 241 => to_unsigned(2978, 12), 242 => to_unsigned(1633, 12), 243 => to_unsigned(109, 12), 244 => to_unsigned(3856, 12), 245 => to_unsigned(485, 12), 246 => to_unsigned(2141, 12), 247 => to_unsigned(2944, 12), 248 => to_unsigned(3587, 12), 249 => to_unsigned(3635, 12), 250 => to_unsigned(1234, 12), 251 => to_unsigned(2699, 12), 252 => to_unsigned(2405, 12), 253 => to_unsigned(1477, 12), 254 => to_unsigned(3680, 12), 255 => to_unsigned(2024, 12), 256 => to_unsigned(3948, 12), 257 => to_unsigned(2979, 12), 258 => to_unsigned(3451, 12), 259 => to_unsigned(2405, 12), 260 => to_unsigned(581, 12), 261 => to_unsigned(2856, 12), 262 => to_unsigned(3762, 12), 263 => to_unsigned(1240, 12), 264 => to_unsigned(3146, 12), 265 => to_unsigned(1770, 12), 266 => to_unsigned(1483, 12), 267 => to_unsigned(3443, 12), 268 => to_unsigned(4031, 12), 269 => to_unsigned(3170, 12), 270 => to_unsigned(2548, 12), 271 => to_unsigned(1433, 12), 272 => to_unsigned(233, 12), 273 => to_unsigned(2213, 12), 274 => to_unsigned(1251, 12), 275 => to_unsigned(2075, 12), 276 => to_unsigned(1733, 12), 277 => to_unsigned(238, 12), 278 => to_unsigned(3811, 12), 279 => to_unsigned(3915, 12), 280 => to_unsigned(3942, 12), 281 => to_unsigned(2130, 12), 282 => to_unsigned(3003, 12), 283 => to_unsigned(2063, 12), 284 => to_unsigned(886, 12), 285 => to_unsigned(602, 12), 286 => to_unsigned(1034, 12), 287 => to_unsigned(524, 12), 288 => to_unsigned(592, 12), 289 => to_unsigned(2659, 12), 290 => to_unsigned(606, 12), 291 => to_unsigned(3117, 12), 292 => to_unsigned(896, 12), 293 => to_unsigned(3530, 12), 294 => to_unsigned(3204, 12), 295 => to_unsigned(2432, 12), 296 => to_unsigned(76, 12), 297 => to_unsigned(1714, 12), 298 => to_unsigned(2045, 12), 299 => to_unsigned(949, 12), 300 => to_unsigned(2431, 12), 301 => to_unsigned(1519, 12), 302 => to_unsigned(3275, 12), 303 => to_unsigned(1352, 12), 304 => to_unsigned(4043, 12), 305 => to_unsigned(1184, 12), 306 => to_unsigned(1055, 12), 307 => to_unsigned(1917, 12), 308 => to_unsigned(2831, 12), 309 => to_unsigned(1831, 12), 310 => to_unsigned(2261, 12), 311 => to_unsigned(3310, 12), 312 => to_unsigned(1074, 12), 313 => to_unsigned(123, 12), 314 => to_unsigned(3725, 12), 315 => to_unsigned(1552, 12), 316 => to_unsigned(3803, 12), 317 => to_unsigned(3790, 12), 318 => to_unsigned(519, 12), 319 => to_unsigned(1555, 12), 320 => to_unsigned(3878, 12), 321 => to_unsigned(1267, 12), 322 => to_unsigned(190, 12), 323 => to_unsigned(1843, 12), 324 => to_unsigned(761, 12), 325 => to_unsigned(2949, 12), 326 => to_unsigned(3161, 12), 327 => to_unsigned(3414, 12), 328 => to_unsigned(1860, 12), 329 => to_unsigned(3614, 12), 330 => to_unsigned(3871, 12), 331 => to_unsigned(2904, 12), 332 => to_unsigned(2182, 12), 333 => to_unsigned(900, 12), 334 => to_unsigned(3649, 12), 335 => to_unsigned(585, 12), 336 => to_unsigned(3564, 12), 337 => to_unsigned(3024, 12), 338 => to_unsigned(2500, 12), 339 => to_unsigned(3780, 12), 340 => to_unsigned(2944, 12), 341 => to_unsigned(2070, 12), 342 => to_unsigned(908, 12), 343 => to_unsigned(402, 12), 344 => to_unsigned(1635, 12), 345 => to_unsigned(3086, 12), 346 => to_unsigned(2413, 12), 347 => to_unsigned(3885, 12), 348 => to_unsigned(3029, 12), 349 => to_unsigned(1062, 12), 350 => to_unsigned(2057, 12), 351 => to_unsigned(3699, 12), 352 => to_unsigned(2857, 12), 353 => to_unsigned(688, 12), 354 => to_unsigned(1525, 12), 355 => to_unsigned(835, 12), 356 => to_unsigned(1549, 12), 357 => to_unsigned(3575, 12), 358 => to_unsigned(2894, 12), 359 => to_unsigned(1591, 12), 360 => to_unsigned(135, 12), 361 => to_unsigned(1465, 12), 362 => to_unsigned(793, 12), 363 => to_unsigned(2534, 12), 364 => to_unsigned(185, 12), 365 => to_unsigned(1039, 12), 366 => to_unsigned(3706, 12), 367 => to_unsigned(1510, 12), 368 => to_unsigned(3328, 12), 369 => to_unsigned(3748, 12), 370 => to_unsigned(1859, 12), 371 => to_unsigned(1526, 12), 372 => to_unsigned(2920, 12), 373 => to_unsigned(3747, 12), 374 => to_unsigned(714, 12), 375 => to_unsigned(1285, 12), 376 => to_unsigned(3020, 12), 377 => to_unsigned(542, 12), 378 => to_unsigned(3188, 12), 379 => to_unsigned(3433, 12), 380 => to_unsigned(1219, 12), 381 => to_unsigned(3691, 12), 382 => to_unsigned(690, 12), 383 => to_unsigned(4025, 12), 384 => to_unsigned(847, 12), 385 => to_unsigned(334, 12), 386 => to_unsigned(561, 12), 387 => to_unsigned(3371, 12), 388 => to_unsigned(3383, 12), 389 => to_unsigned(3392, 12), 390 => to_unsigned(1773, 12), 391 => to_unsigned(3987, 12), 392 => to_unsigned(1563, 12), 393 => to_unsigned(1783, 12), 394 => to_unsigned(216, 12), 395 => to_unsigned(1139, 12), 396 => to_unsigned(3312, 12), 397 => to_unsigned(954, 12), 398 => to_unsigned(2280, 12), 399 => to_unsigned(3368, 12), 400 => to_unsigned(765, 12), 401 => to_unsigned(3981, 12), 402 => to_unsigned(2836, 12), 403 => to_unsigned(3351, 12), 404 => to_unsigned(3985, 12), 405 => to_unsigned(3959, 12), 406 => to_unsigned(1535, 12), 407 => to_unsigned(1825, 12), 408 => to_unsigned(3346, 12), 409 => to_unsigned(36, 12), 410 => to_unsigned(743, 12), 411 => to_unsigned(3130, 12), 412 => to_unsigned(105, 12), 413 => to_unsigned(2142, 12), 414 => to_unsigned(2, 12), 415 => to_unsigned(35, 12), 416 => to_unsigned(1828, 12), 417 => to_unsigned(1847, 12), 418 => to_unsigned(2707, 12), 419 => to_unsigned(2184, 12), 420 => to_unsigned(754, 12), 421 => to_unsigned(23, 12), 422 => to_unsigned(2091, 12), 423 => to_unsigned(386, 12), 424 => to_unsigned(1159, 12), 425 => to_unsigned(1044, 12), 426 => to_unsigned(1266, 12), 427 => to_unsigned(2311, 12), 428 => to_unsigned(2803, 12), 429 => to_unsigned(1912, 12), 430 => to_unsigned(2687, 12), 431 => to_unsigned(1208, 12), 432 => to_unsigned(2224, 12), 433 => to_unsigned(3835, 12), 434 => to_unsigned(2442, 12), 435 => to_unsigned(1334, 12), 436 => to_unsigned(848, 12), 437 => to_unsigned(3838, 12), 438 => to_unsigned(2240, 12), 439 => to_unsigned(1731, 12), 440 => to_unsigned(1319, 12), 441 => to_unsigned(3791, 12), 442 => to_unsigned(415, 12), 443 => to_unsigned(3136, 12), 444 => to_unsigned(2878, 12), 445 => to_unsigned(106, 12), 446 => to_unsigned(360, 12), 447 => to_unsigned(3371, 12), 448 => to_unsigned(1001, 12), 449 => to_unsigned(815, 12), 450 => to_unsigned(1189, 12), 451 => to_unsigned(2636, 12), 452 => to_unsigned(404, 12), 453 => to_unsigned(3498, 12), 454 => to_unsigned(1376, 12), 455 => to_unsigned(94, 12), 456 => to_unsigned(3257, 12), 457 => to_unsigned(169, 12), 458 => to_unsigned(3924, 12), 459 => to_unsigned(3020, 12), 460 => to_unsigned(1610, 12), 461 => to_unsigned(7, 12), 462 => to_unsigned(2635, 12), 463 => to_unsigned(3653, 12), 464 => to_unsigned(518, 12), 465 => to_unsigned(2665, 12), 466 => to_unsigned(1066, 12), 467 => to_unsigned(3803, 12), 468 => to_unsigned(1900, 12), 469 => to_unsigned(3289, 12), 470 => to_unsigned(804, 12), 471 => to_unsigned(1016, 12), 472 => to_unsigned(3396, 12), 473 => to_unsigned(3371, 12), 474 => to_unsigned(1200, 12), 475 => to_unsigned(1668, 12), 476 => to_unsigned(2429, 12), 477 => to_unsigned(1003, 12), 478 => to_unsigned(2597, 12), 479 => to_unsigned(2885, 12), 480 => to_unsigned(1096, 12), 481 => to_unsigned(3406, 12), 482 => to_unsigned(1622, 12), 483 => to_unsigned(984, 12), 484 => to_unsigned(1721, 12), 485 => to_unsigned(3019, 12), 486 => to_unsigned(2955, 12), 487 => to_unsigned(804, 12), 488 => to_unsigned(1270, 12), 489 => to_unsigned(3327, 12), 490 => to_unsigned(3017, 12), 491 => to_unsigned(2863, 12), 492 => to_unsigned(2100, 12), 493 => to_unsigned(3879, 12), 494 => to_unsigned(1088, 12), 495 => to_unsigned(3141, 12), 496 => to_unsigned(1359, 12), 497 => to_unsigned(1397, 12), 498 => to_unsigned(2391, 12), 499 => to_unsigned(1298, 12), 500 => to_unsigned(3449, 12), 501 => to_unsigned(1141, 12), 502 => to_unsigned(2742, 12), 503 => to_unsigned(3849, 12), 504 => to_unsigned(1686, 12), 505 => to_unsigned(1065, 12), 506 => to_unsigned(3985, 12), 507 => to_unsigned(1936, 12), 508 => to_unsigned(890, 12), 509 => to_unsigned(2389, 12), 510 => to_unsigned(2859, 12), 511 => to_unsigned(2994, 12), 512 => to_unsigned(1719, 12), 513 => to_unsigned(1825, 12), 514 => to_unsigned(85, 12), 515 => to_unsigned(586, 12), 516 => to_unsigned(689, 12), 517 => to_unsigned(2127, 12), 518 => to_unsigned(368, 12), 519 => to_unsigned(2712, 12), 520 => to_unsigned(799, 12), 521 => to_unsigned(2084, 12), 522 => to_unsigned(1044, 12), 523 => to_unsigned(3252, 12), 524 => to_unsigned(575, 12), 525 => to_unsigned(637, 12), 526 => to_unsigned(1204, 12), 527 => to_unsigned(1978, 12), 528 => to_unsigned(2659, 12), 529 => to_unsigned(6, 12), 530 => to_unsigned(299, 12), 531 => to_unsigned(1363, 12), 532 => to_unsigned(1996, 12), 533 => to_unsigned(756, 12), 534 => to_unsigned(3359, 12), 535 => to_unsigned(2306, 12), 536 => to_unsigned(1816, 12), 537 => to_unsigned(555, 12), 538 => to_unsigned(1726, 12), 539 => to_unsigned(1601, 12), 540 => to_unsigned(1181, 12), 541 => to_unsigned(1822, 12), 542 => to_unsigned(1434, 12), 543 => to_unsigned(1413, 12), 544 => to_unsigned(2786, 12), 545 => to_unsigned(440, 12), 546 => to_unsigned(969, 12), 547 => to_unsigned(3464, 12), 548 => to_unsigned(376, 12), 549 => to_unsigned(3690, 12), 550 => to_unsigned(313, 12), 551 => to_unsigned(3789, 12), 552 => to_unsigned(382, 12), 553 => to_unsigned(3946, 12), 554 => to_unsigned(3935, 12), 555 => to_unsigned(2480, 12), 556 => to_unsigned(343, 12), 557 => to_unsigned(505, 12), 558 => to_unsigned(424, 12), 559 => to_unsigned(141, 12), 560 => to_unsigned(2114, 12), 561 => to_unsigned(4082, 12), 562 => to_unsigned(214, 12), 563 => to_unsigned(684, 12), 564 => to_unsigned(181, 12), 565 => to_unsigned(3833, 12), 566 => to_unsigned(657, 12), 567 => to_unsigned(2885, 12), 568 => to_unsigned(2621, 12), 569 => to_unsigned(1999, 12), 570 => to_unsigned(3769, 12), 571 => to_unsigned(174, 12), 572 => to_unsigned(1112, 12), 573 => to_unsigned(2579, 12), 574 => to_unsigned(900, 12), 575 => to_unsigned(3943, 12), 576 => to_unsigned(3072, 12), 577 => to_unsigned(2496, 12), 578 => to_unsigned(3815, 12), 579 => to_unsigned(2283, 12), 580 => to_unsigned(3018, 12), 581 => to_unsigned(3192, 12), 582 => to_unsigned(3677, 12), 583 => to_unsigned(1368, 12), 584 => to_unsigned(2185, 12), 585 => to_unsigned(139, 12), 586 => to_unsigned(3796, 12), 587 => to_unsigned(444, 12), 588 => to_unsigned(1601, 12), 589 => to_unsigned(3851, 12), 590 => to_unsigned(2565, 12), 591 => to_unsigned(986, 12), 592 => to_unsigned(2701, 12), 593 => to_unsigned(3587, 12), 594 => to_unsigned(1248, 12), 595 => to_unsigned(3680, 12), 596 => to_unsigned(2308, 12), 597 => to_unsigned(3564, 12), 598 => to_unsigned(2404, 12), 599 => to_unsigned(420, 12), 600 => to_unsigned(3521, 12), 601 => to_unsigned(2977, 12), 602 => to_unsigned(1017, 12), 603 => to_unsigned(3419, 12), 604 => to_unsigned(1848, 12), 605 => to_unsigned(2678, 12), 606 => to_unsigned(2923, 12), 607 => to_unsigned(2423, 12), 608 => to_unsigned(3115, 12), 609 => to_unsigned(3546, 12), 610 => to_unsigned(21, 12), 611 => to_unsigned(808, 12), 612 => to_unsigned(534, 12), 613 => to_unsigned(2403, 12), 614 => to_unsigned(206, 12), 615 => to_unsigned(3275, 12), 616 => to_unsigned(852, 12), 617 => to_unsigned(1207, 12), 618 => to_unsigned(15, 12), 619 => to_unsigned(194, 12), 620 => to_unsigned(82, 12), 621 => to_unsigned(1865, 12), 622 => to_unsigned(222, 12), 623 => to_unsigned(3287, 12), 624 => to_unsigned(310, 12), 625 => to_unsigned(1969, 12), 626 => to_unsigned(1464, 12), 627 => to_unsigned(2329, 12), 628 => to_unsigned(1415, 12), 629 => to_unsigned(3830, 12), 630 => to_unsigned(2186, 12), 631 => to_unsigned(3159, 12), 632 => to_unsigned(1958, 12), 633 => to_unsigned(3140, 12), 634 => to_unsigned(3124, 12), 635 => to_unsigned(784, 12), 636 => to_unsigned(1997, 12), 637 => to_unsigned(1009, 12), 638 => to_unsigned(2558, 12), 639 => to_unsigned(2848, 12), 640 => to_unsigned(2247, 12), 641 => to_unsigned(2414, 12), 642 => to_unsigned(865, 12), 643 => to_unsigned(3871, 12), 644 => to_unsigned(3426, 12), 645 => to_unsigned(924, 12), 646 => to_unsigned(2925, 12), 647 => to_unsigned(766, 12), 648 => to_unsigned(1722, 12), 649 => to_unsigned(429, 12), 650 => to_unsigned(3920, 12), 651 => to_unsigned(2951, 12), 652 => to_unsigned(1462, 12), 653 => to_unsigned(3546, 12), 654 => to_unsigned(1779, 12), 655 => to_unsigned(2073, 12), 656 => to_unsigned(1111, 12), 657 => to_unsigned(1542, 12), 658 => to_unsigned(542, 12), 659 => to_unsigned(3211, 12), 660 => to_unsigned(2161, 12), 661 => to_unsigned(23, 12), 662 => to_unsigned(2516, 12), 663 => to_unsigned(1095, 12), 664 => to_unsigned(320, 12), 665 => to_unsigned(3310, 12), 666 => to_unsigned(3707, 12), 667 => to_unsigned(1486, 12), 668 => to_unsigned(2378, 12), 669 => to_unsigned(1798, 12), 670 => to_unsigned(339, 12), 671 => to_unsigned(3651, 12), 672 => to_unsigned(2268, 12), 673 => to_unsigned(479, 12), 674 => to_unsigned(387, 12), 675 => to_unsigned(677, 12), 676 => to_unsigned(1125, 12), 677 => to_unsigned(3655, 12), 678 => to_unsigned(1224, 12), 679 => to_unsigned(241, 12), 680 => to_unsigned(2348, 12), 681 => to_unsigned(1904, 12), 682 => to_unsigned(260, 12), 683 => to_unsigned(3781, 12), 684 => to_unsigned(2955, 12), 685 => to_unsigned(659, 12), 686 => to_unsigned(1824, 12), 687 => to_unsigned(3062, 12), 688 => to_unsigned(464, 12), 689 => to_unsigned(1577, 12), 690 => to_unsigned(2800, 12), 691 => to_unsigned(1325, 12), 692 => to_unsigned(1734, 12), 693 => to_unsigned(2518, 12), 694 => to_unsigned(1378, 12), 695 => to_unsigned(1345, 12), 696 => to_unsigned(2810, 12), 697 => to_unsigned(3102, 12), 698 => to_unsigned(815, 12), 699 => to_unsigned(2684, 12), 700 => to_unsigned(1141, 12), 701 => to_unsigned(3425, 12), 702 => to_unsigned(2241, 12), 703 => to_unsigned(2465, 12), 704 => to_unsigned(3306, 12), 705 => to_unsigned(2113, 12), 706 => to_unsigned(509, 12), 707 => to_unsigned(1966, 12), 708 => to_unsigned(1554, 12), 709 => to_unsigned(1209, 12), 710 => to_unsigned(3789, 12), 711 => to_unsigned(2071, 12), 712 => to_unsigned(1087, 12), 713 => to_unsigned(528, 12), 714 => to_unsigned(2055, 12), 715 => to_unsigned(354, 12), 716 => to_unsigned(3050, 12), 717 => to_unsigned(3434, 12), 718 => to_unsigned(2850, 12), 719 => to_unsigned(1698, 12), 720 => to_unsigned(1796, 12), 721 => to_unsigned(3676, 12), 722 => to_unsigned(2749, 12), 723 => to_unsigned(3051, 12), 724 => to_unsigned(3624, 12), 725 => to_unsigned(2415, 12), 726 => to_unsigned(3152, 12), 727 => to_unsigned(1146, 12), 728 => to_unsigned(3092, 12), 729 => to_unsigned(1609, 12), 730 => to_unsigned(1851, 12), 731 => to_unsigned(549, 12), 732 => to_unsigned(1315, 12), 733 => to_unsigned(253, 12), 734 => to_unsigned(3934, 12), 735 => to_unsigned(2553, 12), 736 => to_unsigned(293, 12), 737 => to_unsigned(508, 12), 738 => to_unsigned(3762, 12), 739 => to_unsigned(1061, 12), 740 => to_unsigned(3985, 12), 741 => to_unsigned(623, 12), 742 => to_unsigned(690, 12), 743 => to_unsigned(1766, 12), 744 => to_unsigned(2224, 12), 745 => to_unsigned(3513, 12), 746 => to_unsigned(3637, 12), 747 => to_unsigned(1315, 12), 748 => to_unsigned(2609, 12), 749 => to_unsigned(270, 12), 750 => to_unsigned(3112, 12), 751 => to_unsigned(133, 12), 752 => to_unsigned(4006, 12), 753 => to_unsigned(3164, 12), 754 => to_unsigned(90, 12), 755 => to_unsigned(2113, 12), 756 => to_unsigned(955, 12), 757 => to_unsigned(742, 12), 758 => to_unsigned(2677, 12), 759 => to_unsigned(345, 12), 760 => to_unsigned(2772, 12), 761 => to_unsigned(2826, 12), 762 => to_unsigned(1605, 12), 763 => to_unsigned(1086, 12), 764 => to_unsigned(1126, 12), 765 => to_unsigned(3896, 12), 766 => to_unsigned(1089, 12), 767 => to_unsigned(1136, 12), 768 => to_unsigned(1211, 12), 769 => to_unsigned(1642, 12), 770 => to_unsigned(1837, 12), 771 => to_unsigned(260, 12), 772 => to_unsigned(3490, 12), 773 => to_unsigned(1059, 12), 774 => to_unsigned(2608, 12), 775 => to_unsigned(2639, 12), 776 => to_unsigned(1705, 12), 777 => to_unsigned(1512, 12), 778 => to_unsigned(1968, 12), 779 => to_unsigned(2243, 12), 780 => to_unsigned(1395, 12), 781 => to_unsigned(1996, 12), 782 => to_unsigned(2374, 12), 783 => to_unsigned(3964, 12), 784 => to_unsigned(3155, 12), 785 => to_unsigned(4086, 12), 786 => to_unsigned(1346, 12), 787 => to_unsigned(3456, 12), 788 => to_unsigned(3657, 12), 789 => to_unsigned(1105, 12), 790 => to_unsigned(3605, 12), 791 => to_unsigned(1351, 12), 792 => to_unsigned(3761, 12), 793 => to_unsigned(3467, 12), 794 => to_unsigned(84, 12), 795 => to_unsigned(4088, 12), 796 => to_unsigned(1010, 12), 797 => to_unsigned(2443, 12), 798 => to_unsigned(1487, 12), 799 => to_unsigned(3262, 12), 800 => to_unsigned(4055, 12), 801 => to_unsigned(831, 12), 802 => to_unsigned(3919, 12), 803 => to_unsigned(3446, 12), 804 => to_unsigned(1555, 12), 805 => to_unsigned(2662, 12), 806 => to_unsigned(1043, 12), 807 => to_unsigned(2593, 12), 808 => to_unsigned(1135, 12), 809 => to_unsigned(639, 12), 810 => to_unsigned(1684, 12), 811 => to_unsigned(2005, 12), 812 => to_unsigned(2511, 12), 813 => to_unsigned(1133, 12), 814 => to_unsigned(1962, 12), 815 => to_unsigned(135, 12), 816 => to_unsigned(1826, 12), 817 => to_unsigned(653, 12), 818 => to_unsigned(111, 12), 819 => to_unsigned(3183, 12), 820 => to_unsigned(3223, 12), 821 => to_unsigned(1510, 12), 822 => to_unsigned(603, 12), 823 => to_unsigned(1827, 12), 824 => to_unsigned(945, 12), 825 => to_unsigned(1606, 12), 826 => to_unsigned(382, 12), 827 => to_unsigned(114, 12), 828 => to_unsigned(2264, 12), 829 => to_unsigned(3919, 12), 830 => to_unsigned(4036, 12), 831 => to_unsigned(2950, 12), 832 => to_unsigned(2887, 12), 833 => to_unsigned(2497, 12), 834 => to_unsigned(3797, 12), 835 => to_unsigned(3652, 12), 836 => to_unsigned(3940, 12), 837 => to_unsigned(1740, 12), 838 => to_unsigned(1323, 12), 839 => to_unsigned(559, 12), 840 => to_unsigned(1332, 12), 841 => to_unsigned(670, 12), 842 => to_unsigned(1099, 12), 843 => to_unsigned(2198, 12), 844 => to_unsigned(2947, 12), 845 => to_unsigned(4087, 12), 846 => to_unsigned(3037, 12), 847 => to_unsigned(2540, 12), 848 => to_unsigned(3203, 12), 849 => to_unsigned(1969, 12), 850 => to_unsigned(2710, 12), 851 => to_unsigned(3138, 12), 852 => to_unsigned(1573, 12), 853 => to_unsigned(2706, 12), 854 => to_unsigned(1915, 12), 855 => to_unsigned(2232, 12), 856 => to_unsigned(3029, 12), 857 => to_unsigned(3771, 12), 858 => to_unsigned(1859, 12), 859 => to_unsigned(39, 12), 860 => to_unsigned(388, 12), 861 => to_unsigned(844, 12), 862 => to_unsigned(1332, 12), 863 => to_unsigned(817, 12), 864 => to_unsigned(864, 12), 865 => to_unsigned(2642, 12), 866 => to_unsigned(2424, 12), 867 => to_unsigned(1211, 12), 868 => to_unsigned(3747, 12), 869 => to_unsigned(1606, 12), 870 => to_unsigned(860, 12), 871 => to_unsigned(1623, 12), 872 => to_unsigned(2456, 12), 873 => to_unsigned(2651, 12), 874 => to_unsigned(146, 12), 875 => to_unsigned(3728, 12), 876 => to_unsigned(2425, 12), 877 => to_unsigned(2468, 12), 878 => to_unsigned(3632, 12), 879 => to_unsigned(1769, 12), 880 => to_unsigned(1456, 12), 881 => to_unsigned(959, 12), 882 => to_unsigned(2433, 12), 883 => to_unsigned(3764, 12), 884 => to_unsigned(1294, 12), 885 => to_unsigned(2075, 12), 886 => to_unsigned(13, 12), 887 => to_unsigned(1142, 12), 888 => to_unsigned(2738, 12), 889 => to_unsigned(3917, 12), 890 => to_unsigned(1260, 12), 891 => to_unsigned(2842, 12), 892 => to_unsigned(3988, 12), 893 => to_unsigned(3834, 12), 894 => to_unsigned(3982, 12), 895 => to_unsigned(2771, 12), 896 => to_unsigned(4071, 12), 897 => to_unsigned(1242, 12), 898 => to_unsigned(1681, 12), 899 => to_unsigned(85, 12), 900 => to_unsigned(928, 12), 901 => to_unsigned(2392, 12), 902 => to_unsigned(102, 12), 903 => to_unsigned(711, 12), 904 => to_unsigned(3803, 12), 905 => to_unsigned(2632, 12), 906 => to_unsigned(3630, 12), 907 => to_unsigned(3158, 12), 908 => to_unsigned(269, 12), 909 => to_unsigned(621, 12), 910 => to_unsigned(687, 12), 911 => to_unsigned(2334, 12), 912 => to_unsigned(2946, 12), 913 => to_unsigned(1519, 12), 914 => to_unsigned(3609, 12), 915 => to_unsigned(1896, 12), 916 => to_unsigned(3067, 12), 917 => to_unsigned(3559, 12), 918 => to_unsigned(237, 12), 919 => to_unsigned(2932, 12), 920 => to_unsigned(2683, 12), 921 => to_unsigned(3149, 12), 922 => to_unsigned(2526, 12), 923 => to_unsigned(1575, 12), 924 => to_unsigned(3678, 12), 925 => to_unsigned(2733, 12), 926 => to_unsigned(2880, 12), 927 => to_unsigned(291, 12), 928 => to_unsigned(1070, 12), 929 => to_unsigned(2691, 12), 930 => to_unsigned(3757, 12), 931 => to_unsigned(1869, 12), 932 => to_unsigned(3964, 12), 933 => to_unsigned(2313, 12), 934 => to_unsigned(2071, 12), 935 => to_unsigned(1736, 12), 936 => to_unsigned(3117, 12), 937 => to_unsigned(623, 12), 938 => to_unsigned(2490, 12), 939 => to_unsigned(528, 12), 940 => to_unsigned(3516, 12), 941 => to_unsigned(2597, 12), 942 => to_unsigned(3942, 12), 943 => to_unsigned(2093, 12), 944 => to_unsigned(3445, 12), 945 => to_unsigned(3321, 12), 946 => to_unsigned(2978, 12), 947 => to_unsigned(1772, 12), 948 => to_unsigned(3847, 12), 949 => to_unsigned(378, 12), 950 => to_unsigned(479, 12), 951 => to_unsigned(1350, 12), 952 => to_unsigned(1899, 12), 953 => to_unsigned(585, 12), 954 => to_unsigned(3355, 12), 955 => to_unsigned(4042, 12), 956 => to_unsigned(263, 12), 957 => to_unsigned(3051, 12), 958 => to_unsigned(1880, 12), 959 => to_unsigned(1423, 12), 960 => to_unsigned(2812, 12), 961 => to_unsigned(543, 12), 962 => to_unsigned(483, 12), 963 => to_unsigned(227, 12), 964 => to_unsigned(1726, 12), 965 => to_unsigned(742, 12), 966 => to_unsigned(1369, 12), 967 => to_unsigned(1609, 12), 968 => to_unsigned(2222, 12), 969 => to_unsigned(679, 12), 970 => to_unsigned(3323, 12), 971 => to_unsigned(3391, 12), 972 => to_unsigned(1054, 12), 973 => to_unsigned(1053, 12), 974 => to_unsigned(3987, 12), 975 => to_unsigned(161, 12), 976 => to_unsigned(1614, 12), 977 => to_unsigned(1991, 12), 978 => to_unsigned(3685, 12), 979 => to_unsigned(3344, 12), 980 => to_unsigned(3305, 12), 981 => to_unsigned(2174, 12), 982 => to_unsigned(2934, 12), 983 => to_unsigned(508, 12), 984 => to_unsigned(2123, 12), 985 => to_unsigned(730, 12), 986 => to_unsigned(28, 12), 987 => to_unsigned(134, 12), 988 => to_unsigned(1431, 12), 989 => to_unsigned(1233, 12), 990 => to_unsigned(1756, 12), 991 => to_unsigned(4031, 12), 992 => to_unsigned(1902, 12), 993 => to_unsigned(168, 12), 994 => to_unsigned(3363, 12), 995 => to_unsigned(3164, 12), 996 => to_unsigned(2611, 12), 997 => to_unsigned(3473, 12), 998 => to_unsigned(690, 12), 999 => to_unsigned(1714, 12), 1000 => to_unsigned(3997, 12), 1001 => to_unsigned(2892, 12), 1002 => to_unsigned(1021, 12), 1003 => to_unsigned(597, 12), 1004 => to_unsigned(2286, 12), 1005 => to_unsigned(2565, 12), 1006 => to_unsigned(810, 12), 1007 => to_unsigned(644, 12), 1008 => to_unsigned(3242, 12), 1009 => to_unsigned(2809, 12), 1010 => to_unsigned(1304, 12), 1011 => to_unsigned(3335, 12), 1012 => to_unsigned(3737, 12), 1013 => to_unsigned(935, 12), 1014 => to_unsigned(2126, 12), 1015 => to_unsigned(3628, 12), 1016 => to_unsigned(2193, 12), 1017 => to_unsigned(2883, 12), 1018 => to_unsigned(669, 12), 1019 => to_unsigned(1078, 12), 1020 => to_unsigned(301, 12), 1021 => to_unsigned(3811, 12), 1022 => to_unsigned(1889, 12), 1023 => to_unsigned(572, 12), 1024 => to_unsigned(2815, 12), 1025 => to_unsigned(852, 12), 1026 => to_unsigned(3222, 12), 1027 => to_unsigned(1714, 12), 1028 => to_unsigned(2350, 12), 1029 => to_unsigned(2522, 12), 1030 => to_unsigned(3000, 12), 1031 => to_unsigned(3714, 12), 1032 => to_unsigned(2027, 12), 1033 => to_unsigned(1131, 12), 1034 => to_unsigned(428, 12), 1035 => to_unsigned(2350, 12), 1036 => to_unsigned(3090, 12), 1037 => to_unsigned(1026, 12), 1038 => to_unsigned(4080, 12), 1039 => to_unsigned(1793, 12), 1040 => to_unsigned(3130, 12), 1041 => to_unsigned(3922, 12), 1042 => to_unsigned(3264, 12), 1043 => to_unsigned(881, 12), 1044 => to_unsigned(3343, 12), 1045 => to_unsigned(1806, 12), 1046 => to_unsigned(1873, 12), 1047 => to_unsigned(2282, 12), 1048 => to_unsigned(818, 12), 1049 => to_unsigned(1980, 12), 1050 => to_unsigned(2349, 12), 1051 => to_unsigned(2314, 12), 1052 => to_unsigned(1488, 12), 1053 => to_unsigned(236, 12), 1054 => to_unsigned(2794, 12), 1055 => to_unsigned(1988, 12), 1056 => to_unsigned(3944, 12), 1057 => to_unsigned(3850, 12), 1058 => to_unsigned(4068, 12), 1059 => to_unsigned(3766, 12), 1060 => to_unsigned(2678, 12), 1061 => to_unsigned(4023, 12), 1062 => to_unsigned(2484, 12), 1063 => to_unsigned(3034, 12), 1064 => to_unsigned(1774, 12), 1065 => to_unsigned(1739, 12), 1066 => to_unsigned(2352, 12), 1067 => to_unsigned(4022, 12), 1068 => to_unsigned(288, 12), 1069 => to_unsigned(3147, 12), 1070 => to_unsigned(556, 12), 1071 => to_unsigned(2943, 12), 1072 => to_unsigned(3969, 12), 1073 => to_unsigned(200, 12), 1074 => to_unsigned(3398, 12), 1075 => to_unsigned(2494, 12), 1076 => to_unsigned(291, 12), 1077 => to_unsigned(3661, 12), 1078 => to_unsigned(1692, 12), 1079 => to_unsigned(3946, 12), 1080 => to_unsigned(1241, 12), 1081 => to_unsigned(3775, 12), 1082 => to_unsigned(539, 12), 1083 => to_unsigned(3794, 12), 1084 => to_unsigned(894, 12), 1085 => to_unsigned(2070, 12), 1086 => to_unsigned(3946, 12), 1087 => to_unsigned(138, 12), 1088 => to_unsigned(2617, 12), 1089 => to_unsigned(3223, 12), 1090 => to_unsigned(107, 12), 1091 => to_unsigned(825, 12), 1092 => to_unsigned(3358, 12), 1093 => to_unsigned(1070, 12), 1094 => to_unsigned(1667, 12), 1095 => to_unsigned(1286, 12), 1096 => to_unsigned(899, 12), 1097 => to_unsigned(740, 12), 1098 => to_unsigned(3280, 12), 1099 => to_unsigned(3152, 12), 1100 => to_unsigned(1059, 12), 1101 => to_unsigned(2937, 12), 1102 => to_unsigned(3324, 12), 1103 => to_unsigned(1234, 12), 1104 => to_unsigned(2346, 12), 1105 => to_unsigned(3175, 12), 1106 => to_unsigned(3327, 12), 1107 => to_unsigned(1385, 12), 1108 => to_unsigned(3183, 12), 1109 => to_unsigned(3562, 12), 1110 => to_unsigned(1626, 12), 1111 => to_unsigned(3798, 12), 1112 => to_unsigned(2015, 12), 1113 => to_unsigned(3710, 12), 1114 => to_unsigned(1124, 12), 1115 => to_unsigned(1196, 12), 1116 => to_unsigned(1934, 12), 1117 => to_unsigned(2917, 12), 1118 => to_unsigned(3341, 12), 1119 => to_unsigned(3262, 12), 1120 => to_unsigned(2203, 12), 1121 => to_unsigned(1947, 12), 1122 => to_unsigned(2032, 12), 1123 => to_unsigned(1527, 12), 1124 => to_unsigned(1903, 12), 1125 => to_unsigned(1749, 12), 1126 => to_unsigned(2047, 12), 1127 => to_unsigned(2481, 12), 1128 => to_unsigned(1053, 12), 1129 => to_unsigned(1773, 12), 1130 => to_unsigned(946, 12), 1131 => to_unsigned(2506, 12), 1132 => to_unsigned(2737, 12), 1133 => to_unsigned(3370, 12), 1134 => to_unsigned(3377, 12), 1135 => to_unsigned(2922, 12), 1136 => to_unsigned(2273, 12), 1137 => to_unsigned(3300, 12), 1138 => to_unsigned(1121, 12), 1139 => to_unsigned(1431, 12), 1140 => to_unsigned(1975, 12), 1141 => to_unsigned(2762, 12), 1142 => to_unsigned(1783, 12), 1143 => to_unsigned(2390, 12), 1144 => to_unsigned(157, 12), 1145 => to_unsigned(3714, 12), 1146 => to_unsigned(2300, 12), 1147 => to_unsigned(3043, 12), 1148 => to_unsigned(3070, 12), 1149 => to_unsigned(1816, 12), 1150 => to_unsigned(2697, 12), 1151 => to_unsigned(738, 12), 1152 => to_unsigned(672, 12), 1153 => to_unsigned(3305, 12), 1154 => to_unsigned(3761, 12), 1155 => to_unsigned(3287, 12), 1156 => to_unsigned(3326, 12), 1157 => to_unsigned(1951, 12), 1158 => to_unsigned(1344, 12), 1159 => to_unsigned(3770, 12), 1160 => to_unsigned(1477, 12), 1161 => to_unsigned(145, 12), 1162 => to_unsigned(1852, 12), 1163 => to_unsigned(767, 12), 1164 => to_unsigned(1535, 12), 1165 => to_unsigned(1379, 12), 1166 => to_unsigned(2926, 12), 1167 => to_unsigned(1396, 12), 1168 => to_unsigned(1716, 12), 1169 => to_unsigned(1922, 12), 1170 => to_unsigned(1052, 12), 1171 => to_unsigned(2303, 12), 1172 => to_unsigned(3250, 12), 1173 => to_unsigned(2603, 12), 1174 => to_unsigned(1934, 12), 1175 => to_unsigned(3152, 12), 1176 => to_unsigned(1500, 12), 1177 => to_unsigned(1352, 12), 1178 => to_unsigned(1839, 12), 1179 => to_unsigned(3263, 12), 1180 => to_unsigned(3833, 12), 1181 => to_unsigned(3271, 12), 1182 => to_unsigned(241, 12), 1183 => to_unsigned(1394, 12), 1184 => to_unsigned(476, 12), 1185 => to_unsigned(279, 12), 1186 => to_unsigned(776, 12), 1187 => to_unsigned(1996, 12), 1188 => to_unsigned(1333, 12), 1189 => to_unsigned(3348, 12), 1190 => to_unsigned(1658, 12), 1191 => to_unsigned(2677, 12), 1192 => to_unsigned(3801, 12), 1193 => to_unsigned(2718, 12), 1194 => to_unsigned(95, 12), 1195 => to_unsigned(3733, 12), 1196 => to_unsigned(2206, 12), 1197 => to_unsigned(1987, 12), 1198 => to_unsigned(1430, 12), 1199 => to_unsigned(3725, 12), 1200 => to_unsigned(4080, 12), 1201 => to_unsigned(1643, 12), 1202 => to_unsigned(2807, 12), 1203 => to_unsigned(3522, 12), 1204 => to_unsigned(1820, 12), 1205 => to_unsigned(2228, 12), 1206 => to_unsigned(2141, 12), 1207 => to_unsigned(34, 12), 1208 => to_unsigned(3737, 12), 1209 => to_unsigned(2389, 12), 1210 => to_unsigned(1717, 12), 1211 => to_unsigned(71, 12), 1212 => to_unsigned(3586, 12), 1213 => to_unsigned(3183, 12), 1214 => to_unsigned(848, 12), 1215 => to_unsigned(2320, 12), 1216 => to_unsigned(493, 12), 1217 => to_unsigned(3614, 12), 1218 => to_unsigned(3107, 12), 1219 => to_unsigned(2177, 12), 1220 => to_unsigned(1705, 12), 1221 => to_unsigned(90, 12), 1222 => to_unsigned(2736, 12), 1223 => to_unsigned(3001, 12), 1224 => to_unsigned(2424, 12), 1225 => to_unsigned(42, 12), 1226 => to_unsigned(1322, 12), 1227 => to_unsigned(1422, 12), 1228 => to_unsigned(1144, 12), 1229 => to_unsigned(2240, 12), 1230 => to_unsigned(2989, 12), 1231 => to_unsigned(487, 12), 1232 => to_unsigned(1324, 12), 1233 => to_unsigned(2741, 12), 1234 => to_unsigned(283, 12), 1235 => to_unsigned(1549, 12), 1236 => to_unsigned(3233, 12), 1237 => to_unsigned(2111, 12), 1238 => to_unsigned(3287, 12), 1239 => to_unsigned(3167, 12), 1240 => to_unsigned(2085, 12), 1241 => to_unsigned(274, 12), 1242 => to_unsigned(1999, 12), 1243 => to_unsigned(3930, 12), 1244 => to_unsigned(889, 12), 1245 => to_unsigned(1603, 12), 1246 => to_unsigned(1031, 12), 1247 => to_unsigned(1205, 12), 1248 => to_unsigned(3579, 12), 1249 => to_unsigned(139, 12), 1250 => to_unsigned(3553, 12), 1251 => to_unsigned(136, 12), 1252 => to_unsigned(452, 12), 1253 => to_unsigned(44, 12), 1254 => to_unsigned(3608, 12), 1255 => to_unsigned(1994, 12), 1256 => to_unsigned(2588, 12), 1257 => to_unsigned(3124, 12), 1258 => to_unsigned(2784, 12), 1259 => to_unsigned(3598, 12), 1260 => to_unsigned(1835, 12), 1261 => to_unsigned(1736, 12), 1262 => to_unsigned(3849, 12), 1263 => to_unsigned(434, 12), 1264 => to_unsigned(1390, 12), 1265 => to_unsigned(2019, 12), 1266 => to_unsigned(3586, 12), 1267 => to_unsigned(3007, 12), 1268 => to_unsigned(3178, 12), 1269 => to_unsigned(3933, 12), 1270 => to_unsigned(2280, 12), 1271 => to_unsigned(2205, 12), 1272 => to_unsigned(632, 12), 1273 => to_unsigned(585, 12), 1274 => to_unsigned(3936, 12), 1275 => to_unsigned(4037, 12), 1276 => to_unsigned(868, 12), 1277 => to_unsigned(921, 12), 1278 => to_unsigned(2090, 12), 1279 => to_unsigned(3554, 12), 1280 => to_unsigned(1409, 12), 1281 => to_unsigned(3323, 12), 1282 => to_unsigned(827, 12), 1283 => to_unsigned(2153, 12), 1284 => to_unsigned(1358, 12), 1285 => to_unsigned(1152, 12), 1286 => to_unsigned(2831, 12), 1287 => to_unsigned(1993, 12), 1288 => to_unsigned(2167, 12), 1289 => to_unsigned(1760, 12), 1290 => to_unsigned(2445, 12), 1291 => to_unsigned(1872, 12), 1292 => to_unsigned(1603, 12), 1293 => to_unsigned(1126, 12), 1294 => to_unsigned(3509, 12), 1295 => to_unsigned(2827, 12), 1296 => to_unsigned(749, 12), 1297 => to_unsigned(3408, 12), 1298 => to_unsigned(3513, 12), 1299 => to_unsigned(1486, 12), 1300 => to_unsigned(3697, 12), 1301 => to_unsigned(100, 12), 1302 => to_unsigned(2238, 12), 1303 => to_unsigned(3045, 12), 1304 => to_unsigned(2075, 12), 1305 => to_unsigned(3777, 12), 1306 => to_unsigned(1218, 12), 1307 => to_unsigned(2497, 12), 1308 => to_unsigned(1665, 12), 1309 => to_unsigned(1956, 12), 1310 => to_unsigned(228, 12), 1311 => to_unsigned(418, 12), 1312 => to_unsigned(2501, 12), 1313 => to_unsigned(613, 12), 1314 => to_unsigned(3811, 12), 1315 => to_unsigned(1230, 12), 1316 => to_unsigned(3064, 12), 1317 => to_unsigned(2314, 12), 1318 => to_unsigned(2164, 12), 1319 => to_unsigned(2632, 12), 1320 => to_unsigned(2579, 12), 1321 => to_unsigned(3606, 12), 1322 => to_unsigned(2378, 12), 1323 => to_unsigned(592, 12), 1324 => to_unsigned(3037, 12), 1325 => to_unsigned(2491, 12), 1326 => to_unsigned(2870, 12), 1327 => to_unsigned(1656, 12), 1328 => to_unsigned(3759, 12), 1329 => to_unsigned(1991, 12), 1330 => to_unsigned(2717, 12), 1331 => to_unsigned(1736, 12), 1332 => to_unsigned(2650, 12), 1333 => to_unsigned(734, 12), 1334 => to_unsigned(4032, 12), 1335 => to_unsigned(716, 12), 1336 => to_unsigned(3525, 12), 1337 => to_unsigned(3830, 12), 1338 => to_unsigned(240, 12), 1339 => to_unsigned(1622, 12), 1340 => to_unsigned(2538, 12), 1341 => to_unsigned(425, 12), 1342 => to_unsigned(1378, 12), 1343 => to_unsigned(1895, 12), 1344 => to_unsigned(473, 12), 1345 => to_unsigned(1338, 12), 1346 => to_unsigned(1484, 12), 1347 => to_unsigned(2667, 12), 1348 => to_unsigned(1106, 12), 1349 => to_unsigned(299, 12), 1350 => to_unsigned(300, 12), 1351 => to_unsigned(467, 12), 1352 => to_unsigned(373, 12), 1353 => to_unsigned(1498, 12), 1354 => to_unsigned(3670, 12), 1355 => to_unsigned(715, 12), 1356 => to_unsigned(3133, 12), 1357 => to_unsigned(2813, 12), 1358 => to_unsigned(632, 12), 1359 => to_unsigned(856, 12), 1360 => to_unsigned(3975, 12), 1361 => to_unsigned(1558, 12), 1362 => to_unsigned(298, 12), 1363 => to_unsigned(2380, 12), 1364 => to_unsigned(2805, 12), 1365 => to_unsigned(1188, 12), 1366 => to_unsigned(2145, 12), 1367 => to_unsigned(362, 12), 1368 => to_unsigned(2987, 12), 1369 => to_unsigned(3900, 12), 1370 => to_unsigned(1602, 12), 1371 => to_unsigned(456, 12), 1372 => to_unsigned(738, 12), 1373 => to_unsigned(2172, 12), 1374 => to_unsigned(893, 12), 1375 => to_unsigned(2495, 12), 1376 => to_unsigned(223, 12), 1377 => to_unsigned(44, 12), 1378 => to_unsigned(2273, 12), 1379 => to_unsigned(3083, 12), 1380 => to_unsigned(1338, 12), 1381 => to_unsigned(1220, 12), 1382 => to_unsigned(2873, 12), 1383 => to_unsigned(2965, 12), 1384 => to_unsigned(4021, 12), 1385 => to_unsigned(262, 12), 1386 => to_unsigned(2663, 12), 1387 => to_unsigned(3097, 12), 1388 => to_unsigned(803, 12), 1389 => to_unsigned(276, 12), 1390 => to_unsigned(3635, 12), 1391 => to_unsigned(3703, 12), 1392 => to_unsigned(522, 12), 1393 => to_unsigned(1493, 12), 1394 => to_unsigned(541, 12), 1395 => to_unsigned(800, 12), 1396 => to_unsigned(3577, 12), 1397 => to_unsigned(2530, 12), 1398 => to_unsigned(388, 12), 1399 => to_unsigned(3314, 12), 1400 => to_unsigned(2644, 12), 1401 => to_unsigned(1310, 12), 1402 => to_unsigned(942, 12), 1403 => to_unsigned(2062, 12), 1404 => to_unsigned(2428, 12), 1405 => to_unsigned(4059, 12), 1406 => to_unsigned(822, 12), 1407 => to_unsigned(2533, 12), 1408 => to_unsigned(307, 12), 1409 => to_unsigned(3533, 12), 1410 => to_unsigned(3666, 12), 1411 => to_unsigned(350, 12), 1412 => to_unsigned(124, 12), 1413 => to_unsigned(2081, 12), 1414 => to_unsigned(125, 12), 1415 => to_unsigned(719, 12), 1416 => to_unsigned(3045, 12), 1417 => to_unsigned(3498, 12), 1418 => to_unsigned(3125, 12), 1419 => to_unsigned(2480, 12), 1420 => to_unsigned(3844, 12), 1421 => to_unsigned(958, 12), 1422 => to_unsigned(2966, 12), 1423 => to_unsigned(4045, 12), 1424 => to_unsigned(1479, 12), 1425 => to_unsigned(330, 12), 1426 => to_unsigned(3563, 12), 1427 => to_unsigned(304, 12), 1428 => to_unsigned(320, 12), 1429 => to_unsigned(1987, 12), 1430 => to_unsigned(2903, 12), 1431 => to_unsigned(2316, 12), 1432 => to_unsigned(3377, 12), 1433 => to_unsigned(3744, 12), 1434 => to_unsigned(338, 12), 1435 => to_unsigned(2807, 12), 1436 => to_unsigned(2872, 12), 1437 => to_unsigned(1741, 12), 1438 => to_unsigned(1745, 12), 1439 => to_unsigned(2073, 12), 1440 => to_unsigned(3359, 12), 1441 => to_unsigned(798, 12), 1442 => to_unsigned(280, 12), 1443 => to_unsigned(630, 12), 1444 => to_unsigned(367, 12), 1445 => to_unsigned(1533, 12), 1446 => to_unsigned(1584, 12), 1447 => to_unsigned(2952, 12), 1448 => to_unsigned(1748, 12), 1449 => to_unsigned(2351, 12), 1450 => to_unsigned(1910, 12), 1451 => to_unsigned(1, 12), 1452 => to_unsigned(3531, 12), 1453 => to_unsigned(250, 12), 1454 => to_unsigned(2913, 12), 1455 => to_unsigned(138, 12), 1456 => to_unsigned(378, 12), 1457 => to_unsigned(1827, 12), 1458 => to_unsigned(3627, 12), 1459 => to_unsigned(1898, 12), 1460 => to_unsigned(3463, 12), 1461 => to_unsigned(894, 12), 1462 => to_unsigned(2373, 12), 1463 => to_unsigned(2318, 12), 1464 => to_unsigned(1688, 12), 1465 => to_unsigned(2836, 12), 1466 => to_unsigned(3626, 12), 1467 => to_unsigned(901, 12), 1468 => to_unsigned(175, 12), 1469 => to_unsigned(2621, 12), 1470 => to_unsigned(2467, 12), 1471 => to_unsigned(2511, 12), 1472 => to_unsigned(3264, 12), 1473 => to_unsigned(2063, 12), 1474 => to_unsigned(2246, 12), 1475 => to_unsigned(1630, 12), 1476 => to_unsigned(630, 12), 1477 => to_unsigned(1142, 12), 1478 => to_unsigned(1037, 12), 1479 => to_unsigned(3555, 12), 1480 => to_unsigned(3080, 12), 1481 => to_unsigned(2612, 12), 1482 => to_unsigned(1503, 12), 1483 => to_unsigned(3300, 12), 1484 => to_unsigned(4005, 12), 1485 => to_unsigned(2076, 12), 1486 => to_unsigned(2765, 12), 1487 => to_unsigned(3825, 12), 1488 => to_unsigned(1009, 12), 1489 => to_unsigned(2509, 12), 1490 => to_unsigned(2397, 12), 1491 => to_unsigned(655, 12), 1492 => to_unsigned(622, 12), 1493 => to_unsigned(491, 12), 1494 => to_unsigned(412, 12), 1495 => to_unsigned(1169, 12), 1496 => to_unsigned(1700, 12), 1497 => to_unsigned(3088, 12), 1498 => to_unsigned(2427, 12), 1499 => to_unsigned(1781, 12), 1500 => to_unsigned(3506, 12), 1501 => to_unsigned(2948, 12), 1502 => to_unsigned(1131, 12), 1503 => to_unsigned(3276, 12), 1504 => to_unsigned(3791, 12), 1505 => to_unsigned(650, 12), 1506 => to_unsigned(1567, 12), 1507 => to_unsigned(4078, 12), 1508 => to_unsigned(2059, 12), 1509 => to_unsigned(860, 12), 1510 => to_unsigned(154, 12), 1511 => to_unsigned(851, 12), 1512 => to_unsigned(3, 12), 1513 => to_unsigned(101, 12), 1514 => to_unsigned(1603, 12), 1515 => to_unsigned(1896, 12), 1516 => to_unsigned(2894, 12), 1517 => to_unsigned(2261, 12), 1518 => to_unsigned(526, 12), 1519 => to_unsigned(3496, 12), 1520 => to_unsigned(2072, 12), 1521 => to_unsigned(3460, 12), 1522 => to_unsigned(3273, 12), 1523 => to_unsigned(1275, 12), 1524 => to_unsigned(404, 12), 1525 => to_unsigned(3095, 12), 1526 => to_unsigned(1138, 12), 1527 => to_unsigned(1017, 12), 1528 => to_unsigned(2416, 12), 1529 => to_unsigned(2733, 12), 1530 => to_unsigned(1266, 12), 1531 => to_unsigned(519, 12), 1532 => to_unsigned(1304, 12), 1533 => to_unsigned(1245, 12), 1534 => to_unsigned(2306, 12), 1535 => to_unsigned(3444, 12), 1536 => to_unsigned(3058, 12), 1537 => to_unsigned(3369, 12), 1538 => to_unsigned(3783, 12), 1539 => to_unsigned(50, 12), 1540 => to_unsigned(3847, 12), 1541 => to_unsigned(4, 12), 1542 => to_unsigned(2079, 12), 1543 => to_unsigned(1271, 12), 1544 => to_unsigned(687, 12), 1545 => to_unsigned(2715, 12), 1546 => to_unsigned(1035, 12), 1547 => to_unsigned(1095, 12), 1548 => to_unsigned(1025, 12), 1549 => to_unsigned(2221, 12), 1550 => to_unsigned(2871, 12), 1551 => to_unsigned(1878, 12), 1552 => to_unsigned(2581, 12), 1553 => to_unsigned(2590, 12), 1554 => to_unsigned(1141, 12), 1555 => to_unsigned(616, 12), 1556 => to_unsigned(27, 12), 1557 => to_unsigned(3228, 12), 1558 => to_unsigned(4028, 12), 1559 => to_unsigned(1071, 12), 1560 => to_unsigned(596, 12), 1561 => to_unsigned(3521, 12), 1562 => to_unsigned(2996, 12), 1563 => to_unsigned(2527, 12), 1564 => to_unsigned(2125, 12), 1565 => to_unsigned(1005, 12), 1566 => to_unsigned(2373, 12), 1567 => to_unsigned(1457, 12), 1568 => to_unsigned(1834, 12), 1569 => to_unsigned(3896, 12), 1570 => to_unsigned(1290, 12), 1571 => to_unsigned(2826, 12), 1572 => to_unsigned(3249, 12), 1573 => to_unsigned(1464, 12), 1574 => to_unsigned(3114, 12), 1575 => to_unsigned(2941, 12), 1576 => to_unsigned(424, 12), 1577 => to_unsigned(3790, 12), 1578 => to_unsigned(3808, 12), 1579 => to_unsigned(2355, 12), 1580 => to_unsigned(3057, 12), 1581 => to_unsigned(2820, 12), 1582 => to_unsigned(3636, 12), 1583 => to_unsigned(858, 12), 1584 => to_unsigned(3240, 12), 1585 => to_unsigned(1302, 12), 1586 => to_unsigned(1926, 12), 1587 => to_unsigned(2992, 12), 1588 => to_unsigned(703, 12), 1589 => to_unsigned(2502, 12), 1590 => to_unsigned(1520, 12), 1591 => to_unsigned(1272, 12), 1592 => to_unsigned(262, 12), 1593 => to_unsigned(2925, 12), 1594 => to_unsigned(3453, 12), 1595 => to_unsigned(2087, 12), 1596 => to_unsigned(1076, 12), 1597 => to_unsigned(496, 12), 1598 => to_unsigned(1219, 12), 1599 => to_unsigned(1526, 12), 1600 => to_unsigned(1239, 12), 1601 => to_unsigned(1010, 12), 1602 => to_unsigned(2370, 12), 1603 => to_unsigned(3895, 12), 1604 => to_unsigned(773, 12), 1605 => to_unsigned(3795, 12), 1606 => to_unsigned(3333, 12), 1607 => to_unsigned(2547, 12), 1608 => to_unsigned(3915, 12), 1609 => to_unsigned(3740, 12), 1610 => to_unsigned(86, 12), 1611 => to_unsigned(2966, 12), 1612 => to_unsigned(1785, 12), 1613 => to_unsigned(3486, 12), 1614 => to_unsigned(2280, 12), 1615 => to_unsigned(421, 12), 1616 => to_unsigned(2678, 12), 1617 => to_unsigned(3046, 12), 1618 => to_unsigned(1902, 12), 1619 => to_unsigned(15, 12), 1620 => to_unsigned(2328, 12), 1621 => to_unsigned(3994, 12), 1622 => to_unsigned(2405, 12), 1623 => to_unsigned(929, 12), 1624 => to_unsigned(917, 12), 1625 => to_unsigned(3378, 12), 1626 => to_unsigned(582, 12), 1627 => to_unsigned(2067, 12), 1628 => to_unsigned(3337, 12), 1629 => to_unsigned(108, 12), 1630 => to_unsigned(2260, 12), 1631 => to_unsigned(3211, 12), 1632 => to_unsigned(1307, 12), 1633 => to_unsigned(1176, 12), 1634 => to_unsigned(1130, 12), 1635 => to_unsigned(2104, 12), 1636 => to_unsigned(2767, 12), 1637 => to_unsigned(800, 12), 1638 => to_unsigned(3196, 12), 1639 => to_unsigned(3373, 12), 1640 => to_unsigned(1391, 12), 1641 => to_unsigned(2919, 12), 1642 => to_unsigned(3668, 12), 1643 => to_unsigned(3874, 12), 1644 => to_unsigned(451, 12), 1645 => to_unsigned(994, 12), 1646 => to_unsigned(3042, 12), 1647 => to_unsigned(3978, 12), 1648 => to_unsigned(2248, 12), 1649 => to_unsigned(1477, 12), 1650 => to_unsigned(2451, 12), 1651 => to_unsigned(1975, 12), 1652 => to_unsigned(3778, 12), 1653 => to_unsigned(3765, 12), 1654 => to_unsigned(823, 12), 1655 => to_unsigned(2952, 12), 1656 => to_unsigned(2555, 12), 1657 => to_unsigned(2493, 12), 1658 => to_unsigned(2107, 12), 1659 => to_unsigned(3248, 12), 1660 => to_unsigned(2220, 12), 1661 => to_unsigned(2806, 12), 1662 => to_unsigned(1325, 12), 1663 => to_unsigned(3754, 12), 1664 => to_unsigned(1585, 12), 1665 => to_unsigned(3845, 12), 1666 => to_unsigned(2270, 12), 1667 => to_unsigned(206, 12), 1668 => to_unsigned(2572, 12), 1669 => to_unsigned(291, 12), 1670 => to_unsigned(2761, 12), 1671 => to_unsigned(3386, 12), 1672 => to_unsigned(1456, 12), 1673 => to_unsigned(2667, 12), 1674 => to_unsigned(235, 12), 1675 => to_unsigned(1815, 12), 1676 => to_unsigned(2749, 12), 1677 => to_unsigned(1485, 12), 1678 => to_unsigned(460, 12), 1679 => to_unsigned(2641, 12), 1680 => to_unsigned(2632, 12), 1681 => to_unsigned(2068, 12), 1682 => to_unsigned(209, 12), 1683 => to_unsigned(2148, 12), 1684 => to_unsigned(2009, 12), 1685 => to_unsigned(1841, 12), 1686 => to_unsigned(2421, 12), 1687 => to_unsigned(1962, 12), 1688 => to_unsigned(1290, 12), 1689 => to_unsigned(547, 12), 1690 => to_unsigned(577, 12), 1691 => to_unsigned(3593, 12), 1692 => to_unsigned(174, 12), 1693 => to_unsigned(2886, 12), 1694 => to_unsigned(2318, 12), 1695 => to_unsigned(1735, 12), 1696 => to_unsigned(2902, 12), 1697 => to_unsigned(2265, 12), 1698 => to_unsigned(133, 12), 1699 => to_unsigned(3655, 12), 1700 => to_unsigned(730, 12), 1701 => to_unsigned(3564, 12), 1702 => to_unsigned(2561, 12), 1703 => to_unsigned(4084, 12), 1704 => to_unsigned(1223, 12), 1705 => to_unsigned(3237, 12), 1706 => to_unsigned(2340, 12), 1707 => to_unsigned(650, 12), 1708 => to_unsigned(258, 12), 1709 => to_unsigned(2411, 12), 1710 => to_unsigned(1177, 12), 1711 => to_unsigned(879, 12), 1712 => to_unsigned(1324, 12), 1713 => to_unsigned(1246, 12), 1714 => to_unsigned(2930, 12), 1715 => to_unsigned(583, 12), 1716 => to_unsigned(674, 12), 1717 => to_unsigned(3772, 12), 1718 => to_unsigned(3081, 12), 1719 => to_unsigned(2022, 12), 1720 => to_unsigned(1037, 12), 1721 => to_unsigned(3621, 12), 1722 => to_unsigned(2166, 12), 1723 => to_unsigned(4021, 12), 1724 => to_unsigned(445, 12), 1725 => to_unsigned(1877, 12), 1726 => to_unsigned(915, 12), 1727 => to_unsigned(3194, 12), 1728 => to_unsigned(3792, 12), 1729 => to_unsigned(235, 12), 1730 => to_unsigned(2315, 12), 1731 => to_unsigned(3161, 12), 1732 => to_unsigned(3207, 12), 1733 => to_unsigned(2402, 12), 1734 => to_unsigned(178, 12), 1735 => to_unsigned(1562, 12), 1736 => to_unsigned(2653, 12), 1737 => to_unsigned(3017, 12), 1738 => to_unsigned(1161, 12), 1739 => to_unsigned(1206, 12), 1740 => to_unsigned(3506, 12), 1741 => to_unsigned(1034, 12), 1742 => to_unsigned(77, 12), 1743 => to_unsigned(1778, 12), 1744 => to_unsigned(1259, 12), 1745 => to_unsigned(238, 12), 1746 => to_unsigned(1588, 12), 1747 => to_unsigned(2228, 12), 1748 => to_unsigned(3505, 12), 1749 => to_unsigned(2775, 12), 1750 => to_unsigned(1129, 12), 1751 => to_unsigned(3804, 12), 1752 => to_unsigned(77, 12), 1753 => to_unsigned(3414, 12), 1754 => to_unsigned(1527, 12), 1755 => to_unsigned(750, 12), 1756 => to_unsigned(482, 12), 1757 => to_unsigned(1898, 12), 1758 => to_unsigned(2403, 12), 1759 => to_unsigned(87, 12), 1760 => to_unsigned(1742, 12), 1761 => to_unsigned(919, 12), 1762 => to_unsigned(2928, 12), 1763 => to_unsigned(37, 12), 1764 => to_unsigned(1310, 12), 1765 => to_unsigned(3246, 12), 1766 => to_unsigned(1247, 12), 1767 => to_unsigned(1955, 12), 1768 => to_unsigned(3755, 12), 1769 => to_unsigned(647, 12), 1770 => to_unsigned(3602, 12), 1771 => to_unsigned(799, 12), 1772 => to_unsigned(3206, 12), 1773 => to_unsigned(335, 12), 1774 => to_unsigned(99, 12), 1775 => to_unsigned(2489, 12), 1776 => to_unsigned(4069, 12), 1777 => to_unsigned(2431, 12), 1778 => to_unsigned(2870, 12), 1779 => to_unsigned(2320, 12), 1780 => to_unsigned(246, 12), 1781 => to_unsigned(2749, 12), 1782 => to_unsigned(3243, 12), 1783 => to_unsigned(2241, 12), 1784 => to_unsigned(1958, 12), 1785 => to_unsigned(1737, 12), 1786 => to_unsigned(889, 12), 1787 => to_unsigned(3139, 12), 1788 => to_unsigned(1495, 12), 1789 => to_unsigned(1605, 12), 1790 => to_unsigned(1344, 12), 1791 => to_unsigned(1862, 12), 1792 => to_unsigned(1346, 12), 1793 => to_unsigned(3271, 12), 1794 => to_unsigned(3703, 12), 1795 => to_unsigned(3057, 12), 1796 => to_unsigned(1815, 12), 1797 => to_unsigned(1776, 12), 1798 => to_unsigned(352, 12), 1799 => to_unsigned(100, 12), 1800 => to_unsigned(1599, 12), 1801 => to_unsigned(122, 12), 1802 => to_unsigned(3879, 12), 1803 => to_unsigned(582, 12), 1804 => to_unsigned(1800, 12), 1805 => to_unsigned(1106, 12), 1806 => to_unsigned(3320, 12), 1807 => to_unsigned(1158, 12), 1808 => to_unsigned(1056, 12), 1809 => to_unsigned(239, 12), 1810 => to_unsigned(819, 12), 1811 => to_unsigned(3199, 12), 1812 => to_unsigned(3086, 12), 1813 => to_unsigned(2410, 12), 1814 => to_unsigned(287, 12), 1815 => to_unsigned(1507, 12), 1816 => to_unsigned(2042, 12), 1817 => to_unsigned(1753, 12), 1818 => to_unsigned(3315, 12), 1819 => to_unsigned(1932, 12), 1820 => to_unsigned(3480, 12), 1821 => to_unsigned(52, 12), 1822 => to_unsigned(3055, 12), 1823 => to_unsigned(3517, 12), 1824 => to_unsigned(2354, 12), 1825 => to_unsigned(78, 12), 1826 => to_unsigned(3465, 12), 1827 => to_unsigned(1686, 12), 1828 => to_unsigned(3404, 12), 1829 => to_unsigned(3109, 12), 1830 => to_unsigned(1121, 12), 1831 => to_unsigned(2500, 12), 1832 => to_unsigned(2430, 12), 1833 => to_unsigned(2989, 12), 1834 => to_unsigned(814, 12), 1835 => to_unsigned(3091, 12), 1836 => to_unsigned(3112, 12), 1837 => to_unsigned(3908, 12), 1838 => to_unsigned(2698, 12), 1839 => to_unsigned(267, 12), 1840 => to_unsigned(1652, 12), 1841 => to_unsigned(2487, 12), 1842 => to_unsigned(3467, 12), 1843 => to_unsigned(2289, 12), 1844 => to_unsigned(3329, 12), 1845 => to_unsigned(2021, 12), 1846 => to_unsigned(836, 12), 1847 => to_unsigned(2377, 12), 1848 => to_unsigned(2926, 12), 1849 => to_unsigned(2162, 12), 1850 => to_unsigned(1115, 12), 1851 => to_unsigned(495, 12), 1852 => to_unsigned(2783, 12), 1853 => to_unsigned(2356, 12), 1854 => to_unsigned(302, 12), 1855 => to_unsigned(884, 12), 1856 => to_unsigned(1876, 12), 1857 => to_unsigned(1811, 12), 1858 => to_unsigned(421, 12), 1859 => to_unsigned(3483, 12), 1860 => to_unsigned(3894, 12), 1861 => to_unsigned(2838, 12), 1862 => to_unsigned(1567, 12), 1863 => to_unsigned(3867, 12), 1864 => to_unsigned(898, 12), 1865 => to_unsigned(2101, 12), 1866 => to_unsigned(625, 12), 1867 => to_unsigned(2338, 12), 1868 => to_unsigned(3664, 12), 1869 => to_unsigned(2962, 12), 1870 => to_unsigned(2217, 12), 1871 => to_unsigned(1958, 12), 1872 => to_unsigned(1731, 12), 1873 => to_unsigned(4001, 12), 1874 => to_unsigned(583, 12), 1875 => to_unsigned(2706, 12), 1876 => to_unsigned(755, 12), 1877 => to_unsigned(3827, 12), 1878 => to_unsigned(1350, 12), 1879 => to_unsigned(262, 12), 1880 => to_unsigned(2350, 12), 1881 => to_unsigned(983, 12), 1882 => to_unsigned(2264, 12), 1883 => to_unsigned(1728, 12), 1884 => to_unsigned(100, 12), 1885 => to_unsigned(1187, 12), 1886 => to_unsigned(898, 12), 1887 => to_unsigned(636, 12), 1888 => to_unsigned(828, 12), 1889 => to_unsigned(945, 12), 1890 => to_unsigned(3989, 12), 1891 => to_unsigned(3902, 12), 1892 => to_unsigned(1012, 12), 1893 => to_unsigned(942, 12), 1894 => to_unsigned(3913, 12), 1895 => to_unsigned(2709, 12), 1896 => to_unsigned(1600, 12), 1897 => to_unsigned(827, 12), 1898 => to_unsigned(2688, 12), 1899 => to_unsigned(3369, 12), 1900 => to_unsigned(4075, 12), 1901 => to_unsigned(2878, 12), 1902 => to_unsigned(1059, 12), 1903 => to_unsigned(3827, 12), 1904 => to_unsigned(3957, 12), 1905 => to_unsigned(3487, 12), 1906 => to_unsigned(3524, 12), 1907 => to_unsigned(2376, 12), 1908 => to_unsigned(3312, 12), 1909 => to_unsigned(3496, 12), 1910 => to_unsigned(710, 12), 1911 => to_unsigned(3791, 12), 1912 => to_unsigned(628, 12), 1913 => to_unsigned(1276, 12), 1914 => to_unsigned(2020, 12), 1915 => to_unsigned(662, 12), 1916 => to_unsigned(341, 12), 1917 => to_unsigned(2989, 12), 1918 => to_unsigned(1427, 12), 1919 => to_unsigned(2104, 12), 1920 => to_unsigned(3222, 12), 1921 => to_unsigned(2631, 12), 1922 => to_unsigned(1995, 12), 1923 => to_unsigned(2294, 12), 1924 => to_unsigned(2831, 12), 1925 => to_unsigned(715, 12), 1926 => to_unsigned(3246, 12), 1927 => to_unsigned(561, 12), 1928 => to_unsigned(3593, 12), 1929 => to_unsigned(4064, 12), 1930 => to_unsigned(3875, 12), 1931 => to_unsigned(3761, 12), 1932 => to_unsigned(3746, 12), 1933 => to_unsigned(4, 12), 1934 => to_unsigned(1482, 12), 1935 => to_unsigned(1072, 12), 1936 => to_unsigned(2482, 12), 1937 => to_unsigned(53, 12), 1938 => to_unsigned(19, 12), 1939 => to_unsigned(2598, 12), 1940 => to_unsigned(2136, 12), 1941 => to_unsigned(3421, 12), 1942 => to_unsigned(2677, 12), 1943 => to_unsigned(1161, 12), 1944 => to_unsigned(1905, 12), 1945 => to_unsigned(3390, 12), 1946 => to_unsigned(2999, 12), 1947 => to_unsigned(1544, 12), 1948 => to_unsigned(695, 12), 1949 => to_unsigned(2260, 12), 1950 => to_unsigned(1397, 12), 1951 => to_unsigned(3722, 12), 1952 => to_unsigned(2345, 12), 1953 => to_unsigned(2926, 12), 1954 => to_unsigned(1861, 12), 1955 => to_unsigned(590, 12), 1956 => to_unsigned(601, 12), 1957 => to_unsigned(2854, 12), 1958 => to_unsigned(1653, 12), 1959 => to_unsigned(430, 12), 1960 => to_unsigned(4, 12), 1961 => to_unsigned(3410, 12), 1962 => to_unsigned(970, 12), 1963 => to_unsigned(1399, 12), 1964 => to_unsigned(102, 12), 1965 => to_unsigned(1952, 12), 1966 => to_unsigned(2480, 12), 1967 => to_unsigned(1441, 12), 1968 => to_unsigned(862, 12), 1969 => to_unsigned(3537, 12), 1970 => to_unsigned(3333, 12), 1971 => to_unsigned(645, 12), 1972 => to_unsigned(3635, 12), 1973 => to_unsigned(3694, 12), 1974 => to_unsigned(2888, 12), 1975 => to_unsigned(3495, 12), 1976 => to_unsigned(1679, 12), 1977 => to_unsigned(671, 12), 1978 => to_unsigned(3254, 12), 1979 => to_unsigned(3032, 12), 1980 => to_unsigned(2019, 12), 1981 => to_unsigned(1700, 12), 1982 => to_unsigned(1572, 12), 1983 => to_unsigned(243, 12), 1984 => to_unsigned(3834, 12), 1985 => to_unsigned(1863, 12), 1986 => to_unsigned(1744, 12), 1987 => to_unsigned(1602, 12), 1988 => to_unsigned(1330, 12), 1989 => to_unsigned(1348, 12), 1990 => to_unsigned(3449, 12), 1991 => to_unsigned(2674, 12), 1992 => to_unsigned(3809, 12), 1993 => to_unsigned(3972, 12), 1994 => to_unsigned(1247, 12), 1995 => to_unsigned(3720, 12), 1996 => to_unsigned(1035, 12), 1997 => to_unsigned(4025, 12), 1998 => to_unsigned(2311, 12), 1999 => to_unsigned(1565, 12), 2000 => to_unsigned(4047, 12), 2001 => to_unsigned(1845, 12), 2002 => to_unsigned(3232, 12), 2003 => to_unsigned(2961, 12), 2004 => to_unsigned(3469, 12), 2005 => to_unsigned(2564, 12), 2006 => to_unsigned(3752, 12), 2007 => to_unsigned(421, 12), 2008 => to_unsigned(3680, 12), 2009 => to_unsigned(712, 12), 2010 => to_unsigned(1235, 12), 2011 => to_unsigned(450, 12), 2012 => to_unsigned(1606, 12), 2013 => to_unsigned(3503, 12), 2014 => to_unsigned(1264, 12), 2015 => to_unsigned(831, 12), 2016 => to_unsigned(1456, 12), 2017 => to_unsigned(3785, 12), 2018 => to_unsigned(2623, 12), 2019 => to_unsigned(2612, 12), 2020 => to_unsigned(1789, 12), 2021 => to_unsigned(1619, 12), 2022 => to_unsigned(3094, 12), 2023 => to_unsigned(746, 12), 2024 => to_unsigned(2630, 12), 2025 => to_unsigned(2320, 12), 2026 => to_unsigned(3179, 12), 2027 => to_unsigned(2573, 12), 2028 => to_unsigned(1391, 12), 2029 => to_unsigned(528, 12), 2030 => to_unsigned(2883, 12), 2031 => to_unsigned(3920, 12), 2032 => to_unsigned(3906, 12), 2033 => to_unsigned(2486, 12), 2034 => to_unsigned(49, 12), 2035 => to_unsigned(1035, 12), 2036 => to_unsigned(3696, 12), 2037 => to_unsigned(3469, 12), 2038 => to_unsigned(2705, 12), 2039 => to_unsigned(1450, 12), 2040 => to_unsigned(1671, 12), 2041 => to_unsigned(4029, 12), 2042 => to_unsigned(1919, 12), 2043 => to_unsigned(1591, 12), 2044 => to_unsigned(3505, 12), 2045 => to_unsigned(1487, 12), 2046 => to_unsigned(2774, 12), 2047 => to_unsigned(2234, 12)),
            2 => (0 => to_unsigned(2113, 12), 1 => to_unsigned(3129, 12), 2 => to_unsigned(971, 12), 3 => to_unsigned(2463, 12), 4 => to_unsigned(3490, 12), 5 => to_unsigned(3457, 12), 6 => to_unsigned(3688, 12), 7 => to_unsigned(1108, 12), 8 => to_unsigned(3989, 12), 9 => to_unsigned(1137, 12), 10 => to_unsigned(388, 12), 11 => to_unsigned(3762, 12), 12 => to_unsigned(1431, 12), 13 => to_unsigned(726, 12), 14 => to_unsigned(1762, 12), 15 => to_unsigned(3328, 12), 16 => to_unsigned(1539, 12), 17 => to_unsigned(3389, 12), 18 => to_unsigned(2751, 12), 19 => to_unsigned(2771, 12), 20 => to_unsigned(3131, 12), 21 => to_unsigned(803, 12), 22 => to_unsigned(1483, 12), 23 => to_unsigned(806, 12), 24 => to_unsigned(3547, 12), 25 => to_unsigned(2430, 12), 26 => to_unsigned(947, 12), 27 => to_unsigned(82, 12), 28 => to_unsigned(1496, 12), 29 => to_unsigned(330, 12), 30 => to_unsigned(2849, 12), 31 => to_unsigned(2833, 12), 32 => to_unsigned(3795, 12), 33 => to_unsigned(2095, 12), 34 => to_unsigned(611, 12), 35 => to_unsigned(3890, 12), 36 => to_unsigned(2229, 12), 37 => to_unsigned(1459, 12), 38 => to_unsigned(4063, 12), 39 => to_unsigned(1735, 12), 40 => to_unsigned(4071, 12), 41 => to_unsigned(103, 12), 42 => to_unsigned(1611, 12), 43 => to_unsigned(4070, 12), 44 => to_unsigned(451, 12), 45 => to_unsigned(3130, 12), 46 => to_unsigned(3345, 12), 47 => to_unsigned(3886, 12), 48 => to_unsigned(3617, 12), 49 => to_unsigned(1345, 12), 50 => to_unsigned(2014, 12), 51 => to_unsigned(2012, 12), 52 => to_unsigned(2279, 12), 53 => to_unsigned(756, 12), 54 => to_unsigned(2550, 12), 55 => to_unsigned(3958, 12), 56 => to_unsigned(3568, 12), 57 => to_unsigned(3265, 12), 58 => to_unsigned(188, 12), 59 => to_unsigned(1513, 12), 60 => to_unsigned(935, 12), 61 => to_unsigned(2795, 12), 62 => to_unsigned(299, 12), 63 => to_unsigned(751, 12), 64 => to_unsigned(3365, 12), 65 => to_unsigned(3330, 12), 66 => to_unsigned(4038, 12), 67 => to_unsigned(40, 12), 68 => to_unsigned(2460, 12), 69 => to_unsigned(2712, 12), 70 => to_unsigned(2323, 12), 71 => to_unsigned(552, 12), 72 => to_unsigned(1167, 12), 73 => to_unsigned(2202, 12), 74 => to_unsigned(3763, 12), 75 => to_unsigned(539, 12), 76 => to_unsigned(1258, 12), 77 => to_unsigned(3644, 12), 78 => to_unsigned(3513, 12), 79 => to_unsigned(3697, 12), 80 => to_unsigned(960, 12), 81 => to_unsigned(1898, 12), 82 => to_unsigned(1179, 12), 83 => to_unsigned(3497, 12), 84 => to_unsigned(2592, 12), 85 => to_unsigned(2938, 12), 86 => to_unsigned(732, 12), 87 => to_unsigned(1224, 12), 88 => to_unsigned(1385, 12), 89 => to_unsigned(395, 12), 90 => to_unsigned(307, 12), 91 => to_unsigned(2631, 12), 92 => to_unsigned(2096, 12), 93 => to_unsigned(1788, 12), 94 => to_unsigned(1518, 12), 95 => to_unsigned(785, 12), 96 => to_unsigned(2658, 12), 97 => to_unsigned(2503, 12), 98 => to_unsigned(984, 12), 99 => to_unsigned(396, 12), 100 => to_unsigned(2000, 12), 101 => to_unsigned(919, 12), 102 => to_unsigned(149, 12), 103 => to_unsigned(3787, 12), 104 => to_unsigned(3178, 12), 105 => to_unsigned(2143, 12), 106 => to_unsigned(2125, 12), 107 => to_unsigned(923, 12), 108 => to_unsigned(2468, 12), 109 => to_unsigned(2229, 12), 110 => to_unsigned(3837, 12), 111 => to_unsigned(2510, 12), 112 => to_unsigned(2370, 12), 113 => to_unsigned(2698, 12), 114 => to_unsigned(420, 12), 115 => to_unsigned(2134, 12), 116 => to_unsigned(2472, 12), 117 => to_unsigned(1979, 12), 118 => to_unsigned(1224, 12), 119 => to_unsigned(1703, 12), 120 => to_unsigned(1258, 12), 121 => to_unsigned(2781, 12), 122 => to_unsigned(604, 12), 123 => to_unsigned(1811, 12), 124 => to_unsigned(1044, 12), 125 => to_unsigned(2012, 12), 126 => to_unsigned(389, 12), 127 => to_unsigned(3244, 12), 128 => to_unsigned(345, 12), 129 => to_unsigned(2097, 12), 130 => to_unsigned(844, 12), 131 => to_unsigned(3509, 12), 132 => to_unsigned(1385, 12), 133 => to_unsigned(2773, 12), 134 => to_unsigned(2528, 12), 135 => to_unsigned(1661, 12), 136 => to_unsigned(3763, 12), 137 => to_unsigned(3203, 12), 138 => to_unsigned(3122, 12), 139 => to_unsigned(859, 12), 140 => to_unsigned(2809, 12), 141 => to_unsigned(3933, 12), 142 => to_unsigned(3699, 12), 143 => to_unsigned(3209, 12), 144 => to_unsigned(4001, 12), 145 => to_unsigned(2119, 12), 146 => to_unsigned(1840, 12), 147 => to_unsigned(4092, 12), 148 => to_unsigned(2947, 12), 149 => to_unsigned(1819, 12), 150 => to_unsigned(1021, 12), 151 => to_unsigned(3585, 12), 152 => to_unsigned(1366, 12), 153 => to_unsigned(1950, 12), 154 => to_unsigned(2074, 12), 155 => to_unsigned(769, 12), 156 => to_unsigned(3099, 12), 157 => to_unsigned(2615, 12), 158 => to_unsigned(996, 12), 159 => to_unsigned(3135, 12), 160 => to_unsigned(1609, 12), 161 => to_unsigned(1480, 12), 162 => to_unsigned(1655, 12), 163 => to_unsigned(2357, 12), 164 => to_unsigned(3871, 12), 165 => to_unsigned(2077, 12), 166 => to_unsigned(1047, 12), 167 => to_unsigned(3146, 12), 168 => to_unsigned(3861, 12), 169 => to_unsigned(66, 12), 170 => to_unsigned(2690, 12), 171 => to_unsigned(2253, 12), 172 => to_unsigned(2458, 12), 173 => to_unsigned(2769, 12), 174 => to_unsigned(3518, 12), 175 => to_unsigned(482, 12), 176 => to_unsigned(884, 12), 177 => to_unsigned(3818, 12), 178 => to_unsigned(780, 12), 179 => to_unsigned(2748, 12), 180 => to_unsigned(3641, 12), 181 => to_unsigned(113, 12), 182 => to_unsigned(4082, 12), 183 => to_unsigned(158, 12), 184 => to_unsigned(2091, 12), 185 => to_unsigned(2565, 12), 186 => to_unsigned(2062, 12), 187 => to_unsigned(917, 12), 188 => to_unsigned(541, 12), 189 => to_unsigned(447, 12), 190 => to_unsigned(4021, 12), 191 => to_unsigned(3213, 12), 192 => to_unsigned(3805, 12), 193 => to_unsigned(1585, 12), 194 => to_unsigned(1219, 12), 195 => to_unsigned(3817, 12), 196 => to_unsigned(1339, 12), 197 => to_unsigned(3812, 12), 198 => to_unsigned(2040, 12), 199 => to_unsigned(1815, 12), 200 => to_unsigned(3097, 12), 201 => to_unsigned(487, 12), 202 => to_unsigned(672, 12), 203 => to_unsigned(1638, 12), 204 => to_unsigned(1409, 12), 205 => to_unsigned(3891, 12), 206 => to_unsigned(784, 12), 207 => to_unsigned(3150, 12), 208 => to_unsigned(2692, 12), 209 => to_unsigned(3808, 12), 210 => to_unsigned(2056, 12), 211 => to_unsigned(726, 12), 212 => to_unsigned(3077, 12), 213 => to_unsigned(64, 12), 214 => to_unsigned(2026, 12), 215 => to_unsigned(2773, 12), 216 => to_unsigned(3769, 12), 217 => to_unsigned(2317, 12), 218 => to_unsigned(63, 12), 219 => to_unsigned(1635, 12), 220 => to_unsigned(2238, 12), 221 => to_unsigned(3320, 12), 222 => to_unsigned(2275, 12), 223 => to_unsigned(928, 12), 224 => to_unsigned(3826, 12), 225 => to_unsigned(507, 12), 226 => to_unsigned(3287, 12), 227 => to_unsigned(3764, 12), 228 => to_unsigned(1366, 12), 229 => to_unsigned(924, 12), 230 => to_unsigned(3711, 12), 231 => to_unsigned(3212, 12), 232 => to_unsigned(3210, 12), 233 => to_unsigned(39, 12), 234 => to_unsigned(147, 12), 235 => to_unsigned(715, 12), 236 => to_unsigned(747, 12), 237 => to_unsigned(737, 12), 238 => to_unsigned(1521, 12), 239 => to_unsigned(2197, 12), 240 => to_unsigned(1436, 12), 241 => to_unsigned(1686, 12), 242 => to_unsigned(159, 12), 243 => to_unsigned(518, 12), 244 => to_unsigned(1285, 12), 245 => to_unsigned(1818, 12), 246 => to_unsigned(441, 12), 247 => to_unsigned(2525, 12), 248 => to_unsigned(3603, 12), 249 => to_unsigned(2133, 12), 250 => to_unsigned(2219, 12), 251 => to_unsigned(781, 12), 252 => to_unsigned(3188, 12), 253 => to_unsigned(1631, 12), 254 => to_unsigned(3086, 12), 255 => to_unsigned(2571, 12), 256 => to_unsigned(1527, 12), 257 => to_unsigned(1902, 12), 258 => to_unsigned(1736, 12), 259 => to_unsigned(4005, 12), 260 => to_unsigned(3313, 12), 261 => to_unsigned(3945, 12), 262 => to_unsigned(980, 12), 263 => to_unsigned(1553, 12), 264 => to_unsigned(3218, 12), 265 => to_unsigned(1204, 12), 266 => to_unsigned(3425, 12), 267 => to_unsigned(3728, 12), 268 => to_unsigned(3631, 12), 269 => to_unsigned(488, 12), 270 => to_unsigned(2555, 12), 271 => to_unsigned(92, 12), 272 => to_unsigned(2259, 12), 273 => to_unsigned(119, 12), 274 => to_unsigned(223, 12), 275 => to_unsigned(3569, 12), 276 => to_unsigned(2718, 12), 277 => to_unsigned(705, 12), 278 => to_unsigned(2834, 12), 279 => to_unsigned(1328, 12), 280 => to_unsigned(1591, 12), 281 => to_unsigned(700, 12), 282 => to_unsigned(803, 12), 283 => to_unsigned(2545, 12), 284 => to_unsigned(4094, 12), 285 => to_unsigned(3608, 12), 286 => to_unsigned(3281, 12), 287 => to_unsigned(87, 12), 288 => to_unsigned(3655, 12), 289 => to_unsigned(3319, 12), 290 => to_unsigned(2894, 12), 291 => to_unsigned(2828, 12), 292 => to_unsigned(3657, 12), 293 => to_unsigned(2580, 12), 294 => to_unsigned(1004, 12), 295 => to_unsigned(2736, 12), 296 => to_unsigned(1414, 12), 297 => to_unsigned(4048, 12), 298 => to_unsigned(1652, 12), 299 => to_unsigned(366, 12), 300 => to_unsigned(1043, 12), 301 => to_unsigned(1505, 12), 302 => to_unsigned(2575, 12), 303 => to_unsigned(17, 12), 304 => to_unsigned(2419, 12), 305 => to_unsigned(749, 12), 306 => to_unsigned(3185, 12), 307 => to_unsigned(1896, 12), 308 => to_unsigned(1122, 12), 309 => to_unsigned(3677, 12), 310 => to_unsigned(3774, 12), 311 => to_unsigned(442, 12), 312 => to_unsigned(1912, 12), 313 => to_unsigned(3927, 12), 314 => to_unsigned(355, 12), 315 => to_unsigned(3340, 12), 316 => to_unsigned(2994, 12), 317 => to_unsigned(3079, 12), 318 => to_unsigned(1303, 12), 319 => to_unsigned(3220, 12), 320 => to_unsigned(1475, 12), 321 => to_unsigned(2104, 12), 322 => to_unsigned(38, 12), 323 => to_unsigned(2927, 12), 324 => to_unsigned(3973, 12), 325 => to_unsigned(383, 12), 326 => to_unsigned(1776, 12), 327 => to_unsigned(3885, 12), 328 => to_unsigned(2856, 12), 329 => to_unsigned(256, 12), 330 => to_unsigned(1453, 12), 331 => to_unsigned(2457, 12), 332 => to_unsigned(1709, 12), 333 => to_unsigned(2749, 12), 334 => to_unsigned(3323, 12), 335 => to_unsigned(4021, 12), 336 => to_unsigned(675, 12), 337 => to_unsigned(2800, 12), 338 => to_unsigned(1931, 12), 339 => to_unsigned(973, 12), 340 => to_unsigned(2830, 12), 341 => to_unsigned(931, 12), 342 => to_unsigned(1655, 12), 343 => to_unsigned(3352, 12), 344 => to_unsigned(36, 12), 345 => to_unsigned(151, 12), 346 => to_unsigned(4089, 12), 347 => to_unsigned(786, 12), 348 => to_unsigned(2010, 12), 349 => to_unsigned(917, 12), 350 => to_unsigned(2317, 12), 351 => to_unsigned(3393, 12), 352 => to_unsigned(1762, 12), 353 => to_unsigned(3055, 12), 354 => to_unsigned(3159, 12), 355 => to_unsigned(2173, 12), 356 => to_unsigned(44, 12), 357 => to_unsigned(3670, 12), 358 => to_unsigned(2573, 12), 359 => to_unsigned(2990, 12), 360 => to_unsigned(3061, 12), 361 => to_unsigned(1006, 12), 362 => to_unsigned(1534, 12), 363 => to_unsigned(2240, 12), 364 => to_unsigned(2142, 12), 365 => to_unsigned(3858, 12), 366 => to_unsigned(2746, 12), 367 => to_unsigned(1320, 12), 368 => to_unsigned(2746, 12), 369 => to_unsigned(1799, 12), 370 => to_unsigned(1830, 12), 371 => to_unsigned(3545, 12), 372 => to_unsigned(2314, 12), 373 => to_unsigned(1890, 12), 374 => to_unsigned(1975, 12), 375 => to_unsigned(3177, 12), 376 => to_unsigned(3930, 12), 377 => to_unsigned(1971, 12), 378 => to_unsigned(3499, 12), 379 => to_unsigned(922, 12), 380 => to_unsigned(3271, 12), 381 => to_unsigned(414, 12), 382 => to_unsigned(105, 12), 383 => to_unsigned(2734, 12), 384 => to_unsigned(1335, 12), 385 => to_unsigned(1103, 12), 386 => to_unsigned(2601, 12), 387 => to_unsigned(3811, 12), 388 => to_unsigned(3924, 12), 389 => to_unsigned(608, 12), 390 => to_unsigned(2072, 12), 391 => to_unsigned(2415, 12), 392 => to_unsigned(3746, 12), 393 => to_unsigned(59, 12), 394 => to_unsigned(810, 12), 395 => to_unsigned(1287, 12), 396 => to_unsigned(1376, 12), 397 => to_unsigned(1146, 12), 398 => to_unsigned(1048, 12), 399 => to_unsigned(3855, 12), 400 => to_unsigned(2621, 12), 401 => to_unsigned(4076, 12), 402 => to_unsigned(2219, 12), 403 => to_unsigned(935, 12), 404 => to_unsigned(2322, 12), 405 => to_unsigned(3280, 12), 406 => to_unsigned(2239, 12), 407 => to_unsigned(2477, 12), 408 => to_unsigned(804, 12), 409 => to_unsigned(2673, 12), 410 => to_unsigned(1379, 12), 411 => to_unsigned(119, 12), 412 => to_unsigned(4042, 12), 413 => to_unsigned(734, 12), 414 => to_unsigned(316, 12), 415 => to_unsigned(2941, 12), 416 => to_unsigned(3238, 12), 417 => to_unsigned(3666, 12), 418 => to_unsigned(3531, 12), 419 => to_unsigned(1439, 12), 420 => to_unsigned(1172, 12), 421 => to_unsigned(2318, 12), 422 => to_unsigned(2471, 12), 423 => to_unsigned(3397, 12), 424 => to_unsigned(1814, 12), 425 => to_unsigned(2828, 12), 426 => to_unsigned(757, 12), 427 => to_unsigned(4053, 12), 428 => to_unsigned(3410, 12), 429 => to_unsigned(2881, 12), 430 => to_unsigned(2932, 12), 431 => to_unsigned(422, 12), 432 => to_unsigned(1687, 12), 433 => to_unsigned(3090, 12), 434 => to_unsigned(155, 12), 435 => to_unsigned(3376, 12), 436 => to_unsigned(820, 12), 437 => to_unsigned(3892, 12), 438 => to_unsigned(3569, 12), 439 => to_unsigned(2077, 12), 440 => to_unsigned(1687, 12), 441 => to_unsigned(2500, 12), 442 => to_unsigned(3476, 12), 443 => to_unsigned(3503, 12), 444 => to_unsigned(2792, 12), 445 => to_unsigned(203, 12), 446 => to_unsigned(2238, 12), 447 => to_unsigned(3973, 12), 448 => to_unsigned(175, 12), 449 => to_unsigned(1026, 12), 450 => to_unsigned(3029, 12), 451 => to_unsigned(3859, 12), 452 => to_unsigned(890, 12), 453 => to_unsigned(3563, 12), 454 => to_unsigned(3357, 12), 455 => to_unsigned(3040, 12), 456 => to_unsigned(1297, 12), 457 => to_unsigned(3579, 12), 458 => to_unsigned(305, 12), 459 => to_unsigned(376, 12), 460 => to_unsigned(441, 12), 461 => to_unsigned(3582, 12), 462 => to_unsigned(846, 12), 463 => to_unsigned(3297, 12), 464 => to_unsigned(574, 12), 465 => to_unsigned(3797, 12), 466 => to_unsigned(138, 12), 467 => to_unsigned(1939, 12), 468 => to_unsigned(3536, 12), 469 => to_unsigned(2238, 12), 470 => to_unsigned(3228, 12), 471 => to_unsigned(3238, 12), 472 => to_unsigned(1680, 12), 473 => to_unsigned(1192, 12), 474 => to_unsigned(2434, 12), 475 => to_unsigned(1420, 12), 476 => to_unsigned(578, 12), 477 => to_unsigned(1936, 12), 478 => to_unsigned(3045, 12), 479 => to_unsigned(4053, 12), 480 => to_unsigned(2406, 12), 481 => to_unsigned(2471, 12), 482 => to_unsigned(1791, 12), 483 => to_unsigned(137, 12), 484 => to_unsigned(281, 12), 485 => to_unsigned(688, 12), 486 => to_unsigned(974, 12), 487 => to_unsigned(333, 12), 488 => to_unsigned(115, 12), 489 => to_unsigned(2994, 12), 490 => to_unsigned(302, 12), 491 => to_unsigned(751, 12), 492 => to_unsigned(649, 12), 493 => to_unsigned(3262, 12), 494 => to_unsigned(1498, 12), 495 => to_unsigned(368, 12), 496 => to_unsigned(3700, 12), 497 => to_unsigned(83, 12), 498 => to_unsigned(3816, 12), 499 => to_unsigned(903, 12), 500 => to_unsigned(3277, 12), 501 => to_unsigned(3469, 12), 502 => to_unsigned(3226, 12), 503 => to_unsigned(3650, 12), 504 => to_unsigned(2892, 12), 505 => to_unsigned(1930, 12), 506 => to_unsigned(2043, 12), 507 => to_unsigned(1975, 12), 508 => to_unsigned(2689, 12), 509 => to_unsigned(3655, 12), 510 => to_unsigned(3199, 12), 511 => to_unsigned(1073, 12), 512 => to_unsigned(525, 12), 513 => to_unsigned(3028, 12), 514 => to_unsigned(2253, 12), 515 => to_unsigned(3499, 12), 516 => to_unsigned(1268, 12), 517 => to_unsigned(1889, 12), 518 => to_unsigned(3671, 12), 519 => to_unsigned(366, 12), 520 => to_unsigned(2994, 12), 521 => to_unsigned(2908, 12), 522 => to_unsigned(3363, 12), 523 => to_unsigned(1007, 12), 524 => to_unsigned(2794, 12), 525 => to_unsigned(3127, 12), 526 => to_unsigned(4020, 12), 527 => to_unsigned(4078, 12), 528 => to_unsigned(2403, 12), 529 => to_unsigned(2558, 12), 530 => to_unsigned(3994, 12), 531 => to_unsigned(655, 12), 532 => to_unsigned(1961, 12), 533 => to_unsigned(561, 12), 534 => to_unsigned(1917, 12), 535 => to_unsigned(2290, 12), 536 => to_unsigned(2155, 12), 537 => to_unsigned(1305, 12), 538 => to_unsigned(1644, 12), 539 => to_unsigned(1888, 12), 540 => to_unsigned(1756, 12), 541 => to_unsigned(2057, 12), 542 => to_unsigned(3499, 12), 543 => to_unsigned(65, 12), 544 => to_unsigned(104, 12), 545 => to_unsigned(681, 12), 546 => to_unsigned(1660, 12), 547 => to_unsigned(1169, 12), 548 => to_unsigned(3236, 12), 549 => to_unsigned(2463, 12), 550 => to_unsigned(1383, 12), 551 => to_unsigned(1928, 12), 552 => to_unsigned(1355, 12), 553 => to_unsigned(715, 12), 554 => to_unsigned(943, 12), 555 => to_unsigned(721, 12), 556 => to_unsigned(364, 12), 557 => to_unsigned(1527, 12), 558 => to_unsigned(1509, 12), 559 => to_unsigned(627, 12), 560 => to_unsigned(2164, 12), 561 => to_unsigned(701, 12), 562 => to_unsigned(1075, 12), 563 => to_unsigned(1093, 12), 564 => to_unsigned(3905, 12), 565 => to_unsigned(3278, 12), 566 => to_unsigned(3848, 12), 567 => to_unsigned(130, 12), 568 => to_unsigned(3792, 12), 569 => to_unsigned(2963, 12), 570 => to_unsigned(1336, 12), 571 => to_unsigned(2581, 12), 572 => to_unsigned(4015, 12), 573 => to_unsigned(2608, 12), 574 => to_unsigned(1887, 12), 575 => to_unsigned(2121, 12), 576 => to_unsigned(1478, 12), 577 => to_unsigned(1917, 12), 578 => to_unsigned(1824, 12), 579 => to_unsigned(2113, 12), 580 => to_unsigned(2219, 12), 581 => to_unsigned(2099, 12), 582 => to_unsigned(93, 12), 583 => to_unsigned(2972, 12), 584 => to_unsigned(2142, 12), 585 => to_unsigned(3782, 12), 586 => to_unsigned(3297, 12), 587 => to_unsigned(4070, 12), 588 => to_unsigned(4032, 12), 589 => to_unsigned(3897, 12), 590 => to_unsigned(1205, 12), 591 => to_unsigned(532, 12), 592 => to_unsigned(1645, 12), 593 => to_unsigned(3261, 12), 594 => to_unsigned(1530, 12), 595 => to_unsigned(993, 12), 596 => to_unsigned(3009, 12), 597 => to_unsigned(1382, 12), 598 => to_unsigned(1106, 12), 599 => to_unsigned(463, 12), 600 => to_unsigned(3769, 12), 601 => to_unsigned(3730, 12), 602 => to_unsigned(161, 12), 603 => to_unsigned(194, 12), 604 => to_unsigned(3686, 12), 605 => to_unsigned(3457, 12), 606 => to_unsigned(2922, 12), 607 => to_unsigned(3931, 12), 608 => to_unsigned(3279, 12), 609 => to_unsigned(1284, 12), 610 => to_unsigned(2083, 12), 611 => to_unsigned(971, 12), 612 => to_unsigned(2435, 12), 613 => to_unsigned(3595, 12), 614 => to_unsigned(2290, 12), 615 => to_unsigned(3035, 12), 616 => to_unsigned(108, 12), 617 => to_unsigned(4062, 12), 618 => to_unsigned(3253, 12), 619 => to_unsigned(2601, 12), 620 => to_unsigned(242, 12), 621 => to_unsigned(1310, 12), 622 => to_unsigned(1775, 12), 623 => to_unsigned(3054, 12), 624 => to_unsigned(654, 12), 625 => to_unsigned(3301, 12), 626 => to_unsigned(2702, 12), 627 => to_unsigned(1584, 12), 628 => to_unsigned(1927, 12), 629 => to_unsigned(1754, 12), 630 => to_unsigned(849, 12), 631 => to_unsigned(2528, 12), 632 => to_unsigned(3036, 12), 633 => to_unsigned(1898, 12), 634 => to_unsigned(2918, 12), 635 => to_unsigned(2870, 12), 636 => to_unsigned(3551, 12), 637 => to_unsigned(1121, 12), 638 => to_unsigned(3650, 12), 639 => to_unsigned(1548, 12), 640 => to_unsigned(2358, 12), 641 => to_unsigned(1836, 12), 642 => to_unsigned(1838, 12), 643 => to_unsigned(2244, 12), 644 => to_unsigned(2028, 12), 645 => to_unsigned(27, 12), 646 => to_unsigned(2514, 12), 647 => to_unsigned(726, 12), 648 => to_unsigned(2942, 12), 649 => to_unsigned(3359, 12), 650 => to_unsigned(1452, 12), 651 => to_unsigned(3676, 12), 652 => to_unsigned(384, 12), 653 => to_unsigned(394, 12), 654 => to_unsigned(2377, 12), 655 => to_unsigned(406, 12), 656 => to_unsigned(3044, 12), 657 => to_unsigned(2233, 12), 658 => to_unsigned(1414, 12), 659 => to_unsigned(2640, 12), 660 => to_unsigned(3764, 12), 661 => to_unsigned(378, 12), 662 => to_unsigned(2418, 12), 663 => to_unsigned(2028, 12), 664 => to_unsigned(1532, 12), 665 => to_unsigned(210, 12), 666 => to_unsigned(164, 12), 667 => to_unsigned(71, 12), 668 => to_unsigned(1660, 12), 669 => to_unsigned(332, 12), 670 => to_unsigned(3371, 12), 671 => to_unsigned(3813, 12), 672 => to_unsigned(2050, 12), 673 => to_unsigned(3461, 12), 674 => to_unsigned(3190, 12), 675 => to_unsigned(2472, 12), 676 => to_unsigned(1377, 12), 677 => to_unsigned(2097, 12), 678 => to_unsigned(2059, 12), 679 => to_unsigned(2239, 12), 680 => to_unsigned(3581, 12), 681 => to_unsigned(380, 12), 682 => to_unsigned(1034, 12), 683 => to_unsigned(1802, 12), 684 => to_unsigned(1960, 12), 685 => to_unsigned(2467, 12), 686 => to_unsigned(3956, 12), 687 => to_unsigned(369, 12), 688 => to_unsigned(3084, 12), 689 => to_unsigned(4009, 12), 690 => to_unsigned(1534, 12), 691 => to_unsigned(2487, 12), 692 => to_unsigned(2467, 12), 693 => to_unsigned(503, 12), 694 => to_unsigned(4043, 12), 695 => to_unsigned(2907, 12), 696 => to_unsigned(2192, 12), 697 => to_unsigned(2432, 12), 698 => to_unsigned(1692, 12), 699 => to_unsigned(1392, 12), 700 => to_unsigned(1456, 12), 701 => to_unsigned(1903, 12), 702 => to_unsigned(1530, 12), 703 => to_unsigned(3404, 12), 704 => to_unsigned(2933, 12), 705 => to_unsigned(1405, 12), 706 => to_unsigned(741, 12), 707 => to_unsigned(919, 12), 708 => to_unsigned(1318, 12), 709 => to_unsigned(802, 12), 710 => to_unsigned(2945, 12), 711 => to_unsigned(1910, 12), 712 => to_unsigned(954, 12), 713 => to_unsigned(184, 12), 714 => to_unsigned(2094, 12), 715 => to_unsigned(1411, 12), 716 => to_unsigned(3496, 12), 717 => to_unsigned(1932, 12), 718 => to_unsigned(405, 12), 719 => to_unsigned(2368, 12), 720 => to_unsigned(3899, 12), 721 => to_unsigned(1811, 12), 722 => to_unsigned(3700, 12), 723 => to_unsigned(3040, 12), 724 => to_unsigned(685, 12), 725 => to_unsigned(2560, 12), 726 => to_unsigned(2834, 12), 727 => to_unsigned(2751, 12), 728 => to_unsigned(2487, 12), 729 => to_unsigned(465, 12), 730 => to_unsigned(153, 12), 731 => to_unsigned(2737, 12), 732 => to_unsigned(3717, 12), 733 => to_unsigned(904, 12), 734 => to_unsigned(1602, 12), 735 => to_unsigned(102, 12), 736 => to_unsigned(1735, 12), 737 => to_unsigned(58, 12), 738 => to_unsigned(3617, 12), 739 => to_unsigned(3824, 12), 740 => to_unsigned(278, 12), 741 => to_unsigned(905, 12), 742 => to_unsigned(3941, 12), 743 => to_unsigned(2387, 12), 744 => to_unsigned(694, 12), 745 => to_unsigned(2146, 12), 746 => to_unsigned(2428, 12), 747 => to_unsigned(4050, 12), 748 => to_unsigned(3397, 12), 749 => to_unsigned(327, 12), 750 => to_unsigned(3282, 12), 751 => to_unsigned(2185, 12), 752 => to_unsigned(2512, 12), 753 => to_unsigned(3713, 12), 754 => to_unsigned(3038, 12), 755 => to_unsigned(1881, 12), 756 => to_unsigned(2085, 12), 757 => to_unsigned(3384, 12), 758 => to_unsigned(3773, 12), 759 => to_unsigned(1206, 12), 760 => to_unsigned(333, 12), 761 => to_unsigned(217, 12), 762 => to_unsigned(159, 12), 763 => to_unsigned(3652, 12), 764 => to_unsigned(4066, 12), 765 => to_unsigned(4084, 12), 766 => to_unsigned(254, 12), 767 => to_unsigned(2632, 12), 768 => to_unsigned(2176, 12), 769 => to_unsigned(2443, 12), 770 => to_unsigned(17, 12), 771 => to_unsigned(1577, 12), 772 => to_unsigned(3879, 12), 773 => to_unsigned(379, 12), 774 => to_unsigned(3765, 12), 775 => to_unsigned(1135, 12), 776 => to_unsigned(267, 12), 777 => to_unsigned(1501, 12), 778 => to_unsigned(801, 12), 779 => to_unsigned(3901, 12), 780 => to_unsigned(1573, 12), 781 => to_unsigned(2047, 12), 782 => to_unsigned(3813, 12), 783 => to_unsigned(3701, 12), 784 => to_unsigned(2351, 12), 785 => to_unsigned(657, 12), 786 => to_unsigned(4006, 12), 787 => to_unsigned(3033, 12), 788 => to_unsigned(3654, 12), 789 => to_unsigned(3114, 12), 790 => to_unsigned(936, 12), 791 => to_unsigned(2646, 12), 792 => to_unsigned(386, 12), 793 => to_unsigned(3236, 12), 794 => to_unsigned(274, 12), 795 => to_unsigned(3420, 12), 796 => to_unsigned(1090, 12), 797 => to_unsigned(1281, 12), 798 => to_unsigned(1874, 12), 799 => to_unsigned(1938, 12), 800 => to_unsigned(876, 12), 801 => to_unsigned(1410, 12), 802 => to_unsigned(1172, 12), 803 => to_unsigned(1524, 12), 804 => to_unsigned(3791, 12), 805 => to_unsigned(2587, 12), 806 => to_unsigned(504, 12), 807 => to_unsigned(954, 12), 808 => to_unsigned(343, 12), 809 => to_unsigned(2249, 12), 810 => to_unsigned(563, 12), 811 => to_unsigned(1492, 12), 812 => to_unsigned(584, 12), 813 => to_unsigned(410, 12), 814 => to_unsigned(375, 12), 815 => to_unsigned(2244, 12), 816 => to_unsigned(1003, 12), 817 => to_unsigned(895, 12), 818 => to_unsigned(291, 12), 819 => to_unsigned(2441, 12), 820 => to_unsigned(2442, 12), 821 => to_unsigned(2072, 12), 822 => to_unsigned(553, 12), 823 => to_unsigned(1746, 12), 824 => to_unsigned(1105, 12), 825 => to_unsigned(1562, 12), 826 => to_unsigned(2595, 12), 827 => to_unsigned(3476, 12), 828 => to_unsigned(1880, 12), 829 => to_unsigned(3881, 12), 830 => to_unsigned(1382, 12), 831 => to_unsigned(2883, 12), 832 => to_unsigned(4086, 12), 833 => to_unsigned(1695, 12), 834 => to_unsigned(2553, 12), 835 => to_unsigned(2078, 12), 836 => to_unsigned(3769, 12), 837 => to_unsigned(325, 12), 838 => to_unsigned(3953, 12), 839 => to_unsigned(1894, 12), 840 => to_unsigned(2966, 12), 841 => to_unsigned(1515, 12), 842 => to_unsigned(2653, 12), 843 => to_unsigned(3510, 12), 844 => to_unsigned(4074, 12), 845 => to_unsigned(2031, 12), 846 => to_unsigned(1661, 12), 847 => to_unsigned(2031, 12), 848 => to_unsigned(312, 12), 849 => to_unsigned(633, 12), 850 => to_unsigned(2793, 12), 851 => to_unsigned(1245, 12), 852 => to_unsigned(695, 12), 853 => to_unsigned(3077, 12), 854 => to_unsigned(3196, 12), 855 => to_unsigned(55, 12), 856 => to_unsigned(1069, 12), 857 => to_unsigned(44, 12), 858 => to_unsigned(1228, 12), 859 => to_unsigned(1968, 12), 860 => to_unsigned(428, 12), 861 => to_unsigned(1096, 12), 862 => to_unsigned(3918, 12), 863 => to_unsigned(360, 12), 864 => to_unsigned(3380, 12), 865 => to_unsigned(530, 12), 866 => to_unsigned(1757, 12), 867 => to_unsigned(2538, 12), 868 => to_unsigned(806, 12), 869 => to_unsigned(3610, 12), 870 => to_unsigned(594, 12), 871 => to_unsigned(1162, 12), 872 => to_unsigned(3289, 12), 873 => to_unsigned(3714, 12), 874 => to_unsigned(823, 12), 875 => to_unsigned(2270, 12), 876 => to_unsigned(738, 12), 877 => to_unsigned(2329, 12), 878 => to_unsigned(1398, 12), 879 => to_unsigned(3078, 12), 880 => to_unsigned(2663, 12), 881 => to_unsigned(2287, 12), 882 => to_unsigned(290, 12), 883 => to_unsigned(1603, 12), 884 => to_unsigned(3084, 12), 885 => to_unsigned(1552, 12), 886 => to_unsigned(1940, 12), 887 => to_unsigned(1441, 12), 888 => to_unsigned(1483, 12), 889 => to_unsigned(625, 12), 890 => to_unsigned(3868, 12), 891 => to_unsigned(1753, 12), 892 => to_unsigned(103, 12), 893 => to_unsigned(2835, 12), 894 => to_unsigned(1254, 12), 895 => to_unsigned(2012, 12), 896 => to_unsigned(3626, 12), 897 => to_unsigned(694, 12), 898 => to_unsigned(3486, 12), 899 => to_unsigned(1076, 12), 900 => to_unsigned(203, 12), 901 => to_unsigned(1356, 12), 902 => to_unsigned(2540, 12), 903 => to_unsigned(890, 12), 904 => to_unsigned(1568, 12), 905 => to_unsigned(3611, 12), 906 => to_unsigned(300, 12), 907 => to_unsigned(303, 12), 908 => to_unsigned(3310, 12), 909 => to_unsigned(2094, 12), 910 => to_unsigned(1233, 12), 911 => to_unsigned(1870, 12), 912 => to_unsigned(2415, 12), 913 => to_unsigned(1347, 12), 914 => to_unsigned(3185, 12), 915 => to_unsigned(3128, 12), 916 => to_unsigned(3835, 12), 917 => to_unsigned(3137, 12), 918 => to_unsigned(2638, 12), 919 => to_unsigned(1189, 12), 920 => to_unsigned(3907, 12), 921 => to_unsigned(3069, 12), 922 => to_unsigned(154, 12), 923 => to_unsigned(37, 12), 924 => to_unsigned(976, 12), 925 => to_unsigned(2425, 12), 926 => to_unsigned(3096, 12), 927 => to_unsigned(1607, 12), 928 => to_unsigned(3056, 12), 929 => to_unsigned(3146, 12), 930 => to_unsigned(3958, 12), 931 => to_unsigned(489, 12), 932 => to_unsigned(829, 12), 933 => to_unsigned(1243, 12), 934 => to_unsigned(1919, 12), 935 => to_unsigned(3410, 12), 936 => to_unsigned(3655, 12), 937 => to_unsigned(4046, 12), 938 => to_unsigned(2827, 12), 939 => to_unsigned(3937, 12), 940 => to_unsigned(2216, 12), 941 => to_unsigned(1739, 12), 942 => to_unsigned(3791, 12), 943 => to_unsigned(1037, 12), 944 => to_unsigned(2318, 12), 945 => to_unsigned(3586, 12), 946 => to_unsigned(2662, 12), 947 => to_unsigned(2703, 12), 948 => to_unsigned(525, 12), 949 => to_unsigned(3048, 12), 950 => to_unsigned(425, 12), 951 => to_unsigned(650, 12), 952 => to_unsigned(1952, 12), 953 => to_unsigned(3822, 12), 954 => to_unsigned(39, 12), 955 => to_unsigned(39, 12), 956 => to_unsigned(1045, 12), 957 => to_unsigned(430, 12), 958 => to_unsigned(3701, 12), 959 => to_unsigned(149, 12), 960 => to_unsigned(2005, 12), 961 => to_unsigned(1845, 12), 962 => to_unsigned(4072, 12), 963 => to_unsigned(1127, 12), 964 => to_unsigned(3284, 12), 965 => to_unsigned(241, 12), 966 => to_unsigned(1356, 12), 967 => to_unsigned(3440, 12), 968 => to_unsigned(2767, 12), 969 => to_unsigned(3562, 12), 970 => to_unsigned(4071, 12), 971 => to_unsigned(2795, 12), 972 => to_unsigned(1596, 12), 973 => to_unsigned(67, 12), 974 => to_unsigned(3916, 12), 975 => to_unsigned(3077, 12), 976 => to_unsigned(938, 12), 977 => to_unsigned(2214, 12), 978 => to_unsigned(111, 12), 979 => to_unsigned(2200, 12), 980 => to_unsigned(255, 12), 981 => to_unsigned(1891, 12), 982 => to_unsigned(2591, 12), 983 => to_unsigned(851, 12), 984 => to_unsigned(627, 12), 985 => to_unsigned(987, 12), 986 => to_unsigned(1552, 12), 987 => to_unsigned(3787, 12), 988 => to_unsigned(104, 12), 989 => to_unsigned(3837, 12), 990 => to_unsigned(3967, 12), 991 => to_unsigned(1560, 12), 992 => to_unsigned(3824, 12), 993 => to_unsigned(1004, 12), 994 => to_unsigned(107, 12), 995 => to_unsigned(83, 12), 996 => to_unsigned(814, 12), 997 => to_unsigned(3732, 12), 998 => to_unsigned(1064, 12), 999 => to_unsigned(2309, 12), 1000 => to_unsigned(2954, 12), 1001 => to_unsigned(115, 12), 1002 => to_unsigned(1046, 12), 1003 => to_unsigned(1054, 12), 1004 => to_unsigned(3299, 12), 1005 => to_unsigned(2087, 12), 1006 => to_unsigned(2474, 12), 1007 => to_unsigned(3921, 12), 1008 => to_unsigned(1411, 12), 1009 => to_unsigned(432, 12), 1010 => to_unsigned(4005, 12), 1011 => to_unsigned(419, 12), 1012 => to_unsigned(578, 12), 1013 => to_unsigned(1008, 12), 1014 => to_unsigned(1156, 12), 1015 => to_unsigned(184, 12), 1016 => to_unsigned(1508, 12), 1017 => to_unsigned(1172, 12), 1018 => to_unsigned(3121, 12), 1019 => to_unsigned(317, 12), 1020 => to_unsigned(1556, 12), 1021 => to_unsigned(349, 12), 1022 => to_unsigned(504, 12), 1023 => to_unsigned(1231, 12), 1024 => to_unsigned(428, 12), 1025 => to_unsigned(2514, 12), 1026 => to_unsigned(1068, 12), 1027 => to_unsigned(548, 12), 1028 => to_unsigned(2113, 12), 1029 => to_unsigned(995, 12), 1030 => to_unsigned(524, 12), 1031 => to_unsigned(832, 12), 1032 => to_unsigned(2825, 12), 1033 => to_unsigned(398, 12), 1034 => to_unsigned(318, 12), 1035 => to_unsigned(610, 12), 1036 => to_unsigned(3022, 12), 1037 => to_unsigned(815, 12), 1038 => to_unsigned(2550, 12), 1039 => to_unsigned(571, 12), 1040 => to_unsigned(2952, 12), 1041 => to_unsigned(3253, 12), 1042 => to_unsigned(2565, 12), 1043 => to_unsigned(2602, 12), 1044 => to_unsigned(4001, 12), 1045 => to_unsigned(261, 12), 1046 => to_unsigned(2666, 12), 1047 => to_unsigned(163, 12), 1048 => to_unsigned(2567, 12), 1049 => to_unsigned(3108, 12), 1050 => to_unsigned(3387, 12), 1051 => to_unsigned(2195, 12), 1052 => to_unsigned(98, 12), 1053 => to_unsigned(1359, 12), 1054 => to_unsigned(3485, 12), 1055 => to_unsigned(3888, 12), 1056 => to_unsigned(2647, 12), 1057 => to_unsigned(3319, 12), 1058 => to_unsigned(691, 12), 1059 => to_unsigned(1373, 12), 1060 => to_unsigned(3930, 12), 1061 => to_unsigned(839, 12), 1062 => to_unsigned(1110, 12), 1063 => to_unsigned(3378, 12), 1064 => to_unsigned(2773, 12), 1065 => to_unsigned(2789, 12), 1066 => to_unsigned(2437, 12), 1067 => to_unsigned(3613, 12), 1068 => to_unsigned(1436, 12), 1069 => to_unsigned(3414, 12), 1070 => to_unsigned(2561, 12), 1071 => to_unsigned(3197, 12), 1072 => to_unsigned(452, 12), 1073 => to_unsigned(3959, 12), 1074 => to_unsigned(2098, 12), 1075 => to_unsigned(2774, 12), 1076 => to_unsigned(2756, 12), 1077 => to_unsigned(2926, 12), 1078 => to_unsigned(3340, 12), 1079 => to_unsigned(1739, 12), 1080 => to_unsigned(3111, 12), 1081 => to_unsigned(1246, 12), 1082 => to_unsigned(2924, 12), 1083 => to_unsigned(3095, 12), 1084 => to_unsigned(3214, 12), 1085 => to_unsigned(1138, 12), 1086 => to_unsigned(3741, 12), 1087 => to_unsigned(3518, 12), 1088 => to_unsigned(2350, 12), 1089 => to_unsigned(859, 12), 1090 => to_unsigned(3003, 12), 1091 => to_unsigned(3081, 12), 1092 => to_unsigned(606, 12), 1093 => to_unsigned(1095, 12), 1094 => to_unsigned(108, 12), 1095 => to_unsigned(3789, 12), 1096 => to_unsigned(632, 12), 1097 => to_unsigned(2846, 12), 1098 => to_unsigned(785, 12), 1099 => to_unsigned(2755, 12), 1100 => to_unsigned(2766, 12), 1101 => to_unsigned(1470, 12), 1102 => to_unsigned(1390, 12), 1103 => to_unsigned(2392, 12), 1104 => to_unsigned(400, 12), 1105 => to_unsigned(1777, 12), 1106 => to_unsigned(1183, 12), 1107 => to_unsigned(1536, 12), 1108 => to_unsigned(676, 12), 1109 => to_unsigned(2297, 12), 1110 => to_unsigned(677, 12), 1111 => to_unsigned(646, 12), 1112 => to_unsigned(3955, 12), 1113 => to_unsigned(2954, 12), 1114 => to_unsigned(708, 12), 1115 => to_unsigned(381, 12), 1116 => to_unsigned(1757, 12), 1117 => to_unsigned(3819, 12), 1118 => to_unsigned(1021, 12), 1119 => to_unsigned(1585, 12), 1120 => to_unsigned(3180, 12), 1121 => to_unsigned(2775, 12), 1122 => to_unsigned(1920, 12), 1123 => to_unsigned(1976, 12), 1124 => to_unsigned(2396, 12), 1125 => to_unsigned(2780, 12), 1126 => to_unsigned(1769, 12), 1127 => to_unsigned(3338, 12), 1128 => to_unsigned(3639, 12), 1129 => to_unsigned(3317, 12), 1130 => to_unsigned(632, 12), 1131 => to_unsigned(3074, 12), 1132 => to_unsigned(1692, 12), 1133 => to_unsigned(1516, 12), 1134 => to_unsigned(3924, 12), 1135 => to_unsigned(1889, 12), 1136 => to_unsigned(4037, 12), 1137 => to_unsigned(267, 12), 1138 => to_unsigned(4028, 12), 1139 => to_unsigned(785, 12), 1140 => to_unsigned(191, 12), 1141 => to_unsigned(3450, 12), 1142 => to_unsigned(2995, 12), 1143 => to_unsigned(3403, 12), 1144 => to_unsigned(2354, 12), 1145 => to_unsigned(2135, 12), 1146 => to_unsigned(210, 12), 1147 => to_unsigned(3685, 12), 1148 => to_unsigned(1423, 12), 1149 => to_unsigned(3496, 12), 1150 => to_unsigned(380, 12), 1151 => to_unsigned(3205, 12), 1152 => to_unsigned(612, 12), 1153 => to_unsigned(3554, 12), 1154 => to_unsigned(2322, 12), 1155 => to_unsigned(1085, 12), 1156 => to_unsigned(2742, 12), 1157 => to_unsigned(1348, 12), 1158 => to_unsigned(3988, 12), 1159 => to_unsigned(258, 12), 1160 => to_unsigned(621, 12), 1161 => to_unsigned(2323, 12), 1162 => to_unsigned(898, 12), 1163 => to_unsigned(3436, 12), 1164 => to_unsigned(3313, 12), 1165 => to_unsigned(3759, 12), 1166 => to_unsigned(3065, 12), 1167 => to_unsigned(1374, 12), 1168 => to_unsigned(353, 12), 1169 => to_unsigned(959, 12), 1170 => to_unsigned(1929, 12), 1171 => to_unsigned(1547, 12), 1172 => to_unsigned(3974, 12), 1173 => to_unsigned(1587, 12), 1174 => to_unsigned(462, 12), 1175 => to_unsigned(530, 12), 1176 => to_unsigned(325, 12), 1177 => to_unsigned(3932, 12), 1178 => to_unsigned(1916, 12), 1179 => to_unsigned(444, 12), 1180 => to_unsigned(3680, 12), 1181 => to_unsigned(879, 12), 1182 => to_unsigned(2, 12), 1183 => to_unsigned(3820, 12), 1184 => to_unsigned(3877, 12), 1185 => to_unsigned(3747, 12), 1186 => to_unsigned(3139, 12), 1187 => to_unsigned(3018, 12), 1188 => to_unsigned(91, 12), 1189 => to_unsigned(2909, 12), 1190 => to_unsigned(1603, 12), 1191 => to_unsigned(3135, 12), 1192 => to_unsigned(2397, 12), 1193 => to_unsigned(3908, 12), 1194 => to_unsigned(3745, 12), 1195 => to_unsigned(3449, 12), 1196 => to_unsigned(92, 12), 1197 => to_unsigned(3911, 12), 1198 => to_unsigned(4032, 12), 1199 => to_unsigned(2281, 12), 1200 => to_unsigned(2219, 12), 1201 => to_unsigned(2059, 12), 1202 => to_unsigned(3569, 12), 1203 => to_unsigned(1203, 12), 1204 => to_unsigned(779, 12), 1205 => to_unsigned(3670, 12), 1206 => to_unsigned(3000, 12), 1207 => to_unsigned(1316, 12), 1208 => to_unsigned(267, 12), 1209 => to_unsigned(2643, 12), 1210 => to_unsigned(1166, 12), 1211 => to_unsigned(3556, 12), 1212 => to_unsigned(3735, 12), 1213 => to_unsigned(3566, 12), 1214 => to_unsigned(2277, 12), 1215 => to_unsigned(978, 12), 1216 => to_unsigned(2590, 12), 1217 => to_unsigned(994, 12), 1218 => to_unsigned(2303, 12), 1219 => to_unsigned(1, 12), 1220 => to_unsigned(933, 12), 1221 => to_unsigned(3151, 12), 1222 => to_unsigned(1706, 12), 1223 => to_unsigned(2406, 12), 1224 => to_unsigned(1906, 12), 1225 => to_unsigned(1323, 12), 1226 => to_unsigned(185, 12), 1227 => to_unsigned(3104, 12), 1228 => to_unsigned(1517, 12), 1229 => to_unsigned(927, 12), 1230 => to_unsigned(3923, 12), 1231 => to_unsigned(1999, 12), 1232 => to_unsigned(1898, 12), 1233 => to_unsigned(9, 12), 1234 => to_unsigned(3335, 12), 1235 => to_unsigned(253, 12), 1236 => to_unsigned(1576, 12), 1237 => to_unsigned(2267, 12), 1238 => to_unsigned(3971, 12), 1239 => to_unsigned(4028, 12), 1240 => to_unsigned(1371, 12), 1241 => to_unsigned(3859, 12), 1242 => to_unsigned(2165, 12), 1243 => to_unsigned(2967, 12), 1244 => to_unsigned(41, 12), 1245 => to_unsigned(3051, 12), 1246 => to_unsigned(819, 12), 1247 => to_unsigned(2243, 12), 1248 => to_unsigned(1677, 12), 1249 => to_unsigned(2948, 12), 1250 => to_unsigned(2705, 12), 1251 => to_unsigned(776, 12), 1252 => to_unsigned(186, 12), 1253 => to_unsigned(509, 12), 1254 => to_unsigned(3222, 12), 1255 => to_unsigned(900, 12), 1256 => to_unsigned(1348, 12), 1257 => to_unsigned(1956, 12), 1258 => to_unsigned(49, 12), 1259 => to_unsigned(447, 12), 1260 => to_unsigned(2647, 12), 1261 => to_unsigned(1145, 12), 1262 => to_unsigned(1237, 12), 1263 => to_unsigned(1276, 12), 1264 => to_unsigned(3097, 12), 1265 => to_unsigned(1051, 12), 1266 => to_unsigned(1573, 12), 1267 => to_unsigned(457, 12), 1268 => to_unsigned(364, 12), 1269 => to_unsigned(3382, 12), 1270 => to_unsigned(2105, 12), 1271 => to_unsigned(2731, 12), 1272 => to_unsigned(3200, 12), 1273 => to_unsigned(1306, 12), 1274 => to_unsigned(1735, 12), 1275 => to_unsigned(3179, 12), 1276 => to_unsigned(2836, 12), 1277 => to_unsigned(1024, 12), 1278 => to_unsigned(1562, 12), 1279 => to_unsigned(339, 12), 1280 => to_unsigned(3348, 12), 1281 => to_unsigned(1669, 12), 1282 => to_unsigned(2275, 12), 1283 => to_unsigned(69, 12), 1284 => to_unsigned(876, 12), 1285 => to_unsigned(2018, 12), 1286 => to_unsigned(486, 12), 1287 => to_unsigned(2836, 12), 1288 => to_unsigned(2965, 12), 1289 => to_unsigned(4060, 12), 1290 => to_unsigned(1300, 12), 1291 => to_unsigned(3757, 12), 1292 => to_unsigned(2552, 12), 1293 => to_unsigned(300, 12), 1294 => to_unsigned(1389, 12), 1295 => to_unsigned(900, 12), 1296 => to_unsigned(861, 12), 1297 => to_unsigned(1600, 12), 1298 => to_unsigned(1590, 12), 1299 => to_unsigned(3710, 12), 1300 => to_unsigned(1060, 12), 1301 => to_unsigned(3527, 12), 1302 => to_unsigned(3992, 12), 1303 => to_unsigned(3170, 12), 1304 => to_unsigned(2897, 12), 1305 => to_unsigned(1953, 12), 1306 => to_unsigned(195, 12), 1307 => to_unsigned(2240, 12), 1308 => to_unsigned(3188, 12), 1309 => to_unsigned(680, 12), 1310 => to_unsigned(846, 12), 1311 => to_unsigned(1798, 12), 1312 => to_unsigned(1814, 12), 1313 => to_unsigned(2501, 12), 1314 => to_unsigned(3780, 12), 1315 => to_unsigned(3827, 12), 1316 => to_unsigned(2334, 12), 1317 => to_unsigned(1107, 12), 1318 => to_unsigned(2151, 12), 1319 => to_unsigned(3727, 12), 1320 => to_unsigned(3453, 12), 1321 => to_unsigned(314, 12), 1322 => to_unsigned(345, 12), 1323 => to_unsigned(1249, 12), 1324 => to_unsigned(2031, 12), 1325 => to_unsigned(149, 12), 1326 => to_unsigned(2347, 12), 1327 => to_unsigned(318, 12), 1328 => to_unsigned(3918, 12), 1329 => to_unsigned(178, 12), 1330 => to_unsigned(4077, 12), 1331 => to_unsigned(577, 12), 1332 => to_unsigned(3816, 12), 1333 => to_unsigned(1650, 12), 1334 => to_unsigned(2112, 12), 1335 => to_unsigned(827, 12), 1336 => to_unsigned(1548, 12), 1337 => to_unsigned(2997, 12), 1338 => to_unsigned(1256, 12), 1339 => to_unsigned(2500, 12), 1340 => to_unsigned(2096, 12), 1341 => to_unsigned(122, 12), 1342 => to_unsigned(3398, 12), 1343 => to_unsigned(505, 12), 1344 => to_unsigned(4012, 12), 1345 => to_unsigned(3277, 12), 1346 => to_unsigned(3704, 12), 1347 => to_unsigned(2681, 12), 1348 => to_unsigned(3255, 12), 1349 => to_unsigned(1503, 12), 1350 => to_unsigned(2974, 12), 1351 => to_unsigned(4073, 12), 1352 => to_unsigned(583, 12), 1353 => to_unsigned(3428, 12), 1354 => to_unsigned(2619, 12), 1355 => to_unsigned(2838, 12), 1356 => to_unsigned(3346, 12), 1357 => to_unsigned(623, 12), 1358 => to_unsigned(457, 12), 1359 => to_unsigned(2788, 12), 1360 => to_unsigned(1819, 12), 1361 => to_unsigned(2322, 12), 1362 => to_unsigned(2531, 12), 1363 => to_unsigned(2070, 12), 1364 => to_unsigned(3410, 12), 1365 => to_unsigned(3628, 12), 1366 => to_unsigned(1841, 12), 1367 => to_unsigned(2794, 12), 1368 => to_unsigned(1766, 12), 1369 => to_unsigned(3589, 12), 1370 => to_unsigned(4019, 12), 1371 => to_unsigned(3120, 12), 1372 => to_unsigned(1138, 12), 1373 => to_unsigned(1307, 12), 1374 => to_unsigned(3714, 12), 1375 => to_unsigned(2126, 12), 1376 => to_unsigned(304, 12), 1377 => to_unsigned(3161, 12), 1378 => to_unsigned(3777, 12), 1379 => to_unsigned(3231, 12), 1380 => to_unsigned(3811, 12), 1381 => to_unsigned(3958, 12), 1382 => to_unsigned(3605, 12), 1383 => to_unsigned(1888, 12), 1384 => to_unsigned(1223, 12), 1385 => to_unsigned(558, 12), 1386 => to_unsigned(3641, 12), 1387 => to_unsigned(842, 12), 1388 => to_unsigned(3849, 12), 1389 => to_unsigned(3760, 12), 1390 => to_unsigned(1334, 12), 1391 => to_unsigned(2587, 12), 1392 => to_unsigned(2939, 12), 1393 => to_unsigned(1440, 12), 1394 => to_unsigned(2446, 12), 1395 => to_unsigned(3041, 12), 1396 => to_unsigned(1543, 12), 1397 => to_unsigned(2021, 12), 1398 => to_unsigned(2174, 12), 1399 => to_unsigned(2213, 12), 1400 => to_unsigned(1423, 12), 1401 => to_unsigned(3427, 12), 1402 => to_unsigned(594, 12), 1403 => to_unsigned(1613, 12), 1404 => to_unsigned(98, 12), 1405 => to_unsigned(3727, 12), 1406 => to_unsigned(1260, 12), 1407 => to_unsigned(3031, 12), 1408 => to_unsigned(415, 12), 1409 => to_unsigned(3498, 12), 1410 => to_unsigned(1203, 12), 1411 => to_unsigned(3838, 12), 1412 => to_unsigned(2959, 12), 1413 => to_unsigned(3258, 12), 1414 => to_unsigned(1318, 12), 1415 => to_unsigned(163, 12), 1416 => to_unsigned(2442, 12), 1417 => to_unsigned(1065, 12), 1418 => to_unsigned(1623, 12), 1419 => to_unsigned(579, 12), 1420 => to_unsigned(3450, 12), 1421 => to_unsigned(2989, 12), 1422 => to_unsigned(3555, 12), 1423 => to_unsigned(1914, 12), 1424 => to_unsigned(3497, 12), 1425 => to_unsigned(2290, 12), 1426 => to_unsigned(2818, 12), 1427 => to_unsigned(3900, 12), 1428 => to_unsigned(530, 12), 1429 => to_unsigned(3173, 12), 1430 => to_unsigned(227, 12), 1431 => to_unsigned(1869, 12), 1432 => to_unsigned(1179, 12), 1433 => to_unsigned(1023, 12), 1434 => to_unsigned(704, 12), 1435 => to_unsigned(2455, 12), 1436 => to_unsigned(278, 12), 1437 => to_unsigned(2895, 12), 1438 => to_unsigned(1814, 12), 1439 => to_unsigned(2237, 12), 1440 => to_unsigned(2300, 12), 1441 => to_unsigned(235, 12), 1442 => to_unsigned(1677, 12), 1443 => to_unsigned(3666, 12), 1444 => to_unsigned(3179, 12), 1445 => to_unsigned(3736, 12), 1446 => to_unsigned(1504, 12), 1447 => to_unsigned(549, 12), 1448 => to_unsigned(733, 12), 1449 => to_unsigned(2780, 12), 1450 => to_unsigned(3545, 12), 1451 => to_unsigned(453, 12), 1452 => to_unsigned(679, 12), 1453 => to_unsigned(1596, 12), 1454 => to_unsigned(1982, 12), 1455 => to_unsigned(2277, 12), 1456 => to_unsigned(3179, 12), 1457 => to_unsigned(175, 12), 1458 => to_unsigned(4091, 12), 1459 => to_unsigned(2768, 12), 1460 => to_unsigned(163, 12), 1461 => to_unsigned(1129, 12), 1462 => to_unsigned(92, 12), 1463 => to_unsigned(2183, 12), 1464 => to_unsigned(2434, 12), 1465 => to_unsigned(2136, 12), 1466 => to_unsigned(607, 12), 1467 => to_unsigned(3209, 12), 1468 => to_unsigned(251, 12), 1469 => to_unsigned(427, 12), 1470 => to_unsigned(1146, 12), 1471 => to_unsigned(3889, 12), 1472 => to_unsigned(680, 12), 1473 => to_unsigned(1464, 12), 1474 => to_unsigned(597, 12), 1475 => to_unsigned(3124, 12), 1476 => to_unsigned(578, 12), 1477 => to_unsigned(605, 12), 1478 => to_unsigned(3604, 12), 1479 => to_unsigned(1203, 12), 1480 => to_unsigned(1390, 12), 1481 => to_unsigned(1854, 12), 1482 => to_unsigned(482, 12), 1483 => to_unsigned(2382, 12), 1484 => to_unsigned(812, 12), 1485 => to_unsigned(2820, 12), 1486 => to_unsigned(156, 12), 1487 => to_unsigned(2787, 12), 1488 => to_unsigned(1954, 12), 1489 => to_unsigned(3319, 12), 1490 => to_unsigned(435, 12), 1491 => to_unsigned(2884, 12), 1492 => to_unsigned(277, 12), 1493 => to_unsigned(3361, 12), 1494 => to_unsigned(1743, 12), 1495 => to_unsigned(2257, 12), 1496 => to_unsigned(802, 12), 1497 => to_unsigned(1826, 12), 1498 => to_unsigned(1654, 12), 1499 => to_unsigned(2532, 12), 1500 => to_unsigned(726, 12), 1501 => to_unsigned(3532, 12), 1502 => to_unsigned(3418, 12), 1503 => to_unsigned(1904, 12), 1504 => to_unsigned(1184, 12), 1505 => to_unsigned(3970, 12), 1506 => to_unsigned(2976, 12), 1507 => to_unsigned(2209, 12), 1508 => to_unsigned(2569, 12), 1509 => to_unsigned(2247, 12), 1510 => to_unsigned(2455, 12), 1511 => to_unsigned(3527, 12), 1512 => to_unsigned(1163, 12), 1513 => to_unsigned(1750, 12), 1514 => to_unsigned(3235, 12), 1515 => to_unsigned(1176, 12), 1516 => to_unsigned(1225, 12), 1517 => to_unsigned(4053, 12), 1518 => to_unsigned(3118, 12), 1519 => to_unsigned(2839, 12), 1520 => to_unsigned(2731, 12), 1521 => to_unsigned(23, 12), 1522 => to_unsigned(1368, 12), 1523 => to_unsigned(2182, 12), 1524 => to_unsigned(1940, 12), 1525 => to_unsigned(2532, 12), 1526 => to_unsigned(1326, 12), 1527 => to_unsigned(416, 12), 1528 => to_unsigned(3370, 12), 1529 => to_unsigned(3987, 12), 1530 => to_unsigned(2624, 12), 1531 => to_unsigned(446, 12), 1532 => to_unsigned(3844, 12), 1533 => to_unsigned(85, 12), 1534 => to_unsigned(1208, 12), 1535 => to_unsigned(2719, 12), 1536 => to_unsigned(3760, 12), 1537 => to_unsigned(2759, 12), 1538 => to_unsigned(1201, 12), 1539 => to_unsigned(3056, 12), 1540 => to_unsigned(1136, 12), 1541 => to_unsigned(1548, 12), 1542 => to_unsigned(3729, 12), 1543 => to_unsigned(3997, 12), 1544 => to_unsigned(1016, 12), 1545 => to_unsigned(179, 12), 1546 => to_unsigned(3459, 12), 1547 => to_unsigned(1182, 12), 1548 => to_unsigned(90, 12), 1549 => to_unsigned(1581, 12), 1550 => to_unsigned(2711, 12), 1551 => to_unsigned(377, 12), 1552 => to_unsigned(3553, 12), 1553 => to_unsigned(1745, 12), 1554 => to_unsigned(274, 12), 1555 => to_unsigned(1757, 12), 1556 => to_unsigned(2498, 12), 1557 => to_unsigned(3988, 12), 1558 => to_unsigned(3120, 12), 1559 => to_unsigned(3605, 12), 1560 => to_unsigned(1214, 12), 1561 => to_unsigned(1764, 12), 1562 => to_unsigned(285, 12), 1563 => to_unsigned(3396, 12), 1564 => to_unsigned(169, 12), 1565 => to_unsigned(2493, 12), 1566 => to_unsigned(286, 12), 1567 => to_unsigned(114, 12), 1568 => to_unsigned(3435, 12), 1569 => to_unsigned(3562, 12), 1570 => to_unsigned(2690, 12), 1571 => to_unsigned(3592, 12), 1572 => to_unsigned(2299, 12), 1573 => to_unsigned(1996, 12), 1574 => to_unsigned(3321, 12), 1575 => to_unsigned(3974, 12), 1576 => to_unsigned(3754, 12), 1577 => to_unsigned(4013, 12), 1578 => to_unsigned(3891, 12), 1579 => to_unsigned(1625, 12), 1580 => to_unsigned(932, 12), 1581 => to_unsigned(3479, 12), 1582 => to_unsigned(3200, 12), 1583 => to_unsigned(2416, 12), 1584 => to_unsigned(3585, 12), 1585 => to_unsigned(170, 12), 1586 => to_unsigned(2842, 12), 1587 => to_unsigned(2736, 12), 1588 => to_unsigned(1200, 12), 1589 => to_unsigned(3528, 12), 1590 => to_unsigned(1426, 12), 1591 => to_unsigned(3090, 12), 1592 => to_unsigned(269, 12), 1593 => to_unsigned(3207, 12), 1594 => to_unsigned(3436, 12), 1595 => to_unsigned(2789, 12), 1596 => to_unsigned(1411, 12), 1597 => to_unsigned(3476, 12), 1598 => to_unsigned(2998, 12), 1599 => to_unsigned(234, 12), 1600 => to_unsigned(2738, 12), 1601 => to_unsigned(2626, 12), 1602 => to_unsigned(3640, 12), 1603 => to_unsigned(3690, 12), 1604 => to_unsigned(1274, 12), 1605 => to_unsigned(2384, 12), 1606 => to_unsigned(1658, 12), 1607 => to_unsigned(1998, 12), 1608 => to_unsigned(235, 12), 1609 => to_unsigned(3055, 12), 1610 => to_unsigned(1977, 12), 1611 => to_unsigned(3828, 12), 1612 => to_unsigned(396, 12), 1613 => to_unsigned(2216, 12), 1614 => to_unsigned(755, 12), 1615 => to_unsigned(489, 12), 1616 => to_unsigned(1849, 12), 1617 => to_unsigned(1362, 12), 1618 => to_unsigned(915, 12), 1619 => to_unsigned(194, 12), 1620 => to_unsigned(1348, 12), 1621 => to_unsigned(4055, 12), 1622 => to_unsigned(1430, 12), 1623 => to_unsigned(1065, 12), 1624 => to_unsigned(2153, 12), 1625 => to_unsigned(1212, 12), 1626 => to_unsigned(2188, 12), 1627 => to_unsigned(3583, 12), 1628 => to_unsigned(2921, 12), 1629 => to_unsigned(1639, 12), 1630 => to_unsigned(3905, 12), 1631 => to_unsigned(1042, 12), 1632 => to_unsigned(2770, 12), 1633 => to_unsigned(131, 12), 1634 => to_unsigned(1599, 12), 1635 => to_unsigned(661, 12), 1636 => to_unsigned(1447, 12), 1637 => to_unsigned(1544, 12), 1638 => to_unsigned(1857, 12), 1639 => to_unsigned(3445, 12), 1640 => to_unsigned(1765, 12), 1641 => to_unsigned(1577, 12), 1642 => to_unsigned(1184, 12), 1643 => to_unsigned(950, 12), 1644 => to_unsigned(3632, 12), 1645 => to_unsigned(3474, 12), 1646 => to_unsigned(799, 12), 1647 => to_unsigned(1634, 12), 1648 => to_unsigned(1892, 12), 1649 => to_unsigned(3959, 12), 1650 => to_unsigned(3507, 12), 1651 => to_unsigned(2551, 12), 1652 => to_unsigned(2748, 12), 1653 => to_unsigned(3938, 12), 1654 => to_unsigned(3855, 12), 1655 => to_unsigned(276, 12), 1656 => to_unsigned(1169, 12), 1657 => to_unsigned(3751, 12), 1658 => to_unsigned(2370, 12), 1659 => to_unsigned(1997, 12), 1660 => to_unsigned(3134, 12), 1661 => to_unsigned(612, 12), 1662 => to_unsigned(2060, 12), 1663 => to_unsigned(1967, 12), 1664 => to_unsigned(1902, 12), 1665 => to_unsigned(1954, 12), 1666 => to_unsigned(1393, 12), 1667 => to_unsigned(2653, 12), 1668 => to_unsigned(3959, 12), 1669 => to_unsigned(2451, 12), 1670 => to_unsigned(304, 12), 1671 => to_unsigned(265, 12), 1672 => to_unsigned(923, 12), 1673 => to_unsigned(325, 12), 1674 => to_unsigned(3493, 12), 1675 => to_unsigned(1623, 12), 1676 => to_unsigned(574, 12), 1677 => to_unsigned(3582, 12), 1678 => to_unsigned(1779, 12), 1679 => to_unsigned(2584, 12), 1680 => to_unsigned(2105, 12), 1681 => to_unsigned(2570, 12), 1682 => to_unsigned(4088, 12), 1683 => to_unsigned(3658, 12), 1684 => to_unsigned(3464, 12), 1685 => to_unsigned(2819, 12), 1686 => to_unsigned(2768, 12), 1687 => to_unsigned(2076, 12), 1688 => to_unsigned(3637, 12), 1689 => to_unsigned(4076, 12), 1690 => to_unsigned(2155, 12), 1691 => to_unsigned(806, 12), 1692 => to_unsigned(3481, 12), 1693 => to_unsigned(1444, 12), 1694 => to_unsigned(2056, 12), 1695 => to_unsigned(2172, 12), 1696 => to_unsigned(1336, 12), 1697 => to_unsigned(2398, 12), 1698 => to_unsigned(758, 12), 1699 => to_unsigned(1034, 12), 1700 => to_unsigned(2980, 12), 1701 => to_unsigned(341, 12), 1702 => to_unsigned(2855, 12), 1703 => to_unsigned(3484, 12), 1704 => to_unsigned(2413, 12), 1705 => to_unsigned(2865, 12), 1706 => to_unsigned(2147, 12), 1707 => to_unsigned(2209, 12), 1708 => to_unsigned(1648, 12), 1709 => to_unsigned(3067, 12), 1710 => to_unsigned(4011, 12), 1711 => to_unsigned(603, 12), 1712 => to_unsigned(2687, 12), 1713 => to_unsigned(1052, 12), 1714 => to_unsigned(2881, 12), 1715 => to_unsigned(1374, 12), 1716 => to_unsigned(942, 12), 1717 => to_unsigned(1566, 12), 1718 => to_unsigned(240, 12), 1719 => to_unsigned(1998, 12), 1720 => to_unsigned(1729, 12), 1721 => to_unsigned(3571, 12), 1722 => to_unsigned(2976, 12), 1723 => to_unsigned(1518, 12), 1724 => to_unsigned(3594, 12), 1725 => to_unsigned(121, 12), 1726 => to_unsigned(2650, 12), 1727 => to_unsigned(2920, 12), 1728 => to_unsigned(653, 12), 1729 => to_unsigned(138, 12), 1730 => to_unsigned(3772, 12), 1731 => to_unsigned(3005, 12), 1732 => to_unsigned(3477, 12), 1733 => to_unsigned(3504, 12), 1734 => to_unsigned(343, 12), 1735 => to_unsigned(76, 12), 1736 => to_unsigned(3363, 12), 1737 => to_unsigned(365, 12), 1738 => to_unsigned(989, 12), 1739 => to_unsigned(3088, 12), 1740 => to_unsigned(245, 12), 1741 => to_unsigned(107, 12), 1742 => to_unsigned(777, 12), 1743 => to_unsigned(4093, 12), 1744 => to_unsigned(2028, 12), 1745 => to_unsigned(2700, 12), 1746 => to_unsigned(127, 12), 1747 => to_unsigned(782, 12), 1748 => to_unsigned(1580, 12), 1749 => to_unsigned(2445, 12), 1750 => to_unsigned(3420, 12), 1751 => to_unsigned(2954, 12), 1752 => to_unsigned(2458, 12), 1753 => to_unsigned(4060, 12), 1754 => to_unsigned(3902, 12), 1755 => to_unsigned(2304, 12), 1756 => to_unsigned(2162, 12), 1757 => to_unsigned(1243, 12), 1758 => to_unsigned(2931, 12), 1759 => to_unsigned(2759, 12), 1760 => to_unsigned(3245, 12), 1761 => to_unsigned(1843, 12), 1762 => to_unsigned(52, 12), 1763 => to_unsigned(2295, 12), 1764 => to_unsigned(197, 12), 1765 => to_unsigned(2443, 12), 1766 => to_unsigned(2881, 12), 1767 => to_unsigned(306, 12), 1768 => to_unsigned(3412, 12), 1769 => to_unsigned(223, 12), 1770 => to_unsigned(1821, 12), 1771 => to_unsigned(3517, 12), 1772 => to_unsigned(1160, 12), 1773 => to_unsigned(3680, 12), 1774 => to_unsigned(2331, 12), 1775 => to_unsigned(3197, 12), 1776 => to_unsigned(2809, 12), 1777 => to_unsigned(3104, 12), 1778 => to_unsigned(2605, 12), 1779 => to_unsigned(3246, 12), 1780 => to_unsigned(2782, 12), 1781 => to_unsigned(565, 12), 1782 => to_unsigned(2762, 12), 1783 => to_unsigned(2996, 12), 1784 => to_unsigned(347, 12), 1785 => to_unsigned(47, 12), 1786 => to_unsigned(1092, 12), 1787 => to_unsigned(1418, 12), 1788 => to_unsigned(2800, 12), 1789 => to_unsigned(728, 12), 1790 => to_unsigned(3115, 12), 1791 => to_unsigned(2660, 12), 1792 => to_unsigned(384, 12), 1793 => to_unsigned(3253, 12), 1794 => to_unsigned(1561, 12), 1795 => to_unsigned(2180, 12), 1796 => to_unsigned(3462, 12), 1797 => to_unsigned(1050, 12), 1798 => to_unsigned(3589, 12), 1799 => to_unsigned(479, 12), 1800 => to_unsigned(1001, 12), 1801 => to_unsigned(4016, 12), 1802 => to_unsigned(180, 12), 1803 => to_unsigned(3626, 12), 1804 => to_unsigned(442, 12), 1805 => to_unsigned(3984, 12), 1806 => to_unsigned(954, 12), 1807 => to_unsigned(3986, 12), 1808 => to_unsigned(3263, 12), 1809 => to_unsigned(2878, 12), 1810 => to_unsigned(1801, 12), 1811 => to_unsigned(616, 12), 1812 => to_unsigned(1833, 12), 1813 => to_unsigned(3676, 12), 1814 => to_unsigned(1026, 12), 1815 => to_unsigned(1118, 12), 1816 => to_unsigned(3162, 12), 1817 => to_unsigned(1480, 12), 1818 => to_unsigned(1173, 12), 1819 => to_unsigned(3930, 12), 1820 => to_unsigned(795, 12), 1821 => to_unsigned(1703, 12), 1822 => to_unsigned(4012, 12), 1823 => to_unsigned(3449, 12), 1824 => to_unsigned(1406, 12), 1825 => to_unsigned(255, 12), 1826 => to_unsigned(2439, 12), 1827 => to_unsigned(1389, 12), 1828 => to_unsigned(1470, 12), 1829 => to_unsigned(361, 12), 1830 => to_unsigned(3011, 12), 1831 => to_unsigned(2285, 12), 1832 => to_unsigned(2788, 12), 1833 => to_unsigned(35, 12), 1834 => to_unsigned(1048, 12), 1835 => to_unsigned(1937, 12), 1836 => to_unsigned(1449, 12), 1837 => to_unsigned(537, 12), 1838 => to_unsigned(986, 12), 1839 => to_unsigned(2809, 12), 1840 => to_unsigned(995, 12), 1841 => to_unsigned(3542, 12), 1842 => to_unsigned(3344, 12), 1843 => to_unsigned(2827, 12), 1844 => to_unsigned(2263, 12), 1845 => to_unsigned(1204, 12), 1846 => to_unsigned(3072, 12), 1847 => to_unsigned(3762, 12), 1848 => to_unsigned(1110, 12), 1849 => to_unsigned(3149, 12), 1850 => to_unsigned(2864, 12), 1851 => to_unsigned(2818, 12), 1852 => to_unsigned(2467, 12), 1853 => to_unsigned(3393, 12), 1854 => to_unsigned(128, 12), 1855 => to_unsigned(2989, 12), 1856 => to_unsigned(2581, 12), 1857 => to_unsigned(3082, 12), 1858 => to_unsigned(1094, 12), 1859 => to_unsigned(478, 12), 1860 => to_unsigned(1716, 12), 1861 => to_unsigned(228, 12), 1862 => to_unsigned(2167, 12), 1863 => to_unsigned(865, 12), 1864 => to_unsigned(811, 12), 1865 => to_unsigned(1093, 12), 1866 => to_unsigned(847, 12), 1867 => to_unsigned(1186, 12), 1868 => to_unsigned(3056, 12), 1869 => to_unsigned(2953, 12), 1870 => to_unsigned(2796, 12), 1871 => to_unsigned(1898, 12), 1872 => to_unsigned(3228, 12), 1873 => to_unsigned(1771, 12), 1874 => to_unsigned(4078, 12), 1875 => to_unsigned(1449, 12), 1876 => to_unsigned(2661, 12), 1877 => to_unsigned(3926, 12), 1878 => to_unsigned(1795, 12), 1879 => to_unsigned(2178, 12), 1880 => to_unsigned(2392, 12), 1881 => to_unsigned(2118, 12), 1882 => to_unsigned(3845, 12), 1883 => to_unsigned(1335, 12), 1884 => to_unsigned(173, 12), 1885 => to_unsigned(123, 12), 1886 => to_unsigned(2413, 12), 1887 => to_unsigned(2114, 12), 1888 => to_unsigned(1486, 12), 1889 => to_unsigned(1670, 12), 1890 => to_unsigned(3140, 12), 1891 => to_unsigned(3725, 12), 1892 => to_unsigned(914, 12), 1893 => to_unsigned(674, 12), 1894 => to_unsigned(1264, 12), 1895 => to_unsigned(180, 12), 1896 => to_unsigned(171, 12), 1897 => to_unsigned(171, 12), 1898 => to_unsigned(3926, 12), 1899 => to_unsigned(617, 12), 1900 => to_unsigned(2271, 12), 1901 => to_unsigned(3044, 12), 1902 => to_unsigned(1053, 12), 1903 => to_unsigned(3260, 12), 1904 => to_unsigned(3845, 12), 1905 => to_unsigned(480, 12), 1906 => to_unsigned(1563, 12), 1907 => to_unsigned(1574, 12), 1908 => to_unsigned(38, 12), 1909 => to_unsigned(3349, 12), 1910 => to_unsigned(2621, 12), 1911 => to_unsigned(3995, 12), 1912 => to_unsigned(538, 12), 1913 => to_unsigned(1947, 12), 1914 => to_unsigned(796, 12), 1915 => to_unsigned(1653, 12), 1916 => to_unsigned(2838, 12), 1917 => to_unsigned(2668, 12), 1918 => to_unsigned(3033, 12), 1919 => to_unsigned(1915, 12), 1920 => to_unsigned(3041, 12), 1921 => to_unsigned(501, 12), 1922 => to_unsigned(3014, 12), 1923 => to_unsigned(2524, 12), 1924 => to_unsigned(334, 12), 1925 => to_unsigned(370, 12), 1926 => to_unsigned(2056, 12), 1927 => to_unsigned(2599, 12), 1928 => to_unsigned(694, 12), 1929 => to_unsigned(3381, 12), 1930 => to_unsigned(3534, 12), 1931 => to_unsigned(2167, 12), 1932 => to_unsigned(3594, 12), 1933 => to_unsigned(1443, 12), 1934 => to_unsigned(3475, 12), 1935 => to_unsigned(4001, 12), 1936 => to_unsigned(2703, 12), 1937 => to_unsigned(3070, 12), 1938 => to_unsigned(3792, 12), 1939 => to_unsigned(565, 12), 1940 => to_unsigned(3177, 12), 1941 => to_unsigned(3910, 12), 1942 => to_unsigned(3756, 12), 1943 => to_unsigned(272, 12), 1944 => to_unsigned(2193, 12), 1945 => to_unsigned(876, 12), 1946 => to_unsigned(954, 12), 1947 => to_unsigned(605, 12), 1948 => to_unsigned(2456, 12), 1949 => to_unsigned(2207, 12), 1950 => to_unsigned(2275, 12), 1951 => to_unsigned(3556, 12), 1952 => to_unsigned(3312, 12), 1953 => to_unsigned(14, 12), 1954 => to_unsigned(3402, 12), 1955 => to_unsigned(412, 12), 1956 => to_unsigned(263, 12), 1957 => to_unsigned(3000, 12), 1958 => to_unsigned(346, 12), 1959 => to_unsigned(1342, 12), 1960 => to_unsigned(935, 12), 1961 => to_unsigned(1565, 12), 1962 => to_unsigned(908, 12), 1963 => to_unsigned(1380, 12), 1964 => to_unsigned(2252, 12), 1965 => to_unsigned(3940, 12), 1966 => to_unsigned(2793, 12), 1967 => to_unsigned(193, 12), 1968 => to_unsigned(529, 12), 1969 => to_unsigned(3043, 12), 1970 => to_unsigned(2925, 12), 1971 => to_unsigned(801, 12), 1972 => to_unsigned(860, 12), 1973 => to_unsigned(1396, 12), 1974 => to_unsigned(2589, 12), 1975 => to_unsigned(3641, 12), 1976 => to_unsigned(1402, 12), 1977 => to_unsigned(3288, 12), 1978 => to_unsigned(2010, 12), 1979 => to_unsigned(1953, 12), 1980 => to_unsigned(253, 12), 1981 => to_unsigned(3313, 12), 1982 => to_unsigned(1480, 12), 1983 => to_unsigned(937, 12), 1984 => to_unsigned(3384, 12), 1985 => to_unsigned(2645, 12), 1986 => to_unsigned(3218, 12), 1987 => to_unsigned(1079, 12), 1988 => to_unsigned(2888, 12), 1989 => to_unsigned(1843, 12), 1990 => to_unsigned(1937, 12), 1991 => to_unsigned(2579, 12), 1992 => to_unsigned(3778, 12), 1993 => to_unsigned(551, 12), 1994 => to_unsigned(571, 12), 1995 => to_unsigned(19, 12), 1996 => to_unsigned(2981, 12), 1997 => to_unsigned(180, 12), 1998 => to_unsigned(3725, 12), 1999 => to_unsigned(539, 12), 2000 => to_unsigned(3705, 12), 2001 => to_unsigned(254, 12), 2002 => to_unsigned(3920, 12), 2003 => to_unsigned(785, 12), 2004 => to_unsigned(2126, 12), 2005 => to_unsigned(2045, 12), 2006 => to_unsigned(3735, 12), 2007 => to_unsigned(1946, 12), 2008 => to_unsigned(3036, 12), 2009 => to_unsigned(407, 12), 2010 => to_unsigned(3428, 12), 2011 => to_unsigned(2561, 12), 2012 => to_unsigned(4028, 12), 2013 => to_unsigned(1495, 12), 2014 => to_unsigned(1869, 12), 2015 => to_unsigned(2151, 12), 2016 => to_unsigned(4043, 12), 2017 => to_unsigned(14, 12), 2018 => to_unsigned(3585, 12), 2019 => to_unsigned(689, 12), 2020 => to_unsigned(17, 12), 2021 => to_unsigned(3370, 12), 2022 => to_unsigned(1161, 12), 2023 => to_unsigned(2320, 12), 2024 => to_unsigned(1931, 12), 2025 => to_unsigned(331, 12), 2026 => to_unsigned(2726, 12), 2027 => to_unsigned(1670, 12), 2028 => to_unsigned(453, 12), 2029 => to_unsigned(1848, 12), 2030 => to_unsigned(1820, 12), 2031 => to_unsigned(2538, 12), 2032 => to_unsigned(1481, 12), 2033 => to_unsigned(2862, 12), 2034 => to_unsigned(938, 12), 2035 => to_unsigned(2361, 12), 2036 => to_unsigned(1145, 12), 2037 => to_unsigned(167, 12), 2038 => to_unsigned(110, 12), 2039 => to_unsigned(2043, 12), 2040 => to_unsigned(3691, 12), 2041 => to_unsigned(932, 12), 2042 => to_unsigned(2441, 12), 2043 => to_unsigned(3588, 12), 2044 => to_unsigned(3031, 12), 2045 => to_unsigned(3943, 12), 2046 => to_unsigned(2413, 12), 2047 => to_unsigned(2784, 12)),
            3 => (0 => to_unsigned(3317, 12), 1 => to_unsigned(2957, 12), 2 => to_unsigned(2287, 12), 3 => to_unsigned(3360, 12), 4 => to_unsigned(67, 12), 5 => to_unsigned(1521, 12), 6 => to_unsigned(3247, 12), 7 => to_unsigned(2909, 12), 8 => to_unsigned(2001, 12), 9 => to_unsigned(3992, 12), 10 => to_unsigned(72, 12), 11 => to_unsigned(2692, 12), 12 => to_unsigned(263, 12), 13 => to_unsigned(3550, 12), 14 => to_unsigned(2067, 12), 15 => to_unsigned(459, 12), 16 => to_unsigned(3332, 12), 17 => to_unsigned(2755, 12), 18 => to_unsigned(949, 12), 19 => to_unsigned(3689, 12), 20 => to_unsigned(706, 12), 21 => to_unsigned(3081, 12), 22 => to_unsigned(721, 12), 23 => to_unsigned(3740, 12), 24 => to_unsigned(3055, 12), 25 => to_unsigned(3808, 12), 26 => to_unsigned(94, 12), 27 => to_unsigned(1571, 12), 28 => to_unsigned(452, 12), 29 => to_unsigned(2324, 12), 30 => to_unsigned(2557, 12), 31 => to_unsigned(2223, 12), 32 => to_unsigned(996, 12), 33 => to_unsigned(1886, 12), 34 => to_unsigned(234, 12), 35 => to_unsigned(925, 12), 36 => to_unsigned(3620, 12), 37 => to_unsigned(187, 12), 38 => to_unsigned(4004, 12), 39 => to_unsigned(2136, 12), 40 => to_unsigned(1929, 12), 41 => to_unsigned(3278, 12), 42 => to_unsigned(3123, 12), 43 => to_unsigned(1412, 12), 44 => to_unsigned(463, 12), 45 => to_unsigned(3832, 12), 46 => to_unsigned(1161, 12), 47 => to_unsigned(3551, 12), 48 => to_unsigned(2229, 12), 49 => to_unsigned(1775, 12), 50 => to_unsigned(3931, 12), 51 => to_unsigned(2835, 12), 52 => to_unsigned(1317, 12), 53 => to_unsigned(1899, 12), 54 => to_unsigned(1491, 12), 55 => to_unsigned(2065, 12), 56 => to_unsigned(2186, 12), 57 => to_unsigned(1769, 12), 58 => to_unsigned(315, 12), 59 => to_unsigned(398, 12), 60 => to_unsigned(60, 12), 61 => to_unsigned(1840, 12), 62 => to_unsigned(1279, 12), 63 => to_unsigned(27, 12), 64 => to_unsigned(466, 12), 65 => to_unsigned(2309, 12), 66 => to_unsigned(1197, 12), 67 => to_unsigned(1156, 12), 68 => to_unsigned(2984, 12), 69 => to_unsigned(2530, 12), 70 => to_unsigned(3525, 12), 71 => to_unsigned(1417, 12), 72 => to_unsigned(3105, 12), 73 => to_unsigned(3156, 12), 74 => to_unsigned(2344, 12), 75 => to_unsigned(1367, 12), 76 => to_unsigned(427, 12), 77 => to_unsigned(1460, 12), 78 => to_unsigned(3791, 12), 79 => to_unsigned(1543, 12), 80 => to_unsigned(2421, 12), 81 => to_unsigned(2733, 12), 82 => to_unsigned(2214, 12), 83 => to_unsigned(2864, 12), 84 => to_unsigned(920, 12), 85 => to_unsigned(2263, 12), 86 => to_unsigned(3013, 12), 87 => to_unsigned(381, 12), 88 => to_unsigned(1612, 12), 89 => to_unsigned(212, 12), 90 => to_unsigned(1790, 12), 91 => to_unsigned(1804, 12), 92 => to_unsigned(3420, 12), 93 => to_unsigned(547, 12), 94 => to_unsigned(2517, 12), 95 => to_unsigned(1925, 12), 96 => to_unsigned(294, 12), 97 => to_unsigned(1972, 12), 98 => to_unsigned(2129, 12), 99 => to_unsigned(1207, 12), 100 => to_unsigned(252, 12), 101 => to_unsigned(500, 12), 102 => to_unsigned(2369, 12), 103 => to_unsigned(1203, 12), 104 => to_unsigned(3852, 12), 105 => to_unsigned(8, 12), 106 => to_unsigned(2755, 12), 107 => to_unsigned(573, 12), 108 => to_unsigned(3748, 12), 109 => to_unsigned(3213, 12), 110 => to_unsigned(2775, 12), 111 => to_unsigned(2375, 12), 112 => to_unsigned(3495, 12), 113 => to_unsigned(3125, 12), 114 => to_unsigned(606, 12), 115 => to_unsigned(1828, 12), 116 => to_unsigned(2990, 12), 117 => to_unsigned(1992, 12), 118 => to_unsigned(3914, 12), 119 => to_unsigned(1541, 12), 120 => to_unsigned(2087, 12), 121 => to_unsigned(3714, 12), 122 => to_unsigned(275, 12), 123 => to_unsigned(2617, 12), 124 => to_unsigned(1539, 12), 125 => to_unsigned(1530, 12), 126 => to_unsigned(4023, 12), 127 => to_unsigned(600, 12), 128 => to_unsigned(3402, 12), 129 => to_unsigned(2390, 12), 130 => to_unsigned(1537, 12), 131 => to_unsigned(1427, 12), 132 => to_unsigned(2332, 12), 133 => to_unsigned(3451, 12), 134 => to_unsigned(3954, 12), 135 => to_unsigned(3229, 12), 136 => to_unsigned(3937, 12), 137 => to_unsigned(2070, 12), 138 => to_unsigned(1927, 12), 139 => to_unsigned(1160, 12), 140 => to_unsigned(878, 12), 141 => to_unsigned(1648, 12), 142 => to_unsigned(681, 12), 143 => to_unsigned(989, 12), 144 => to_unsigned(2771, 12), 145 => to_unsigned(1046, 12), 146 => to_unsigned(1769, 12), 147 => to_unsigned(1864, 12), 148 => to_unsigned(3761, 12), 149 => to_unsigned(583, 12), 150 => to_unsigned(64, 12), 151 => to_unsigned(3100, 12), 152 => to_unsigned(3269, 12), 153 => to_unsigned(2451, 12), 154 => to_unsigned(2289, 12), 155 => to_unsigned(2311, 12), 156 => to_unsigned(572, 12), 157 => to_unsigned(2747, 12), 158 => to_unsigned(2854, 12), 159 => to_unsigned(360, 12), 160 => to_unsigned(985, 12), 161 => to_unsigned(645, 12), 162 => to_unsigned(1827, 12), 163 => to_unsigned(216, 12), 164 => to_unsigned(2166, 12), 165 => to_unsigned(522, 12), 166 => to_unsigned(3900, 12), 167 => to_unsigned(1131, 12), 168 => to_unsigned(201, 12), 169 => to_unsigned(4004, 12), 170 => to_unsigned(698, 12), 171 => to_unsigned(789, 12), 172 => to_unsigned(272, 12), 173 => to_unsigned(1069, 12), 174 => to_unsigned(1651, 12), 175 => to_unsigned(3044, 12), 176 => to_unsigned(3280, 12), 177 => to_unsigned(3434, 12), 178 => to_unsigned(902, 12), 179 => to_unsigned(437, 12), 180 => to_unsigned(2729, 12), 181 => to_unsigned(1817, 12), 182 => to_unsigned(244, 12), 183 => to_unsigned(1442, 12), 184 => to_unsigned(67, 12), 185 => to_unsigned(3323, 12), 186 => to_unsigned(1686, 12), 187 => to_unsigned(2141, 12), 188 => to_unsigned(3764, 12), 189 => to_unsigned(408, 12), 190 => to_unsigned(1969, 12), 191 => to_unsigned(2849, 12), 192 => to_unsigned(2019, 12), 193 => to_unsigned(3416, 12), 194 => to_unsigned(3366, 12), 195 => to_unsigned(1099, 12), 196 => to_unsigned(702, 12), 197 => to_unsigned(618, 12), 198 => to_unsigned(4003, 12), 199 => to_unsigned(3800, 12), 200 => to_unsigned(3001, 12), 201 => to_unsigned(3825, 12), 202 => to_unsigned(1543, 12), 203 => to_unsigned(2148, 12), 204 => to_unsigned(1675, 12), 205 => to_unsigned(3200, 12), 206 => to_unsigned(420, 12), 207 => to_unsigned(5, 12), 208 => to_unsigned(2057, 12), 209 => to_unsigned(889, 12), 210 => to_unsigned(3653, 12), 211 => to_unsigned(682, 12), 212 => to_unsigned(2318, 12), 213 => to_unsigned(1110, 12), 214 => to_unsigned(1318, 12), 215 => to_unsigned(1313, 12), 216 => to_unsigned(1059, 12), 217 => to_unsigned(3720, 12), 218 => to_unsigned(3551, 12), 219 => to_unsigned(2, 12), 220 => to_unsigned(2999, 12), 221 => to_unsigned(2084, 12), 222 => to_unsigned(1980, 12), 223 => to_unsigned(20, 12), 224 => to_unsigned(2963, 12), 225 => to_unsigned(2157, 12), 226 => to_unsigned(1694, 12), 227 => to_unsigned(329, 12), 228 => to_unsigned(3988, 12), 229 => to_unsigned(3233, 12), 230 => to_unsigned(1895, 12), 231 => to_unsigned(2018, 12), 232 => to_unsigned(4058, 12), 233 => to_unsigned(1618, 12), 234 => to_unsigned(740, 12), 235 => to_unsigned(2226, 12), 236 => to_unsigned(291, 12), 237 => to_unsigned(190, 12), 238 => to_unsigned(2793, 12), 239 => to_unsigned(3786, 12), 240 => to_unsigned(1611, 12), 241 => to_unsigned(581, 12), 242 => to_unsigned(826, 12), 243 => to_unsigned(2808, 12), 244 => to_unsigned(3804, 12), 245 => to_unsigned(356, 12), 246 => to_unsigned(2507, 12), 247 => to_unsigned(2918, 12), 248 => to_unsigned(3510, 12), 249 => to_unsigned(1488, 12), 250 => to_unsigned(675, 12), 251 => to_unsigned(3412, 12), 252 => to_unsigned(3938, 12), 253 => to_unsigned(1868, 12), 254 => to_unsigned(3459, 12), 255 => to_unsigned(2749, 12), 256 => to_unsigned(253, 12), 257 => to_unsigned(2214, 12), 258 => to_unsigned(1001, 12), 259 => to_unsigned(3708, 12), 260 => to_unsigned(3655, 12), 261 => to_unsigned(1519, 12), 262 => to_unsigned(1803, 12), 263 => to_unsigned(1237, 12), 264 => to_unsigned(3957, 12), 265 => to_unsigned(1621, 12), 266 => to_unsigned(3790, 12), 267 => to_unsigned(139, 12), 268 => to_unsigned(1281, 12), 269 => to_unsigned(2700, 12), 270 => to_unsigned(554, 12), 271 => to_unsigned(3863, 12), 272 => to_unsigned(2245, 12), 273 => to_unsigned(1968, 12), 274 => to_unsigned(879, 12), 275 => to_unsigned(3621, 12), 276 => to_unsigned(1164, 12), 277 => to_unsigned(1587, 12), 278 => to_unsigned(1362, 12), 279 => to_unsigned(2584, 12), 280 => to_unsigned(3092, 12), 281 => to_unsigned(1552, 12), 282 => to_unsigned(3087, 12), 283 => to_unsigned(3726, 12), 284 => to_unsigned(869, 12), 285 => to_unsigned(2212, 12), 286 => to_unsigned(2428, 12), 287 => to_unsigned(2391, 12), 288 => to_unsigned(3747, 12), 289 => to_unsigned(3732, 12), 290 => to_unsigned(310, 12), 291 => to_unsigned(2154, 12), 292 => to_unsigned(255, 12), 293 => to_unsigned(3319, 12), 294 => to_unsigned(3978, 12), 295 => to_unsigned(1223, 12), 296 => to_unsigned(1213, 12), 297 => to_unsigned(1140, 12), 298 => to_unsigned(1959, 12), 299 => to_unsigned(3477, 12), 300 => to_unsigned(1473, 12), 301 => to_unsigned(1908, 12), 302 => to_unsigned(2314, 12), 303 => to_unsigned(2653, 12), 304 => to_unsigned(3227, 12), 305 => to_unsigned(436, 12), 306 => to_unsigned(611, 12), 307 => to_unsigned(2413, 12), 308 => to_unsigned(544, 12), 309 => to_unsigned(135, 12), 310 => to_unsigned(1446, 12), 311 => to_unsigned(633, 12), 312 => to_unsigned(1198, 12), 313 => to_unsigned(2614, 12), 314 => to_unsigned(406, 12), 315 => to_unsigned(3304, 12), 316 => to_unsigned(1812, 12), 317 => to_unsigned(68, 12), 318 => to_unsigned(766, 12), 319 => to_unsigned(2006, 12), 320 => to_unsigned(1892, 12), 321 => to_unsigned(1184, 12), 322 => to_unsigned(3648, 12), 323 => to_unsigned(2899, 12), 324 => to_unsigned(3728, 12), 325 => to_unsigned(3371, 12), 326 => to_unsigned(1481, 12), 327 => to_unsigned(3395, 12), 328 => to_unsigned(3152, 12), 329 => to_unsigned(3569, 12), 330 => to_unsigned(2550, 12), 331 => to_unsigned(719, 12), 332 => to_unsigned(721, 12), 333 => to_unsigned(844, 12), 334 => to_unsigned(1570, 12), 335 => to_unsigned(811, 12), 336 => to_unsigned(312, 12), 337 => to_unsigned(2968, 12), 338 => to_unsigned(3904, 12), 339 => to_unsigned(2736, 12), 340 => to_unsigned(1952, 12), 341 => to_unsigned(2440, 12), 342 => to_unsigned(1635, 12), 343 => to_unsigned(2191, 12), 344 => to_unsigned(2032, 12), 345 => to_unsigned(1954, 12), 346 => to_unsigned(1530, 12), 347 => to_unsigned(3557, 12), 348 => to_unsigned(3831, 12), 349 => to_unsigned(792, 12), 350 => to_unsigned(3668, 12), 351 => to_unsigned(1452, 12), 352 => to_unsigned(3671, 12), 353 => to_unsigned(559, 12), 354 => to_unsigned(978, 12), 355 => to_unsigned(3333, 12), 356 => to_unsigned(1268, 12), 357 => to_unsigned(309, 12), 358 => to_unsigned(3138, 12), 359 => to_unsigned(4076, 12), 360 => to_unsigned(1136, 12), 361 => to_unsigned(3764, 12), 362 => to_unsigned(2965, 12), 363 => to_unsigned(2788, 12), 364 => to_unsigned(859, 12), 365 => to_unsigned(843, 12), 366 => to_unsigned(2636, 12), 367 => to_unsigned(2927, 12), 368 => to_unsigned(887, 12), 369 => to_unsigned(633, 12), 370 => to_unsigned(3774, 12), 371 => to_unsigned(1512, 12), 372 => to_unsigned(2222, 12), 373 => to_unsigned(781, 12), 374 => to_unsigned(3610, 12), 375 => to_unsigned(299, 12), 376 => to_unsigned(481, 12), 377 => to_unsigned(3753, 12), 378 => to_unsigned(2188, 12), 379 => to_unsigned(38, 12), 380 => to_unsigned(2066, 12), 381 => to_unsigned(3241, 12), 382 => to_unsigned(3739, 12), 383 => to_unsigned(3461, 12), 384 => to_unsigned(3900, 12), 385 => to_unsigned(2058, 12), 386 => to_unsigned(3295, 12), 387 => to_unsigned(961, 12), 388 => to_unsigned(282, 12), 389 => to_unsigned(2709, 12), 390 => to_unsigned(2199, 12), 391 => to_unsigned(1461, 12), 392 => to_unsigned(85, 12), 393 => to_unsigned(1023, 12), 394 => to_unsigned(2511, 12), 395 => to_unsigned(1072, 12), 396 => to_unsigned(2980, 12), 397 => to_unsigned(2177, 12), 398 => to_unsigned(2871, 12), 399 => to_unsigned(342, 12), 400 => to_unsigned(967, 12), 401 => to_unsigned(2749, 12), 402 => to_unsigned(3758, 12), 403 => to_unsigned(2545, 12), 404 => to_unsigned(585, 12), 405 => to_unsigned(2760, 12), 406 => to_unsigned(2060, 12), 407 => to_unsigned(956, 12), 408 => to_unsigned(1627, 12), 409 => to_unsigned(3331, 12), 410 => to_unsigned(917, 12), 411 => to_unsigned(77, 12), 412 => to_unsigned(2229, 12), 413 => to_unsigned(3494, 12), 414 => to_unsigned(1252, 12), 415 => to_unsigned(570, 12), 416 => to_unsigned(3764, 12), 417 => to_unsigned(739, 12), 418 => to_unsigned(3137, 12), 419 => to_unsigned(107, 12), 420 => to_unsigned(948, 12), 421 => to_unsigned(3408, 12), 422 => to_unsigned(1738, 12), 423 => to_unsigned(2061, 12), 424 => to_unsigned(2568, 12), 425 => to_unsigned(2418, 12), 426 => to_unsigned(2885, 12), 427 => to_unsigned(232, 12), 428 => to_unsigned(2102, 12), 429 => to_unsigned(2515, 12), 430 => to_unsigned(3057, 12), 431 => to_unsigned(751, 12), 432 => to_unsigned(3963, 12), 433 => to_unsigned(3250, 12), 434 => to_unsigned(4002, 12), 435 => to_unsigned(735, 12), 436 => to_unsigned(294, 12), 437 => to_unsigned(3922, 12), 438 => to_unsigned(966, 12), 439 => to_unsigned(1899, 12), 440 => to_unsigned(1678, 12), 441 => to_unsigned(3231, 12), 442 => to_unsigned(758, 12), 443 => to_unsigned(3440, 12), 444 => to_unsigned(2476, 12), 445 => to_unsigned(2208, 12), 446 => to_unsigned(3103, 12), 447 => to_unsigned(593, 12), 448 => to_unsigned(1856, 12), 449 => to_unsigned(2427, 12), 450 => to_unsigned(2708, 12), 451 => to_unsigned(266, 12), 452 => to_unsigned(2386, 12), 453 => to_unsigned(931, 12), 454 => to_unsigned(2271, 12), 455 => to_unsigned(950, 12), 456 => to_unsigned(116, 12), 457 => to_unsigned(2589, 12), 458 => to_unsigned(2784, 12), 459 => to_unsigned(940, 12), 460 => to_unsigned(3214, 12), 461 => to_unsigned(2512, 12), 462 => to_unsigned(2208, 12), 463 => to_unsigned(476, 12), 464 => to_unsigned(950, 12), 465 => to_unsigned(1265, 12), 466 => to_unsigned(3278, 12), 467 => to_unsigned(1959, 12), 468 => to_unsigned(3316, 12), 469 => to_unsigned(691, 12), 470 => to_unsigned(2105, 12), 471 => to_unsigned(920, 12), 472 => to_unsigned(1647, 12), 473 => to_unsigned(2448, 12), 474 => to_unsigned(3829, 12), 475 => to_unsigned(1386, 12), 476 => to_unsigned(2453, 12), 477 => to_unsigned(2029, 12), 478 => to_unsigned(779, 12), 479 => to_unsigned(3109, 12), 480 => to_unsigned(2210, 12), 481 => to_unsigned(3617, 12), 482 => to_unsigned(1302, 12), 483 => to_unsigned(102, 12), 484 => to_unsigned(2576, 12), 485 => to_unsigned(3701, 12), 486 => to_unsigned(3364, 12), 487 => to_unsigned(2752, 12), 488 => to_unsigned(2458, 12), 489 => to_unsigned(77, 12), 490 => to_unsigned(3929, 12), 491 => to_unsigned(3838, 12), 492 => to_unsigned(590, 12), 493 => to_unsigned(1951, 12), 494 => to_unsigned(800, 12), 495 => to_unsigned(2585, 12), 496 => to_unsigned(496, 12), 497 => to_unsigned(3828, 12), 498 => to_unsigned(135, 12), 499 => to_unsigned(1599, 12), 500 => to_unsigned(1484, 12), 501 => to_unsigned(144, 12), 502 => to_unsigned(2344, 12), 503 => to_unsigned(3589, 12), 504 => to_unsigned(1651, 12), 505 => to_unsigned(169, 12), 506 => to_unsigned(1709, 12), 507 => to_unsigned(2517, 12), 508 => to_unsigned(3354, 12), 509 => to_unsigned(329, 12), 510 => to_unsigned(3837, 12), 511 => to_unsigned(3766, 12), 512 => to_unsigned(1864, 12), 513 => to_unsigned(3909, 12), 514 => to_unsigned(2780, 12), 515 => to_unsigned(1554, 12), 516 => to_unsigned(1692, 12), 517 => to_unsigned(2340, 12), 518 => to_unsigned(2603, 12), 519 => to_unsigned(3674, 12), 520 => to_unsigned(3076, 12), 521 => to_unsigned(357, 12), 522 => to_unsigned(2372, 12), 523 => to_unsigned(2759, 12), 524 => to_unsigned(3384, 12), 525 => to_unsigned(4084, 12), 526 => to_unsigned(2754, 12), 527 => to_unsigned(3978, 12), 528 => to_unsigned(2665, 12), 529 => to_unsigned(3303, 12), 530 => to_unsigned(3165, 12), 531 => to_unsigned(3770, 12), 532 => to_unsigned(648, 12), 533 => to_unsigned(3054, 12), 534 => to_unsigned(2841, 12), 535 => to_unsigned(422, 12), 536 => to_unsigned(656, 12), 537 => to_unsigned(3855, 12), 538 => to_unsigned(298, 12), 539 => to_unsigned(1667, 12), 540 => to_unsigned(3510, 12), 541 => to_unsigned(3092, 12), 542 => to_unsigned(2334, 12), 543 => to_unsigned(1370, 12), 544 => to_unsigned(1642, 12), 545 => to_unsigned(2739, 12), 546 => to_unsigned(402, 12), 547 => to_unsigned(199, 12), 548 => to_unsigned(3996, 12), 549 => to_unsigned(1127, 12), 550 => to_unsigned(1268, 12), 551 => to_unsigned(3923, 12), 552 => to_unsigned(1398, 12), 553 => to_unsigned(3614, 12), 554 => to_unsigned(3443, 12), 555 => to_unsigned(2625, 12), 556 => to_unsigned(981, 12), 557 => to_unsigned(866, 12), 558 => to_unsigned(1733, 12), 559 => to_unsigned(196, 12), 560 => to_unsigned(1314, 12), 561 => to_unsigned(1078, 12), 562 => to_unsigned(602, 12), 563 => to_unsigned(2028, 12), 564 => to_unsigned(2537, 12), 565 => to_unsigned(3505, 12), 566 => to_unsigned(3095, 12), 567 => to_unsigned(3943, 12), 568 => to_unsigned(389, 12), 569 => to_unsigned(286, 12), 570 => to_unsigned(2798, 12), 571 => to_unsigned(3736, 12), 572 => to_unsigned(2337, 12), 573 => to_unsigned(3817, 12), 574 => to_unsigned(3228, 12), 575 => to_unsigned(3336, 12), 576 => to_unsigned(1907, 12), 577 => to_unsigned(2235, 12), 578 => to_unsigned(352, 12), 579 => to_unsigned(3438, 12), 580 => to_unsigned(857, 12), 581 => to_unsigned(2696, 12), 582 => to_unsigned(3081, 12), 583 => to_unsigned(3610, 12), 584 => to_unsigned(3782, 12), 585 => to_unsigned(3692, 12), 586 => to_unsigned(1267, 12), 587 => to_unsigned(3190, 12), 588 => to_unsigned(87, 12), 589 => to_unsigned(2218, 12), 590 => to_unsigned(2975, 12), 591 => to_unsigned(3228, 12), 592 => to_unsigned(2511, 12), 593 => to_unsigned(2372, 12), 594 => to_unsigned(863, 12), 595 => to_unsigned(2040, 12), 596 => to_unsigned(2773, 12), 597 => to_unsigned(77, 12), 598 => to_unsigned(1688, 12), 599 => to_unsigned(1982, 12), 600 => to_unsigned(1084, 12), 601 => to_unsigned(2656, 12), 602 => to_unsigned(3032, 12), 603 => to_unsigned(1220, 12), 604 => to_unsigned(3482, 12), 605 => to_unsigned(612, 12), 606 => to_unsigned(3125, 12), 607 => to_unsigned(1785, 12), 608 => to_unsigned(3829, 12), 609 => to_unsigned(1427, 12), 610 => to_unsigned(2882, 12), 611 => to_unsigned(496, 12), 612 => to_unsigned(3669, 12), 613 => to_unsigned(1733, 12), 614 => to_unsigned(1950, 12), 615 => to_unsigned(2948, 12), 616 => to_unsigned(1562, 12), 617 => to_unsigned(1758, 12), 618 => to_unsigned(2959, 12), 619 => to_unsigned(3339, 12), 620 => to_unsigned(2777, 12), 621 => to_unsigned(678, 12), 622 => to_unsigned(437, 12), 623 => to_unsigned(3566, 12), 624 => to_unsigned(362, 12), 625 => to_unsigned(634, 12), 626 => to_unsigned(73, 12), 627 => to_unsigned(1304, 12), 628 => to_unsigned(2905, 12), 629 => to_unsigned(1846, 12), 630 => to_unsigned(195, 12), 631 => to_unsigned(1513, 12), 632 => to_unsigned(3766, 12), 633 => to_unsigned(1370, 12), 634 => to_unsigned(930, 12), 635 => to_unsigned(3863, 12), 636 => to_unsigned(2143, 12), 637 => to_unsigned(3010, 12), 638 => to_unsigned(3016, 12), 639 => to_unsigned(75, 12), 640 => to_unsigned(2797, 12), 641 => to_unsigned(482, 12), 642 => to_unsigned(2787, 12), 643 => to_unsigned(585, 12), 644 => to_unsigned(825, 12), 645 => to_unsigned(1978, 12), 646 => to_unsigned(3277, 12), 647 => to_unsigned(2601, 12), 648 => to_unsigned(4071, 12), 649 => to_unsigned(959, 12), 650 => to_unsigned(491, 12), 651 => to_unsigned(3214, 12), 652 => to_unsigned(2183, 12), 653 => to_unsigned(4047, 12), 654 => to_unsigned(1187, 12), 655 => to_unsigned(1078, 12), 656 => to_unsigned(413, 12), 657 => to_unsigned(2427, 12), 658 => to_unsigned(2349, 12), 659 => to_unsigned(1090, 12), 660 => to_unsigned(824, 12), 661 => to_unsigned(274, 12), 662 => to_unsigned(745, 12), 663 => to_unsigned(2272, 12), 664 => to_unsigned(1227, 12), 665 => to_unsigned(1184, 12), 666 => to_unsigned(2109, 12), 667 => to_unsigned(1332, 12), 668 => to_unsigned(2310, 12), 669 => to_unsigned(626, 12), 670 => to_unsigned(489, 12), 671 => to_unsigned(2697, 12), 672 => to_unsigned(1002, 12), 673 => to_unsigned(486, 12), 674 => to_unsigned(3756, 12), 675 => to_unsigned(2571, 12), 676 => to_unsigned(3556, 12), 677 => to_unsigned(2414, 12), 678 => to_unsigned(2985, 12), 679 => to_unsigned(992, 12), 680 => to_unsigned(725, 12), 681 => to_unsigned(1619, 12), 682 => to_unsigned(3098, 12), 683 => to_unsigned(364, 12), 684 => to_unsigned(3545, 12), 685 => to_unsigned(1265, 12), 686 => to_unsigned(872, 12), 687 => to_unsigned(831, 12), 688 => to_unsigned(2855, 12), 689 => to_unsigned(2985, 12), 690 => to_unsigned(574, 12), 691 => to_unsigned(1312, 12), 692 => to_unsigned(1534, 12), 693 => to_unsigned(2105, 12), 694 => to_unsigned(1029, 12), 695 => to_unsigned(1114, 12), 696 => to_unsigned(1817, 12), 697 => to_unsigned(1184, 12), 698 => to_unsigned(748, 12), 699 => to_unsigned(2257, 12), 700 => to_unsigned(260, 12), 701 => to_unsigned(2629, 12), 702 => to_unsigned(100, 12), 703 => to_unsigned(947, 12), 704 => to_unsigned(2065, 12), 705 => to_unsigned(2098, 12), 706 => to_unsigned(767, 12), 707 => to_unsigned(2035, 12), 708 => to_unsigned(268, 12), 709 => to_unsigned(1036, 12), 710 => to_unsigned(3713, 12), 711 => to_unsigned(3890, 12), 712 => to_unsigned(3813, 12), 713 => to_unsigned(312, 12), 714 => to_unsigned(3442, 12), 715 => to_unsigned(3456, 12), 716 => to_unsigned(2775, 12), 717 => to_unsigned(1798, 12), 718 => to_unsigned(2826, 12), 719 => to_unsigned(3055, 12), 720 => to_unsigned(1225, 12), 721 => to_unsigned(1968, 12), 722 => to_unsigned(3797, 12), 723 => to_unsigned(1784, 12), 724 => to_unsigned(3931, 12), 725 => to_unsigned(1591, 12), 726 => to_unsigned(1910, 12), 727 => to_unsigned(2384, 12), 728 => to_unsigned(1254, 12), 729 => to_unsigned(347, 12), 730 => to_unsigned(1401, 12), 731 => to_unsigned(3453, 12), 732 => to_unsigned(1958, 12), 733 => to_unsigned(974, 12), 734 => to_unsigned(3499, 12), 735 => to_unsigned(556, 12), 736 => to_unsigned(2634, 12), 737 => to_unsigned(3058, 12), 738 => to_unsigned(1909, 12), 739 => to_unsigned(2077, 12), 740 => to_unsigned(3813, 12), 741 => to_unsigned(27, 12), 742 => to_unsigned(1308, 12), 743 => to_unsigned(2006, 12), 744 => to_unsigned(999, 12), 745 => to_unsigned(3924, 12), 746 => to_unsigned(3680, 12), 747 => to_unsigned(3189, 12), 748 => to_unsigned(2764, 12), 749 => to_unsigned(1977, 12), 750 => to_unsigned(2036, 12), 751 => to_unsigned(1437, 12), 752 => to_unsigned(3194, 12), 753 => to_unsigned(3633, 12), 754 => to_unsigned(2627, 12), 755 => to_unsigned(431, 12), 756 => to_unsigned(843, 12), 757 => to_unsigned(1302, 12), 758 => to_unsigned(3401, 12), 759 => to_unsigned(3383, 12), 760 => to_unsigned(2524, 12), 761 => to_unsigned(1004, 12), 762 => to_unsigned(529, 12), 763 => to_unsigned(662, 12), 764 => to_unsigned(198, 12), 765 => to_unsigned(79, 12), 766 => to_unsigned(2919, 12), 767 => to_unsigned(1555, 12), 768 => to_unsigned(90, 12), 769 => to_unsigned(1367, 12), 770 => to_unsigned(3947, 12), 771 => to_unsigned(2875, 12), 772 => to_unsigned(3535, 12), 773 => to_unsigned(2930, 12), 774 => to_unsigned(3412, 12), 775 => to_unsigned(1969, 12), 776 => to_unsigned(1717, 12), 777 => to_unsigned(3501, 12), 778 => to_unsigned(1196, 12), 779 => to_unsigned(3294, 12), 780 => to_unsigned(1707, 12), 781 => to_unsigned(1889, 12), 782 => to_unsigned(1536, 12), 783 => to_unsigned(1743, 12), 784 => to_unsigned(1386, 12), 785 => to_unsigned(2271, 12), 786 => to_unsigned(1372, 12), 787 => to_unsigned(391, 12), 788 => to_unsigned(2269, 12), 789 => to_unsigned(1805, 12), 790 => to_unsigned(3418, 12), 791 => to_unsigned(1766, 12), 792 => to_unsigned(2628, 12), 793 => to_unsigned(1645, 12), 794 => to_unsigned(2787, 12), 795 => to_unsigned(1633, 12), 796 => to_unsigned(2990, 12), 797 => to_unsigned(521, 12), 798 => to_unsigned(2886, 12), 799 => to_unsigned(3749, 12), 800 => to_unsigned(547, 12), 801 => to_unsigned(1806, 12), 802 => to_unsigned(3218, 12), 803 => to_unsigned(820, 12), 804 => to_unsigned(2975, 12), 805 => to_unsigned(2445, 12), 806 => to_unsigned(1908, 12), 807 => to_unsigned(2245, 12), 808 => to_unsigned(3923, 12), 809 => to_unsigned(2989, 12), 810 => to_unsigned(1196, 12), 811 => to_unsigned(589, 12), 812 => to_unsigned(830, 12), 813 => to_unsigned(1780, 12), 814 => to_unsigned(3313, 12), 815 => to_unsigned(693, 12), 816 => to_unsigned(3483, 12), 817 => to_unsigned(1304, 12), 818 => to_unsigned(673, 12), 819 => to_unsigned(1668, 12), 820 => to_unsigned(950, 12), 821 => to_unsigned(1273, 12), 822 => to_unsigned(300, 12), 823 => to_unsigned(76, 12), 824 => to_unsigned(1819, 12), 825 => to_unsigned(333, 12), 826 => to_unsigned(590, 12), 827 => to_unsigned(65, 12), 828 => to_unsigned(3014, 12), 829 => to_unsigned(1559, 12), 830 => to_unsigned(3334, 12), 831 => to_unsigned(2276, 12), 832 => to_unsigned(2746, 12), 833 => to_unsigned(2755, 12), 834 => to_unsigned(259, 12), 835 => to_unsigned(1331, 12), 836 => to_unsigned(3715, 12), 837 => to_unsigned(1852, 12), 838 => to_unsigned(2918, 12), 839 => to_unsigned(748, 12), 840 => to_unsigned(2372, 12), 841 => to_unsigned(3899, 12), 842 => to_unsigned(286, 12), 843 => to_unsigned(778, 12), 844 => to_unsigned(2374, 12), 845 => to_unsigned(1510, 12), 846 => to_unsigned(1183, 12), 847 => to_unsigned(1199, 12), 848 => to_unsigned(2168, 12), 849 => to_unsigned(2784, 12), 850 => to_unsigned(4008, 12), 851 => to_unsigned(2111, 12), 852 => to_unsigned(1944, 12), 853 => to_unsigned(1461, 12), 854 => to_unsigned(25, 12), 855 => to_unsigned(2906, 12), 856 => to_unsigned(1501, 12), 857 => to_unsigned(2806, 12), 858 => to_unsigned(3909, 12), 859 => to_unsigned(1484, 12), 860 => to_unsigned(1027, 12), 861 => to_unsigned(3155, 12), 862 => to_unsigned(1252, 12), 863 => to_unsigned(1, 12), 864 => to_unsigned(1669, 12), 865 => to_unsigned(2091, 12), 866 => to_unsigned(107, 12), 867 => to_unsigned(3855, 12), 868 => to_unsigned(140, 12), 869 => to_unsigned(2359, 12), 870 => to_unsigned(3323, 12), 871 => to_unsigned(1657, 12), 872 => to_unsigned(437, 12), 873 => to_unsigned(427, 12), 874 => to_unsigned(1160, 12), 875 => to_unsigned(486, 12), 876 => to_unsigned(3253, 12), 877 => to_unsigned(607, 12), 878 => to_unsigned(3014, 12), 879 => to_unsigned(2729, 12), 880 => to_unsigned(1656, 12), 881 => to_unsigned(2055, 12), 882 => to_unsigned(1072, 12), 883 => to_unsigned(2485, 12), 884 => to_unsigned(871, 12), 885 => to_unsigned(3277, 12), 886 => to_unsigned(3336, 12), 887 => to_unsigned(2221, 12), 888 => to_unsigned(1877, 12), 889 => to_unsigned(3590, 12), 890 => to_unsigned(3579, 12), 891 => to_unsigned(3979, 12), 892 => to_unsigned(3785, 12), 893 => to_unsigned(2209, 12), 894 => to_unsigned(652, 12), 895 => to_unsigned(3571, 12), 896 => to_unsigned(2799, 12), 897 => to_unsigned(498, 12), 898 => to_unsigned(1919, 12), 899 => to_unsigned(1956, 12), 900 => to_unsigned(3330, 12), 901 => to_unsigned(3547, 12), 902 => to_unsigned(3355, 12), 903 => to_unsigned(375, 12), 904 => to_unsigned(3172, 12), 905 => to_unsigned(1912, 12), 906 => to_unsigned(1466, 12), 907 => to_unsigned(1807, 12), 908 => to_unsigned(3113, 12), 909 => to_unsigned(1830, 12), 910 => to_unsigned(296, 12), 911 => to_unsigned(3733, 12), 912 => to_unsigned(3314, 12), 913 => to_unsigned(3313, 12), 914 => to_unsigned(2527, 12), 915 => to_unsigned(2184, 12), 916 => to_unsigned(684, 12), 917 => to_unsigned(994, 12), 918 => to_unsigned(2248, 12), 919 => to_unsigned(2882, 12), 920 => to_unsigned(1168, 12), 921 => to_unsigned(2216, 12), 922 => to_unsigned(1419, 12), 923 => to_unsigned(4042, 12), 924 => to_unsigned(396, 12), 925 => to_unsigned(1042, 12), 926 => to_unsigned(629, 12), 927 => to_unsigned(2163, 12), 928 => to_unsigned(1561, 12), 929 => to_unsigned(2116, 12), 930 => to_unsigned(2996, 12), 931 => to_unsigned(1921, 12), 932 => to_unsigned(1157, 12), 933 => to_unsigned(834, 12), 934 => to_unsigned(3842, 12), 935 => to_unsigned(1068, 12), 936 => to_unsigned(373, 12), 937 => to_unsigned(2539, 12), 938 => to_unsigned(39, 12), 939 => to_unsigned(3121, 12), 940 => to_unsigned(1938, 12), 941 => to_unsigned(2384, 12), 942 => to_unsigned(2065, 12), 943 => to_unsigned(879, 12), 944 => to_unsigned(1461, 12), 945 => to_unsigned(3924, 12), 946 => to_unsigned(3052, 12), 947 => to_unsigned(1230, 12), 948 => to_unsigned(3924, 12), 949 => to_unsigned(289, 12), 950 => to_unsigned(969, 12), 951 => to_unsigned(3720, 12), 952 => to_unsigned(2289, 12), 953 => to_unsigned(2776, 12), 954 => to_unsigned(3225, 12), 955 => to_unsigned(418, 12), 956 => to_unsigned(3551, 12), 957 => to_unsigned(3683, 12), 958 => to_unsigned(3090, 12), 959 => to_unsigned(3323, 12), 960 => to_unsigned(4094, 12), 961 => to_unsigned(3717, 12), 962 => to_unsigned(3756, 12), 963 => to_unsigned(2455, 12), 964 => to_unsigned(2744, 12), 965 => to_unsigned(417, 12), 966 => to_unsigned(1520, 12), 967 => to_unsigned(3934, 12), 968 => to_unsigned(1186, 12), 969 => to_unsigned(541, 12), 970 => to_unsigned(2942, 12), 971 => to_unsigned(3852, 12), 972 => to_unsigned(3370, 12), 973 => to_unsigned(3655, 12), 974 => to_unsigned(2547, 12), 975 => to_unsigned(836, 12), 976 => to_unsigned(3307, 12), 977 => to_unsigned(2987, 12), 978 => to_unsigned(3648, 12), 979 => to_unsigned(1088, 12), 980 => to_unsigned(2854, 12), 981 => to_unsigned(2225, 12), 982 => to_unsigned(713, 12), 983 => to_unsigned(2260, 12), 984 => to_unsigned(2632, 12), 985 => to_unsigned(3632, 12), 986 => to_unsigned(2630, 12), 987 => to_unsigned(1908, 12), 988 => to_unsigned(1847, 12), 989 => to_unsigned(788, 12), 990 => to_unsigned(2412, 12), 991 => to_unsigned(3001, 12), 992 => to_unsigned(3073, 12), 993 => to_unsigned(1385, 12), 994 => to_unsigned(1796, 12), 995 => to_unsigned(348, 12), 996 => to_unsigned(3137, 12), 997 => to_unsigned(3411, 12), 998 => to_unsigned(3246, 12), 999 => to_unsigned(2782, 12), 1000 => to_unsigned(1346, 12), 1001 => to_unsigned(2448, 12), 1002 => to_unsigned(2607, 12), 1003 => to_unsigned(1742, 12), 1004 => to_unsigned(2518, 12), 1005 => to_unsigned(248, 12), 1006 => to_unsigned(3344, 12), 1007 => to_unsigned(587, 12), 1008 => to_unsigned(1998, 12), 1009 => to_unsigned(1428, 12), 1010 => to_unsigned(3999, 12), 1011 => to_unsigned(2250, 12), 1012 => to_unsigned(3432, 12), 1013 => to_unsigned(633, 12), 1014 => to_unsigned(2190, 12), 1015 => to_unsigned(166, 12), 1016 => to_unsigned(2699, 12), 1017 => to_unsigned(3085, 12), 1018 => to_unsigned(1582, 12), 1019 => to_unsigned(2555, 12), 1020 => to_unsigned(3328, 12), 1021 => to_unsigned(936, 12), 1022 => to_unsigned(3079, 12), 1023 => to_unsigned(396, 12), 1024 => to_unsigned(1148, 12), 1025 => to_unsigned(769, 12), 1026 => to_unsigned(3218, 12), 1027 => to_unsigned(44, 12), 1028 => to_unsigned(1347, 12), 1029 => to_unsigned(2478, 12), 1030 => to_unsigned(2370, 12), 1031 => to_unsigned(918, 12), 1032 => to_unsigned(636, 12), 1033 => to_unsigned(1525, 12), 1034 => to_unsigned(1946, 12), 1035 => to_unsigned(445, 12), 1036 => to_unsigned(3346, 12), 1037 => to_unsigned(2210, 12), 1038 => to_unsigned(2505, 12), 1039 => to_unsigned(1018, 12), 1040 => to_unsigned(2611, 12), 1041 => to_unsigned(2539, 12), 1042 => to_unsigned(323, 12), 1043 => to_unsigned(3020, 12), 1044 => to_unsigned(809, 12), 1045 => to_unsigned(1830, 12), 1046 => to_unsigned(2928, 12), 1047 => to_unsigned(1007, 12), 1048 => to_unsigned(2333, 12), 1049 => to_unsigned(981, 12), 1050 => to_unsigned(1601, 12), 1051 => to_unsigned(3546, 12), 1052 => to_unsigned(2100, 12), 1053 => to_unsigned(3103, 12), 1054 => to_unsigned(2203, 12), 1055 => to_unsigned(895, 12), 1056 => to_unsigned(520, 12), 1057 => to_unsigned(2705, 12), 1058 => to_unsigned(280, 12), 1059 => to_unsigned(1542, 12), 1060 => to_unsigned(2670, 12), 1061 => to_unsigned(6, 12), 1062 => to_unsigned(3162, 12), 1063 => to_unsigned(2187, 12), 1064 => to_unsigned(444, 12), 1065 => to_unsigned(3671, 12), 1066 => to_unsigned(495, 12), 1067 => to_unsigned(1228, 12), 1068 => to_unsigned(3167, 12), 1069 => to_unsigned(3807, 12), 1070 => to_unsigned(2384, 12), 1071 => to_unsigned(999, 12), 1072 => to_unsigned(2077, 12), 1073 => to_unsigned(2031, 12), 1074 => to_unsigned(727, 12), 1075 => to_unsigned(3181, 12), 1076 => to_unsigned(1316, 12), 1077 => to_unsigned(240, 12), 1078 => to_unsigned(3929, 12), 1079 => to_unsigned(1497, 12), 1080 => to_unsigned(2405, 12), 1081 => to_unsigned(1425, 12), 1082 => to_unsigned(1938, 12), 1083 => to_unsigned(685, 12), 1084 => to_unsigned(1142, 12), 1085 => to_unsigned(1430, 12), 1086 => to_unsigned(2363, 12), 1087 => to_unsigned(3074, 12), 1088 => to_unsigned(3941, 12), 1089 => to_unsigned(3246, 12), 1090 => to_unsigned(3802, 12), 1091 => to_unsigned(1545, 12), 1092 => to_unsigned(2728, 12), 1093 => to_unsigned(434, 12), 1094 => to_unsigned(1473, 12), 1095 => to_unsigned(1179, 12), 1096 => to_unsigned(3555, 12), 1097 => to_unsigned(2476, 12), 1098 => to_unsigned(3306, 12), 1099 => to_unsigned(1965, 12), 1100 => to_unsigned(2380, 12), 1101 => to_unsigned(1798, 12), 1102 => to_unsigned(111, 12), 1103 => to_unsigned(3280, 12), 1104 => to_unsigned(83, 12), 1105 => to_unsigned(1076, 12), 1106 => to_unsigned(3624, 12), 1107 => to_unsigned(3247, 12), 1108 => to_unsigned(881, 12), 1109 => to_unsigned(671, 12), 1110 => to_unsigned(1215, 12), 1111 => to_unsigned(3522, 12), 1112 => to_unsigned(4088, 12), 1113 => to_unsigned(3662, 12), 1114 => to_unsigned(1804, 12), 1115 => to_unsigned(3656, 12), 1116 => to_unsigned(2328, 12), 1117 => to_unsigned(115, 12), 1118 => to_unsigned(1037, 12), 1119 => to_unsigned(2185, 12), 1120 => to_unsigned(3686, 12), 1121 => to_unsigned(3538, 12), 1122 => to_unsigned(1609, 12), 1123 => to_unsigned(1961, 12), 1124 => to_unsigned(2414, 12), 1125 => to_unsigned(1379, 12), 1126 => to_unsigned(2882, 12), 1127 => to_unsigned(3385, 12), 1128 => to_unsigned(2600, 12), 1129 => to_unsigned(2647, 12), 1130 => to_unsigned(3766, 12), 1131 => to_unsigned(1380, 12), 1132 => to_unsigned(716, 12), 1133 => to_unsigned(2146, 12), 1134 => to_unsigned(3548, 12), 1135 => to_unsigned(3440, 12), 1136 => to_unsigned(269, 12), 1137 => to_unsigned(292, 12), 1138 => to_unsigned(2027, 12), 1139 => to_unsigned(1610, 12), 1140 => to_unsigned(3919, 12), 1141 => to_unsigned(298, 12), 1142 => to_unsigned(1508, 12), 1143 => to_unsigned(3494, 12), 1144 => to_unsigned(1886, 12), 1145 => to_unsigned(3499, 12), 1146 => to_unsigned(1813, 12), 1147 => to_unsigned(835, 12), 1148 => to_unsigned(2764, 12), 1149 => to_unsigned(1554, 12), 1150 => to_unsigned(3217, 12), 1151 => to_unsigned(3678, 12), 1152 => to_unsigned(2746, 12), 1153 => to_unsigned(3750, 12), 1154 => to_unsigned(3412, 12), 1155 => to_unsigned(3793, 12), 1156 => to_unsigned(45, 12), 1157 => to_unsigned(4017, 12), 1158 => to_unsigned(288, 12), 1159 => to_unsigned(370, 12), 1160 => to_unsigned(2877, 12), 1161 => to_unsigned(260, 12), 1162 => to_unsigned(291, 12), 1163 => to_unsigned(2774, 12), 1164 => to_unsigned(3251, 12), 1165 => to_unsigned(2691, 12), 1166 => to_unsigned(4007, 12), 1167 => to_unsigned(180, 12), 1168 => to_unsigned(3739, 12), 1169 => to_unsigned(3733, 12), 1170 => to_unsigned(2791, 12), 1171 => to_unsigned(58, 12), 1172 => to_unsigned(2581, 12), 1173 => to_unsigned(3602, 12), 1174 => to_unsigned(1815, 12), 1175 => to_unsigned(1522, 12), 1176 => to_unsigned(719, 12), 1177 => to_unsigned(383, 12), 1178 => to_unsigned(2713, 12), 1179 => to_unsigned(310, 12), 1180 => to_unsigned(2766, 12), 1181 => to_unsigned(32, 12), 1182 => to_unsigned(1304, 12), 1183 => to_unsigned(2556, 12), 1184 => to_unsigned(1028, 12), 1185 => to_unsigned(2174, 12), 1186 => to_unsigned(1872, 12), 1187 => to_unsigned(1385, 12), 1188 => to_unsigned(1251, 12), 1189 => to_unsigned(4050, 12), 1190 => to_unsigned(3844, 12), 1191 => to_unsigned(2551, 12), 1192 => to_unsigned(727, 12), 1193 => to_unsigned(502, 12), 1194 => to_unsigned(2034, 12), 1195 => to_unsigned(3161, 12), 1196 => to_unsigned(2088, 12), 1197 => to_unsigned(2780, 12), 1198 => to_unsigned(3405, 12), 1199 => to_unsigned(1935, 12), 1200 => to_unsigned(1074, 12), 1201 => to_unsigned(712, 12), 1202 => to_unsigned(4019, 12), 1203 => to_unsigned(1979, 12), 1204 => to_unsigned(2140, 12), 1205 => to_unsigned(2627, 12), 1206 => to_unsigned(1536, 12), 1207 => to_unsigned(2833, 12), 1208 => to_unsigned(2797, 12), 1209 => to_unsigned(879, 12), 1210 => to_unsigned(1869, 12), 1211 => to_unsigned(1673, 12), 1212 => to_unsigned(3724, 12), 1213 => to_unsigned(2440, 12), 1214 => to_unsigned(3578, 12), 1215 => to_unsigned(2622, 12), 1216 => to_unsigned(1491, 12), 1217 => to_unsigned(2628, 12), 1218 => to_unsigned(3309, 12), 1219 => to_unsigned(1291, 12), 1220 => to_unsigned(1565, 12), 1221 => to_unsigned(3871, 12), 1222 => to_unsigned(25, 12), 1223 => to_unsigned(616, 12), 1224 => to_unsigned(3488, 12), 1225 => to_unsigned(1642, 12), 1226 => to_unsigned(3421, 12), 1227 => to_unsigned(2808, 12), 1228 => to_unsigned(389, 12), 1229 => to_unsigned(1280, 12), 1230 => to_unsigned(3725, 12), 1231 => to_unsigned(2807, 12), 1232 => to_unsigned(1866, 12), 1233 => to_unsigned(1499, 12), 1234 => to_unsigned(3100, 12), 1235 => to_unsigned(2500, 12), 1236 => to_unsigned(1199, 12), 1237 => to_unsigned(2482, 12), 1238 => to_unsigned(1141, 12), 1239 => to_unsigned(2469, 12), 1240 => to_unsigned(1567, 12), 1241 => to_unsigned(2528, 12), 1242 => to_unsigned(273, 12), 1243 => to_unsigned(1784, 12), 1244 => to_unsigned(1577, 12), 1245 => to_unsigned(4018, 12), 1246 => to_unsigned(3704, 12), 1247 => to_unsigned(2675, 12), 1248 => to_unsigned(304, 12), 1249 => to_unsigned(2432, 12), 1250 => to_unsigned(1734, 12), 1251 => to_unsigned(383, 12), 1252 => to_unsigned(1641, 12), 1253 => to_unsigned(858, 12), 1254 => to_unsigned(460, 12), 1255 => to_unsigned(2682, 12), 1256 => to_unsigned(43, 12), 1257 => to_unsigned(537, 12), 1258 => to_unsigned(854, 12), 1259 => to_unsigned(684, 12), 1260 => to_unsigned(2914, 12), 1261 => to_unsigned(3873, 12), 1262 => to_unsigned(3489, 12), 1263 => to_unsigned(1100, 12), 1264 => to_unsigned(86, 12), 1265 => to_unsigned(3874, 12), 1266 => to_unsigned(2940, 12), 1267 => to_unsigned(1109, 12), 1268 => to_unsigned(1290, 12), 1269 => to_unsigned(3650, 12), 1270 => to_unsigned(1212, 12), 1271 => to_unsigned(3658, 12), 1272 => to_unsigned(3873, 12), 1273 => to_unsigned(3870, 12), 1274 => to_unsigned(496, 12), 1275 => to_unsigned(2375, 12), 1276 => to_unsigned(3951, 12), 1277 => to_unsigned(3740, 12), 1278 => to_unsigned(3295, 12), 1279 => to_unsigned(3196, 12), 1280 => to_unsigned(3338, 12), 1281 => to_unsigned(1670, 12), 1282 => to_unsigned(1848, 12), 1283 => to_unsigned(3299, 12), 1284 => to_unsigned(3671, 12), 1285 => to_unsigned(131, 12), 1286 => to_unsigned(3953, 12), 1287 => to_unsigned(3852, 12), 1288 => to_unsigned(2396, 12), 1289 => to_unsigned(1155, 12), 1290 => to_unsigned(3624, 12), 1291 => to_unsigned(2428, 12), 1292 => to_unsigned(983, 12), 1293 => to_unsigned(643, 12), 1294 => to_unsigned(2902, 12), 1295 => to_unsigned(928, 12), 1296 => to_unsigned(3735, 12), 1297 => to_unsigned(2082, 12), 1298 => to_unsigned(1261, 12), 1299 => to_unsigned(1277, 12), 1300 => to_unsigned(3961, 12), 1301 => to_unsigned(916, 12), 1302 => to_unsigned(704, 12), 1303 => to_unsigned(3955, 12), 1304 => to_unsigned(1255, 12), 1305 => to_unsigned(2335, 12), 1306 => to_unsigned(3431, 12), 1307 => to_unsigned(1808, 12), 1308 => to_unsigned(572, 12), 1309 => to_unsigned(214, 12), 1310 => to_unsigned(3292, 12), 1311 => to_unsigned(3691, 12), 1312 => to_unsigned(814, 12), 1313 => to_unsigned(1778, 12), 1314 => to_unsigned(3198, 12), 1315 => to_unsigned(987, 12), 1316 => to_unsigned(3145, 12), 1317 => to_unsigned(1708, 12), 1318 => to_unsigned(2271, 12), 1319 => to_unsigned(3125, 12), 1320 => to_unsigned(2319, 12), 1321 => to_unsigned(1829, 12), 1322 => to_unsigned(1526, 12), 1323 => to_unsigned(1857, 12), 1324 => to_unsigned(2276, 12), 1325 => to_unsigned(1423, 12), 1326 => to_unsigned(1652, 12), 1327 => to_unsigned(2558, 12), 1328 => to_unsigned(407, 12), 1329 => to_unsigned(965, 12), 1330 => to_unsigned(1811, 12), 1331 => to_unsigned(3551, 12), 1332 => to_unsigned(2689, 12), 1333 => to_unsigned(3771, 12), 1334 => to_unsigned(3092, 12), 1335 => to_unsigned(1995, 12), 1336 => to_unsigned(2029, 12), 1337 => to_unsigned(390, 12), 1338 => to_unsigned(3383, 12), 1339 => to_unsigned(904, 12), 1340 => to_unsigned(2562, 12), 1341 => to_unsigned(4026, 12), 1342 => to_unsigned(162, 12), 1343 => to_unsigned(2670, 12), 1344 => to_unsigned(367, 12), 1345 => to_unsigned(1167, 12), 1346 => to_unsigned(1866, 12), 1347 => to_unsigned(1456, 12), 1348 => to_unsigned(2414, 12), 1349 => to_unsigned(3434, 12), 1350 => to_unsigned(1912, 12), 1351 => to_unsigned(591, 12), 1352 => to_unsigned(4009, 12), 1353 => to_unsigned(1908, 12), 1354 => to_unsigned(1850, 12), 1355 => to_unsigned(3494, 12), 1356 => to_unsigned(2898, 12), 1357 => to_unsigned(4038, 12), 1358 => to_unsigned(289, 12), 1359 => to_unsigned(1631, 12), 1360 => to_unsigned(184, 12), 1361 => to_unsigned(331, 12), 1362 => to_unsigned(2929, 12), 1363 => to_unsigned(1051, 12), 1364 => to_unsigned(2327, 12), 1365 => to_unsigned(458, 12), 1366 => to_unsigned(555, 12), 1367 => to_unsigned(2034, 12), 1368 => to_unsigned(3444, 12), 1369 => to_unsigned(3188, 12), 1370 => to_unsigned(822, 12), 1371 => to_unsigned(3880, 12), 1372 => to_unsigned(2229, 12), 1373 => to_unsigned(1477, 12), 1374 => to_unsigned(46, 12), 1375 => to_unsigned(3452, 12), 1376 => to_unsigned(1154, 12), 1377 => to_unsigned(3872, 12), 1378 => to_unsigned(1645, 12), 1379 => to_unsigned(3920, 12), 1380 => to_unsigned(729, 12), 1381 => to_unsigned(3771, 12), 1382 => to_unsigned(3646, 12), 1383 => to_unsigned(1932, 12), 1384 => to_unsigned(338, 12), 1385 => to_unsigned(3094, 12), 1386 => to_unsigned(431, 12), 1387 => to_unsigned(1674, 12), 1388 => to_unsigned(1584, 12), 1389 => to_unsigned(2334, 12), 1390 => to_unsigned(3139, 12), 1391 => to_unsigned(3208, 12), 1392 => to_unsigned(1199, 12), 1393 => to_unsigned(925, 12), 1394 => to_unsigned(4092, 12), 1395 => to_unsigned(1458, 12), 1396 => to_unsigned(1997, 12), 1397 => to_unsigned(3993, 12), 1398 => to_unsigned(3354, 12), 1399 => to_unsigned(2093, 12), 1400 => to_unsigned(2904, 12), 1401 => to_unsigned(844, 12), 1402 => to_unsigned(203, 12), 1403 => to_unsigned(3640, 12), 1404 => to_unsigned(1315, 12), 1405 => to_unsigned(2470, 12), 1406 => to_unsigned(66, 12), 1407 => to_unsigned(2984, 12), 1408 => to_unsigned(1353, 12), 1409 => to_unsigned(3884, 12), 1410 => to_unsigned(2504, 12), 1411 => to_unsigned(650, 12), 1412 => to_unsigned(2577, 12), 1413 => to_unsigned(3497, 12), 1414 => to_unsigned(2193, 12), 1415 => to_unsigned(2576, 12), 1416 => to_unsigned(3232, 12), 1417 => to_unsigned(101, 12), 1418 => to_unsigned(3205, 12), 1419 => to_unsigned(1097, 12), 1420 => to_unsigned(1669, 12), 1421 => to_unsigned(2319, 12), 1422 => to_unsigned(2325, 12), 1423 => to_unsigned(2978, 12), 1424 => to_unsigned(3750, 12), 1425 => to_unsigned(1662, 12), 1426 => to_unsigned(2976, 12), 1427 => to_unsigned(790, 12), 1428 => to_unsigned(2185, 12), 1429 => to_unsigned(1807, 12), 1430 => to_unsigned(2448, 12), 1431 => to_unsigned(1434, 12), 1432 => to_unsigned(2923, 12), 1433 => to_unsigned(659, 12), 1434 => to_unsigned(2560, 12), 1435 => to_unsigned(2925, 12), 1436 => to_unsigned(2205, 12), 1437 => to_unsigned(1023, 12), 1438 => to_unsigned(1794, 12), 1439 => to_unsigned(2748, 12), 1440 => to_unsigned(3666, 12), 1441 => to_unsigned(3241, 12), 1442 => to_unsigned(2837, 12), 1443 => to_unsigned(1639, 12), 1444 => to_unsigned(2482, 12), 1445 => to_unsigned(2709, 12), 1446 => to_unsigned(1221, 12), 1447 => to_unsigned(626, 12), 1448 => to_unsigned(320, 12), 1449 => to_unsigned(583, 12), 1450 => to_unsigned(1249, 12), 1451 => to_unsigned(3913, 12), 1452 => to_unsigned(2899, 12), 1453 => to_unsigned(3250, 12), 1454 => to_unsigned(1404, 12), 1455 => to_unsigned(2951, 12), 1456 => to_unsigned(952, 12), 1457 => to_unsigned(4079, 12), 1458 => to_unsigned(662, 12), 1459 => to_unsigned(328, 12), 1460 => to_unsigned(3136, 12), 1461 => to_unsigned(730, 12), 1462 => to_unsigned(2965, 12), 1463 => to_unsigned(1072, 12), 1464 => to_unsigned(2786, 12), 1465 => to_unsigned(588, 12), 1466 => to_unsigned(4041, 12), 1467 => to_unsigned(3219, 12), 1468 => to_unsigned(3479, 12), 1469 => to_unsigned(1586, 12), 1470 => to_unsigned(2932, 12), 1471 => to_unsigned(353, 12), 1472 => to_unsigned(2668, 12), 1473 => to_unsigned(2910, 12), 1474 => to_unsigned(140, 12), 1475 => to_unsigned(3363, 12), 1476 => to_unsigned(1487, 12), 1477 => to_unsigned(1327, 12), 1478 => to_unsigned(1440, 12), 1479 => to_unsigned(2787, 12), 1480 => to_unsigned(467, 12), 1481 => to_unsigned(878, 12), 1482 => to_unsigned(669, 12), 1483 => to_unsigned(745, 12), 1484 => to_unsigned(3229, 12), 1485 => to_unsigned(3108, 12), 1486 => to_unsigned(3370, 12), 1487 => to_unsigned(4024, 12), 1488 => to_unsigned(3508, 12), 1489 => to_unsigned(2589, 12), 1490 => to_unsigned(4018, 12), 1491 => to_unsigned(2630, 12), 1492 => to_unsigned(1364, 12), 1493 => to_unsigned(338, 12), 1494 => to_unsigned(3395, 12), 1495 => to_unsigned(3797, 12), 1496 => to_unsigned(73, 12), 1497 => to_unsigned(4090, 12), 1498 => to_unsigned(3147, 12), 1499 => to_unsigned(2235, 12), 1500 => to_unsigned(2410, 12), 1501 => to_unsigned(1245, 12), 1502 => to_unsigned(3340, 12), 1503 => to_unsigned(1143, 12), 1504 => to_unsigned(1001, 12), 1505 => to_unsigned(2768, 12), 1506 => to_unsigned(225, 12), 1507 => to_unsigned(1079, 12), 1508 => to_unsigned(3839, 12), 1509 => to_unsigned(1065, 12), 1510 => to_unsigned(1330, 12), 1511 => to_unsigned(2423, 12), 1512 => to_unsigned(3573, 12), 1513 => to_unsigned(1178, 12), 1514 => to_unsigned(3418, 12), 1515 => to_unsigned(3465, 12), 1516 => to_unsigned(2435, 12), 1517 => to_unsigned(1936, 12), 1518 => to_unsigned(2497, 12), 1519 => to_unsigned(621, 12), 1520 => to_unsigned(3753, 12), 1521 => to_unsigned(3232, 12), 1522 => to_unsigned(1977, 12), 1523 => to_unsigned(1224, 12), 1524 => to_unsigned(2988, 12), 1525 => to_unsigned(627, 12), 1526 => to_unsigned(598, 12), 1527 => to_unsigned(765, 12), 1528 => to_unsigned(3768, 12), 1529 => to_unsigned(1387, 12), 1530 => to_unsigned(3035, 12), 1531 => to_unsigned(2309, 12), 1532 => to_unsigned(669, 12), 1533 => to_unsigned(3574, 12), 1534 => to_unsigned(2154, 12), 1535 => to_unsigned(3928, 12), 1536 => to_unsigned(3729, 12), 1537 => to_unsigned(3875, 12), 1538 => to_unsigned(1835, 12), 1539 => to_unsigned(1459, 12), 1540 => to_unsigned(3915, 12), 1541 => to_unsigned(989, 12), 1542 => to_unsigned(703, 12), 1543 => to_unsigned(2744, 12), 1544 => to_unsigned(1255, 12), 1545 => to_unsigned(2451, 12), 1546 => to_unsigned(2398, 12), 1547 => to_unsigned(660, 12), 1548 => to_unsigned(2215, 12), 1549 => to_unsigned(1936, 12), 1550 => to_unsigned(4042, 12), 1551 => to_unsigned(495, 12), 1552 => to_unsigned(3620, 12), 1553 => to_unsigned(485, 12), 1554 => to_unsigned(2133, 12), 1555 => to_unsigned(3966, 12), 1556 => to_unsigned(682, 12), 1557 => to_unsigned(3136, 12), 1558 => to_unsigned(3410, 12), 1559 => to_unsigned(3347, 12), 1560 => to_unsigned(698, 12), 1561 => to_unsigned(2572, 12), 1562 => to_unsigned(3421, 12), 1563 => to_unsigned(3456, 12), 1564 => to_unsigned(454, 12), 1565 => to_unsigned(3562, 12), 1566 => to_unsigned(1898, 12), 1567 => to_unsigned(3347, 12), 1568 => to_unsigned(3977, 12), 1569 => to_unsigned(2448, 12), 1570 => to_unsigned(142, 12), 1571 => to_unsigned(61, 12), 1572 => to_unsigned(1650, 12), 1573 => to_unsigned(3777, 12), 1574 => to_unsigned(285, 12), 1575 => to_unsigned(817, 12), 1576 => to_unsigned(147, 12), 1577 => to_unsigned(1045, 12), 1578 => to_unsigned(3642, 12), 1579 => to_unsigned(3839, 12), 1580 => to_unsigned(920, 12), 1581 => to_unsigned(3692, 12), 1582 => to_unsigned(3156, 12), 1583 => to_unsigned(2269, 12), 1584 => to_unsigned(627, 12), 1585 => to_unsigned(550, 12), 1586 => to_unsigned(581, 12), 1587 => to_unsigned(2641, 12), 1588 => to_unsigned(1672, 12), 1589 => to_unsigned(2222, 12), 1590 => to_unsigned(3827, 12), 1591 => to_unsigned(1375, 12), 1592 => to_unsigned(3947, 12), 1593 => to_unsigned(2654, 12), 1594 => to_unsigned(4066, 12), 1595 => to_unsigned(3068, 12), 1596 => to_unsigned(597, 12), 1597 => to_unsigned(3237, 12), 1598 => to_unsigned(303, 12), 1599 => to_unsigned(2678, 12), 1600 => to_unsigned(2520, 12), 1601 => to_unsigned(1846, 12), 1602 => to_unsigned(2530, 12), 1603 => to_unsigned(1842, 12), 1604 => to_unsigned(3066, 12), 1605 => to_unsigned(3587, 12), 1606 => to_unsigned(651, 12), 1607 => to_unsigned(383, 12), 1608 => to_unsigned(671, 12), 1609 => to_unsigned(879, 12), 1610 => to_unsigned(3730, 12), 1611 => to_unsigned(538, 12), 1612 => to_unsigned(2468, 12), 1613 => to_unsigned(3048, 12), 1614 => to_unsigned(3194, 12), 1615 => to_unsigned(3689, 12), 1616 => to_unsigned(3768, 12), 1617 => to_unsigned(2622, 12), 1618 => to_unsigned(1301, 12), 1619 => to_unsigned(2142, 12), 1620 => to_unsigned(2881, 12), 1621 => to_unsigned(2285, 12), 1622 => to_unsigned(1461, 12), 1623 => to_unsigned(2971, 12), 1624 => to_unsigned(2348, 12), 1625 => to_unsigned(525, 12), 1626 => to_unsigned(2962, 12), 1627 => to_unsigned(1909, 12), 1628 => to_unsigned(2883, 12), 1629 => to_unsigned(3094, 12), 1630 => to_unsigned(3056, 12), 1631 => to_unsigned(1403, 12), 1632 => to_unsigned(1764, 12), 1633 => to_unsigned(1135, 12), 1634 => to_unsigned(3297, 12), 1635 => to_unsigned(2835, 12), 1636 => to_unsigned(119, 12), 1637 => to_unsigned(478, 12), 1638 => to_unsigned(310, 12), 1639 => to_unsigned(2704, 12), 1640 => to_unsigned(1679, 12), 1641 => to_unsigned(4015, 12), 1642 => to_unsigned(2206, 12), 1643 => to_unsigned(256, 12), 1644 => to_unsigned(938, 12), 1645 => to_unsigned(3707, 12), 1646 => to_unsigned(16, 12), 1647 => to_unsigned(727, 12), 1648 => to_unsigned(1488, 12), 1649 => to_unsigned(204, 12), 1650 => to_unsigned(2876, 12), 1651 => to_unsigned(3689, 12), 1652 => to_unsigned(3967, 12), 1653 => to_unsigned(2734, 12), 1654 => to_unsigned(448, 12), 1655 => to_unsigned(1653, 12), 1656 => to_unsigned(2551, 12), 1657 => to_unsigned(2666, 12), 1658 => to_unsigned(2926, 12), 1659 => to_unsigned(256, 12), 1660 => to_unsigned(3905, 12), 1661 => to_unsigned(2715, 12), 1662 => to_unsigned(1570, 12), 1663 => to_unsigned(534, 12), 1664 => to_unsigned(4018, 12), 1665 => to_unsigned(864, 12), 1666 => to_unsigned(3052, 12), 1667 => to_unsigned(3979, 12), 1668 => to_unsigned(711, 12), 1669 => to_unsigned(2157, 12), 1670 => to_unsigned(1372, 12), 1671 => to_unsigned(3699, 12), 1672 => to_unsigned(160, 12), 1673 => to_unsigned(1121, 12), 1674 => to_unsigned(921, 12), 1675 => to_unsigned(374, 12), 1676 => to_unsigned(3610, 12), 1677 => to_unsigned(3205, 12), 1678 => to_unsigned(1681, 12), 1679 => to_unsigned(3170, 12), 1680 => to_unsigned(3256, 12), 1681 => to_unsigned(3494, 12), 1682 => to_unsigned(260, 12), 1683 => to_unsigned(2479, 12), 1684 => to_unsigned(1020, 12), 1685 => to_unsigned(3122, 12), 1686 => to_unsigned(3954, 12), 1687 => to_unsigned(428, 12), 1688 => to_unsigned(2157, 12), 1689 => to_unsigned(2774, 12), 1690 => to_unsigned(27, 12), 1691 => to_unsigned(3002, 12), 1692 => to_unsigned(1344, 12), 1693 => to_unsigned(2484, 12), 1694 => to_unsigned(3458, 12), 1695 => to_unsigned(3650, 12), 1696 => to_unsigned(1526, 12), 1697 => to_unsigned(148, 12), 1698 => to_unsigned(2360, 12), 1699 => to_unsigned(3027, 12), 1700 => to_unsigned(1822, 12), 1701 => to_unsigned(3100, 12), 1702 => to_unsigned(3168, 12), 1703 => to_unsigned(1819, 12), 1704 => to_unsigned(1327, 12), 1705 => to_unsigned(479, 12), 1706 => to_unsigned(1854, 12), 1707 => to_unsigned(3940, 12), 1708 => to_unsigned(740, 12), 1709 => to_unsigned(2890, 12), 1710 => to_unsigned(2409, 12), 1711 => to_unsigned(3244, 12), 1712 => to_unsigned(3874, 12), 1713 => to_unsigned(3957, 12), 1714 => to_unsigned(1598, 12), 1715 => to_unsigned(3051, 12), 1716 => to_unsigned(284, 12), 1717 => to_unsigned(3276, 12), 1718 => to_unsigned(2494, 12), 1719 => to_unsigned(3259, 12), 1720 => to_unsigned(2043, 12), 1721 => to_unsigned(714, 12), 1722 => to_unsigned(904, 12), 1723 => to_unsigned(1666, 12), 1724 => to_unsigned(61, 12), 1725 => to_unsigned(1694, 12), 1726 => to_unsigned(2162, 12), 1727 => to_unsigned(2921, 12), 1728 => to_unsigned(203, 12), 1729 => to_unsigned(2833, 12), 1730 => to_unsigned(1429, 12), 1731 => to_unsigned(2086, 12), 1732 => to_unsigned(2256, 12), 1733 => to_unsigned(2488, 12), 1734 => to_unsigned(594, 12), 1735 => to_unsigned(1708, 12), 1736 => to_unsigned(2853, 12), 1737 => to_unsigned(1899, 12), 1738 => to_unsigned(1496, 12), 1739 => to_unsigned(3830, 12), 1740 => to_unsigned(2476, 12), 1741 => to_unsigned(3180, 12), 1742 => to_unsigned(1865, 12), 1743 => to_unsigned(1511, 12), 1744 => to_unsigned(229, 12), 1745 => to_unsigned(3119, 12), 1746 => to_unsigned(2160, 12), 1747 => to_unsigned(1365, 12), 1748 => to_unsigned(3667, 12), 1749 => to_unsigned(1854, 12), 1750 => to_unsigned(636, 12), 1751 => to_unsigned(3264, 12), 1752 => to_unsigned(2094, 12), 1753 => to_unsigned(972, 12), 1754 => to_unsigned(3227, 12), 1755 => to_unsigned(99, 12), 1756 => to_unsigned(1329, 12), 1757 => to_unsigned(3528, 12), 1758 => to_unsigned(3532, 12), 1759 => to_unsigned(1548, 12), 1760 => to_unsigned(2416, 12), 1761 => to_unsigned(22, 12), 1762 => to_unsigned(1121, 12), 1763 => to_unsigned(1740, 12), 1764 => to_unsigned(3774, 12), 1765 => to_unsigned(518, 12), 1766 => to_unsigned(2027, 12), 1767 => to_unsigned(2517, 12), 1768 => to_unsigned(3724, 12), 1769 => to_unsigned(3925, 12), 1770 => to_unsigned(429, 12), 1771 => to_unsigned(1164, 12), 1772 => to_unsigned(379, 12), 1773 => to_unsigned(1387, 12), 1774 => to_unsigned(1581, 12), 1775 => to_unsigned(1198, 12), 1776 => to_unsigned(1104, 12), 1777 => to_unsigned(1949, 12), 1778 => to_unsigned(1777, 12), 1779 => to_unsigned(669, 12), 1780 => to_unsigned(1921, 12), 1781 => to_unsigned(2174, 12), 1782 => to_unsigned(2619, 12), 1783 => to_unsigned(3042, 12), 1784 => to_unsigned(2332, 12), 1785 => to_unsigned(1206, 12), 1786 => to_unsigned(1385, 12), 1787 => to_unsigned(3749, 12), 1788 => to_unsigned(3090, 12), 1789 => to_unsigned(92, 12), 1790 => to_unsigned(3630, 12), 1791 => to_unsigned(3536, 12), 1792 => to_unsigned(3824, 12), 1793 => to_unsigned(3428, 12), 1794 => to_unsigned(137, 12), 1795 => to_unsigned(3993, 12), 1796 => to_unsigned(225, 12), 1797 => to_unsigned(2584, 12), 1798 => to_unsigned(215, 12), 1799 => to_unsigned(1661, 12), 1800 => to_unsigned(2241, 12), 1801 => to_unsigned(1132, 12), 1802 => to_unsigned(2540, 12), 1803 => to_unsigned(2504, 12), 1804 => to_unsigned(3412, 12), 1805 => to_unsigned(1758, 12), 1806 => to_unsigned(3517, 12), 1807 => to_unsigned(2331, 12), 1808 => to_unsigned(2587, 12), 1809 => to_unsigned(3627, 12), 1810 => to_unsigned(1520, 12), 1811 => to_unsigned(460, 12), 1812 => to_unsigned(993, 12), 1813 => to_unsigned(689, 12), 1814 => to_unsigned(3838, 12), 1815 => to_unsigned(329, 12), 1816 => to_unsigned(3098, 12), 1817 => to_unsigned(173, 12), 1818 => to_unsigned(2694, 12), 1819 => to_unsigned(1486, 12), 1820 => to_unsigned(599, 12), 1821 => to_unsigned(201, 12), 1822 => to_unsigned(1538, 12), 1823 => to_unsigned(1393, 12), 1824 => to_unsigned(2868, 12), 1825 => to_unsigned(2916, 12), 1826 => to_unsigned(1778, 12), 1827 => to_unsigned(2020, 12), 1828 => to_unsigned(1702, 12), 1829 => to_unsigned(3886, 12), 1830 => to_unsigned(2643, 12), 1831 => to_unsigned(2750, 12), 1832 => to_unsigned(2877, 12), 1833 => to_unsigned(1948, 12), 1834 => to_unsigned(1874, 12), 1835 => to_unsigned(4020, 12), 1836 => to_unsigned(3284, 12), 1837 => to_unsigned(1278, 12), 1838 => to_unsigned(3714, 12), 1839 => to_unsigned(2112, 12), 1840 => to_unsigned(1626, 12), 1841 => to_unsigned(1500, 12), 1842 => to_unsigned(3997, 12), 1843 => to_unsigned(2174, 12), 1844 => to_unsigned(1726, 12), 1845 => to_unsigned(3368, 12), 1846 => to_unsigned(317, 12), 1847 => to_unsigned(3778, 12), 1848 => to_unsigned(3897, 12), 1849 => to_unsigned(2059, 12), 1850 => to_unsigned(1562, 12), 1851 => to_unsigned(2348, 12), 1852 => to_unsigned(960, 12), 1853 => to_unsigned(3486, 12), 1854 => to_unsigned(1424, 12), 1855 => to_unsigned(565, 12), 1856 => to_unsigned(1173, 12), 1857 => to_unsigned(3784, 12), 1858 => to_unsigned(824, 12), 1859 => to_unsigned(2024, 12), 1860 => to_unsigned(3467, 12), 1861 => to_unsigned(2200, 12), 1862 => to_unsigned(2170, 12), 1863 => to_unsigned(559, 12), 1864 => to_unsigned(2867, 12), 1865 => to_unsigned(3409, 12), 1866 => to_unsigned(2980, 12), 1867 => to_unsigned(879, 12), 1868 => to_unsigned(2232, 12), 1869 => to_unsigned(2531, 12), 1870 => to_unsigned(3596, 12), 1871 => to_unsigned(656, 12), 1872 => to_unsigned(2196, 12), 1873 => to_unsigned(3022, 12), 1874 => to_unsigned(3487, 12), 1875 => to_unsigned(3366, 12), 1876 => to_unsigned(2914, 12), 1877 => to_unsigned(1398, 12), 1878 => to_unsigned(3556, 12), 1879 => to_unsigned(2901, 12), 1880 => to_unsigned(4050, 12), 1881 => to_unsigned(690, 12), 1882 => to_unsigned(4001, 12), 1883 => to_unsigned(174, 12), 1884 => to_unsigned(2624, 12), 1885 => to_unsigned(783, 12), 1886 => to_unsigned(1919, 12), 1887 => to_unsigned(2293, 12), 1888 => to_unsigned(2013, 12), 1889 => to_unsigned(3892, 12), 1890 => to_unsigned(2904, 12), 1891 => to_unsigned(623, 12), 1892 => to_unsigned(314, 12), 1893 => to_unsigned(1680, 12), 1894 => to_unsigned(3570, 12), 1895 => to_unsigned(2048, 12), 1896 => to_unsigned(3571, 12), 1897 => to_unsigned(2922, 12), 1898 => to_unsigned(920, 12), 1899 => to_unsigned(1238, 12), 1900 => to_unsigned(985, 12), 1901 => to_unsigned(937, 12), 1902 => to_unsigned(3307, 12), 1903 => to_unsigned(3143, 12), 1904 => to_unsigned(2817, 12), 1905 => to_unsigned(2035, 12), 1906 => to_unsigned(656, 12), 1907 => to_unsigned(3790, 12), 1908 => to_unsigned(2071, 12), 1909 => to_unsigned(3197, 12), 1910 => to_unsigned(1164, 12), 1911 => to_unsigned(565, 12), 1912 => to_unsigned(3730, 12), 1913 => to_unsigned(3177, 12), 1914 => to_unsigned(3445, 12), 1915 => to_unsigned(2642, 12), 1916 => to_unsigned(676, 12), 1917 => to_unsigned(2260, 12), 1918 => to_unsigned(835, 12), 1919 => to_unsigned(3684, 12), 1920 => to_unsigned(3765, 12), 1921 => to_unsigned(2231, 12), 1922 => to_unsigned(1895, 12), 1923 => to_unsigned(3217, 12), 1924 => to_unsigned(382, 12), 1925 => to_unsigned(371, 12), 1926 => to_unsigned(854, 12), 1927 => to_unsigned(3282, 12), 1928 => to_unsigned(291, 12), 1929 => to_unsigned(996, 12), 1930 => to_unsigned(1058, 12), 1931 => to_unsigned(4089, 12), 1932 => to_unsigned(1540, 12), 1933 => to_unsigned(2398, 12), 1934 => to_unsigned(1578, 12), 1935 => to_unsigned(1077, 12), 1936 => to_unsigned(353, 12), 1937 => to_unsigned(119, 12), 1938 => to_unsigned(1511, 12), 1939 => to_unsigned(1551, 12), 1940 => to_unsigned(3355, 12), 1941 => to_unsigned(3141, 12), 1942 => to_unsigned(2391, 12), 1943 => to_unsigned(467, 12), 1944 => to_unsigned(633, 12), 1945 => to_unsigned(269, 12), 1946 => to_unsigned(2167, 12), 1947 => to_unsigned(1593, 12), 1948 => to_unsigned(3860, 12), 1949 => to_unsigned(3482, 12), 1950 => to_unsigned(1375, 12), 1951 => to_unsigned(2703, 12), 1952 => to_unsigned(2513, 12), 1953 => to_unsigned(1958, 12), 1954 => to_unsigned(338, 12), 1955 => to_unsigned(1897, 12), 1956 => to_unsigned(4006, 12), 1957 => to_unsigned(2064, 12), 1958 => to_unsigned(217, 12), 1959 => to_unsigned(1962, 12), 1960 => to_unsigned(3341, 12), 1961 => to_unsigned(2798, 12), 1962 => to_unsigned(3375, 12), 1963 => to_unsigned(1163, 12), 1964 => to_unsigned(3627, 12), 1965 => to_unsigned(2450, 12), 1966 => to_unsigned(3729, 12), 1967 => to_unsigned(4062, 12), 1968 => to_unsigned(1380, 12), 1969 => to_unsigned(1241, 12), 1970 => to_unsigned(2053, 12), 1971 => to_unsigned(1204, 12), 1972 => to_unsigned(3160, 12), 1973 => to_unsigned(2149, 12), 1974 => to_unsigned(1461, 12), 1975 => to_unsigned(2980, 12), 1976 => to_unsigned(515, 12), 1977 => to_unsigned(2690, 12), 1978 => to_unsigned(2012, 12), 1979 => to_unsigned(1793, 12), 1980 => to_unsigned(1811, 12), 1981 => to_unsigned(242, 12), 1982 => to_unsigned(797, 12), 1983 => to_unsigned(246, 12), 1984 => to_unsigned(553, 12), 1985 => to_unsigned(3684, 12), 1986 => to_unsigned(3634, 12), 1987 => to_unsigned(94, 12), 1988 => to_unsigned(940, 12), 1989 => to_unsigned(3904, 12), 1990 => to_unsigned(1119, 12), 1991 => to_unsigned(3902, 12), 1992 => to_unsigned(894, 12), 1993 => to_unsigned(85, 12), 1994 => to_unsigned(1499, 12), 1995 => to_unsigned(2900, 12), 1996 => to_unsigned(2544, 12), 1997 => to_unsigned(3826, 12), 1998 => to_unsigned(3395, 12), 1999 => to_unsigned(768, 12), 2000 => to_unsigned(2796, 12), 2001 => to_unsigned(1886, 12), 2002 => to_unsigned(2351, 12), 2003 => to_unsigned(3350, 12), 2004 => to_unsigned(3272, 12), 2005 => to_unsigned(73, 12), 2006 => to_unsigned(1126, 12), 2007 => to_unsigned(501, 12), 2008 => to_unsigned(220, 12), 2009 => to_unsigned(3193, 12), 2010 => to_unsigned(2183, 12), 2011 => to_unsigned(1378, 12), 2012 => to_unsigned(2220, 12), 2013 => to_unsigned(2660, 12), 2014 => to_unsigned(2923, 12), 2015 => to_unsigned(1021, 12), 2016 => to_unsigned(973, 12), 2017 => to_unsigned(730, 12), 2018 => to_unsigned(2234, 12), 2019 => to_unsigned(656, 12), 2020 => to_unsigned(4028, 12), 2021 => to_unsigned(1395, 12), 2022 => to_unsigned(2309, 12), 2023 => to_unsigned(2350, 12), 2024 => to_unsigned(1261, 12), 2025 => to_unsigned(1021, 12), 2026 => to_unsigned(3181, 12), 2027 => to_unsigned(2118, 12), 2028 => to_unsigned(2730, 12), 2029 => to_unsigned(2476, 12), 2030 => to_unsigned(717, 12), 2031 => to_unsigned(3417, 12), 2032 => to_unsigned(406, 12), 2033 => to_unsigned(2235, 12), 2034 => to_unsigned(1868, 12), 2035 => to_unsigned(567, 12), 2036 => to_unsigned(152, 12), 2037 => to_unsigned(3197, 12), 2038 => to_unsigned(2820, 12), 2039 => to_unsigned(16, 12), 2040 => to_unsigned(444, 12), 2041 => to_unsigned(1095, 12), 2042 => to_unsigned(1572, 12), 2043 => to_unsigned(3034, 12), 2044 => to_unsigned(473, 12), 2045 => to_unsigned(2806, 12), 2046 => to_unsigned(3261, 12), 2047 => to_unsigned(894, 12)),
            4 => (0 => to_unsigned(409, 12), 1 => to_unsigned(1631, 12), 2 => to_unsigned(2650, 12), 3 => to_unsigned(2176, 12), 4 => to_unsigned(2608, 12), 5 => to_unsigned(1905, 12), 6 => to_unsigned(1534, 12), 7 => to_unsigned(3110, 12), 8 => to_unsigned(735, 12), 9 => to_unsigned(1674, 12), 10 => to_unsigned(3494, 12), 11 => to_unsigned(770, 12), 12 => to_unsigned(273, 12), 13 => to_unsigned(3332, 12), 14 => to_unsigned(3899, 12), 15 => to_unsigned(2868, 12), 16 => to_unsigned(3041, 12), 17 => to_unsigned(1539, 12), 18 => to_unsigned(3583, 12), 19 => to_unsigned(2485, 12), 20 => to_unsigned(466, 12), 21 => to_unsigned(971, 12), 22 => to_unsigned(515, 12), 23 => to_unsigned(519, 12), 24 => to_unsigned(1762, 12), 25 => to_unsigned(1150, 12), 26 => to_unsigned(1483, 12), 27 => to_unsigned(2350, 12), 28 => to_unsigned(3006, 12), 29 => to_unsigned(612, 12), 30 => to_unsigned(290, 12), 31 => to_unsigned(1840, 12), 32 => to_unsigned(1399, 12), 33 => to_unsigned(1330, 12), 34 => to_unsigned(757, 12), 35 => to_unsigned(696, 12), 36 => to_unsigned(3379, 12), 37 => to_unsigned(3860, 12), 38 => to_unsigned(3213, 12), 39 => to_unsigned(2764, 12), 40 => to_unsigned(559, 12), 41 => to_unsigned(1527, 12), 42 => to_unsigned(1179, 12), 43 => to_unsigned(776, 12), 44 => to_unsigned(1881, 12), 45 => to_unsigned(3252, 12), 46 => to_unsigned(1485, 12), 47 => to_unsigned(3713, 12), 48 => to_unsigned(543, 12), 49 => to_unsigned(1779, 12), 50 => to_unsigned(3214, 12), 51 => to_unsigned(2848, 12), 52 => to_unsigned(2997, 12), 53 => to_unsigned(2559, 12), 54 => to_unsigned(506, 12), 55 => to_unsigned(2981, 12), 56 => to_unsigned(2906, 12), 57 => to_unsigned(2712, 12), 58 => to_unsigned(2772, 12), 59 => to_unsigned(2231, 12), 60 => to_unsigned(273, 12), 61 => to_unsigned(1147, 12), 62 => to_unsigned(954, 12), 63 => to_unsigned(1242, 12), 64 => to_unsigned(972, 12), 65 => to_unsigned(301, 12), 66 => to_unsigned(1537, 12), 67 => to_unsigned(1154, 12), 68 => to_unsigned(3283, 12), 69 => to_unsigned(3482, 12), 70 => to_unsigned(1723, 12), 71 => to_unsigned(2085, 12), 72 => to_unsigned(3783, 12), 73 => to_unsigned(1430, 12), 74 => to_unsigned(1220, 12), 75 => to_unsigned(2421, 12), 76 => to_unsigned(1242, 12), 77 => to_unsigned(3815, 12), 78 => to_unsigned(3370, 12), 79 => to_unsigned(2189, 12), 80 => to_unsigned(3396, 12), 81 => to_unsigned(2902, 12), 82 => to_unsigned(1460, 12), 83 => to_unsigned(2596, 12), 84 => to_unsigned(1355, 12), 85 => to_unsigned(1675, 12), 86 => to_unsigned(1480, 12), 87 => to_unsigned(1015, 12), 88 => to_unsigned(4014, 12), 89 => to_unsigned(1067, 12), 90 => to_unsigned(1843, 12), 91 => to_unsigned(1126, 12), 92 => to_unsigned(3688, 12), 93 => to_unsigned(1384, 12), 94 => to_unsigned(3195, 12), 95 => to_unsigned(2780, 12), 96 => to_unsigned(1630, 12), 97 => to_unsigned(1239, 12), 98 => to_unsigned(2318, 12), 99 => to_unsigned(250, 12), 100 => to_unsigned(3391, 12), 101 => to_unsigned(2207, 12), 102 => to_unsigned(2750, 12), 103 => to_unsigned(3286, 12), 104 => to_unsigned(2410, 12), 105 => to_unsigned(2705, 12), 106 => to_unsigned(1268, 12), 107 => to_unsigned(110, 12), 108 => to_unsigned(2767, 12), 109 => to_unsigned(3700, 12), 110 => to_unsigned(306, 12), 111 => to_unsigned(804, 12), 112 => to_unsigned(1357, 12), 113 => to_unsigned(961, 12), 114 => to_unsigned(264, 12), 115 => to_unsigned(2493, 12), 116 => to_unsigned(3326, 12), 117 => to_unsigned(525, 12), 118 => to_unsigned(2768, 12), 119 => to_unsigned(529, 12), 120 => to_unsigned(3917, 12), 121 => to_unsigned(3836, 12), 122 => to_unsigned(826, 12), 123 => to_unsigned(1554, 12), 124 => to_unsigned(3050, 12), 125 => to_unsigned(2333, 12), 126 => to_unsigned(1062, 12), 127 => to_unsigned(4077, 12), 128 => to_unsigned(910, 12), 129 => to_unsigned(1455, 12), 130 => to_unsigned(3429, 12), 131 => to_unsigned(3892, 12), 132 => to_unsigned(3567, 12), 133 => to_unsigned(3495, 12), 134 => to_unsigned(3062, 12), 135 => to_unsigned(393, 12), 136 => to_unsigned(1343, 12), 137 => to_unsigned(1013, 12), 138 => to_unsigned(3847, 12), 139 => to_unsigned(3025, 12), 140 => to_unsigned(1982, 12), 141 => to_unsigned(225, 12), 142 => to_unsigned(924, 12), 143 => to_unsigned(3653, 12), 144 => to_unsigned(2016, 12), 145 => to_unsigned(3434, 12), 146 => to_unsigned(719, 12), 147 => to_unsigned(1077, 12), 148 => to_unsigned(769, 12), 149 => to_unsigned(789, 12), 150 => to_unsigned(2472, 12), 151 => to_unsigned(3588, 12), 152 => to_unsigned(1508, 12), 153 => to_unsigned(2277, 12), 154 => to_unsigned(4077, 12), 155 => to_unsigned(1109, 12), 156 => to_unsigned(1196, 12), 157 => to_unsigned(3035, 12), 158 => to_unsigned(759, 12), 159 => to_unsigned(2140, 12), 160 => to_unsigned(864, 12), 161 => to_unsigned(547, 12), 162 => to_unsigned(270, 12), 163 => to_unsigned(1232, 12), 164 => to_unsigned(1971, 12), 165 => to_unsigned(2730, 12), 166 => to_unsigned(3241, 12), 167 => to_unsigned(4041, 12), 168 => to_unsigned(1269, 12), 169 => to_unsigned(2191, 12), 170 => to_unsigned(2132, 12), 171 => to_unsigned(539, 12), 172 => to_unsigned(566, 12), 173 => to_unsigned(2992, 12), 174 => to_unsigned(665, 12), 175 => to_unsigned(2640, 12), 176 => to_unsigned(3520, 12), 177 => to_unsigned(2560, 12), 178 => to_unsigned(1229, 12), 179 => to_unsigned(2041, 12), 180 => to_unsigned(355, 12), 181 => to_unsigned(2045, 12), 182 => to_unsigned(2438, 12), 183 => to_unsigned(1771, 12), 184 => to_unsigned(2232, 12), 185 => to_unsigned(743, 12), 186 => to_unsigned(383, 12), 187 => to_unsigned(1688, 12), 188 => to_unsigned(32, 12), 189 => to_unsigned(1265, 12), 190 => to_unsigned(2304, 12), 191 => to_unsigned(552, 12), 192 => to_unsigned(1208, 12), 193 => to_unsigned(2038, 12), 194 => to_unsigned(228, 12), 195 => to_unsigned(3622, 12), 196 => to_unsigned(697, 12), 197 => to_unsigned(1229, 12), 198 => to_unsigned(771, 12), 199 => to_unsigned(3750, 12), 200 => to_unsigned(2761, 12), 201 => to_unsigned(3132, 12), 202 => to_unsigned(1420, 12), 203 => to_unsigned(3318, 12), 204 => to_unsigned(2636, 12), 205 => to_unsigned(1058, 12), 206 => to_unsigned(3918, 12), 207 => to_unsigned(2279, 12), 208 => to_unsigned(973, 12), 209 => to_unsigned(3327, 12), 210 => to_unsigned(3940, 12), 211 => to_unsigned(1541, 12), 212 => to_unsigned(2368, 12), 213 => to_unsigned(2669, 12), 214 => to_unsigned(3854, 12), 215 => to_unsigned(2457, 12), 216 => to_unsigned(474, 12), 217 => to_unsigned(3951, 12), 218 => to_unsigned(1203, 12), 219 => to_unsigned(2042, 12), 220 => to_unsigned(2550, 12), 221 => to_unsigned(1724, 12), 222 => to_unsigned(3193, 12), 223 => to_unsigned(2061, 12), 224 => to_unsigned(1430, 12), 225 => to_unsigned(3066, 12), 226 => to_unsigned(1379, 12), 227 => to_unsigned(1102, 12), 228 => to_unsigned(464, 12), 229 => to_unsigned(3854, 12), 230 => to_unsigned(1147, 12), 231 => to_unsigned(145, 12), 232 => to_unsigned(3665, 12), 233 => to_unsigned(2820, 12), 234 => to_unsigned(380, 12), 235 => to_unsigned(52, 12), 236 => to_unsigned(400, 12), 237 => to_unsigned(1597, 12), 238 => to_unsigned(2850, 12), 239 => to_unsigned(3682, 12), 240 => to_unsigned(1795, 12), 241 => to_unsigned(380, 12), 242 => to_unsigned(2381, 12), 243 => to_unsigned(520, 12), 244 => to_unsigned(3555, 12), 245 => to_unsigned(315, 12), 246 => to_unsigned(2240, 12), 247 => to_unsigned(3867, 12), 248 => to_unsigned(1371, 12), 249 => to_unsigned(73, 12), 250 => to_unsigned(2753, 12), 251 => to_unsigned(1706, 12), 252 => to_unsigned(999, 12), 253 => to_unsigned(1827, 12), 254 => to_unsigned(1955, 12), 255 => to_unsigned(229, 12), 256 => to_unsigned(3811, 12), 257 => to_unsigned(2712, 12), 258 => to_unsigned(1814, 12), 259 => to_unsigned(2533, 12), 260 => to_unsigned(2585, 12), 261 => to_unsigned(1220, 12), 262 => to_unsigned(2061, 12), 263 => to_unsigned(894, 12), 264 => to_unsigned(333, 12), 265 => to_unsigned(1366, 12), 266 => to_unsigned(1962, 12), 267 => to_unsigned(150, 12), 268 => to_unsigned(680, 12), 269 => to_unsigned(999, 12), 270 => to_unsigned(291, 12), 271 => to_unsigned(524, 12), 272 => to_unsigned(400, 12), 273 => to_unsigned(471, 12), 274 => to_unsigned(1980, 12), 275 => to_unsigned(451, 12), 276 => to_unsigned(3786, 12), 277 => to_unsigned(423, 12), 278 => to_unsigned(2442, 12), 279 => to_unsigned(3345, 12), 280 => to_unsigned(1367, 12), 281 => to_unsigned(1303, 12), 282 => to_unsigned(3898, 12), 283 => to_unsigned(478, 12), 284 => to_unsigned(2711, 12), 285 => to_unsigned(3803, 12), 286 => to_unsigned(1034, 12), 287 => to_unsigned(2580, 12), 288 => to_unsigned(9, 12), 289 => to_unsigned(1285, 12), 290 => to_unsigned(3934, 12), 291 => to_unsigned(2781, 12), 292 => to_unsigned(2139, 12), 293 => to_unsigned(1938, 12), 294 => to_unsigned(755, 12), 295 => to_unsigned(327, 12), 296 => to_unsigned(2154, 12), 297 => to_unsigned(3918, 12), 298 => to_unsigned(2688, 12), 299 => to_unsigned(1011, 12), 300 => to_unsigned(1152, 12), 301 => to_unsigned(2558, 12), 302 => to_unsigned(138, 12), 303 => to_unsigned(1527, 12), 304 => to_unsigned(2064, 12), 305 => to_unsigned(2131, 12), 306 => to_unsigned(688, 12), 307 => to_unsigned(1230, 12), 308 => to_unsigned(3376, 12), 309 => to_unsigned(1322, 12), 310 => to_unsigned(232, 12), 311 => to_unsigned(1282, 12), 312 => to_unsigned(303, 12), 313 => to_unsigned(2944, 12), 314 => to_unsigned(1541, 12), 315 => to_unsigned(1586, 12), 316 => to_unsigned(3413, 12), 317 => to_unsigned(2681, 12), 318 => to_unsigned(3160, 12), 319 => to_unsigned(173, 12), 320 => to_unsigned(2430, 12), 321 => to_unsigned(2404, 12), 322 => to_unsigned(1087, 12), 323 => to_unsigned(300, 12), 324 => to_unsigned(1321, 12), 325 => to_unsigned(3109, 12), 326 => to_unsigned(1929, 12), 327 => to_unsigned(989, 12), 328 => to_unsigned(2141, 12), 329 => to_unsigned(2384, 12), 330 => to_unsigned(3034, 12), 331 => to_unsigned(3446, 12), 332 => to_unsigned(1859, 12), 333 => to_unsigned(4026, 12), 334 => to_unsigned(3863, 12), 335 => to_unsigned(901, 12), 336 => to_unsigned(3499, 12), 337 => to_unsigned(476, 12), 338 => to_unsigned(1739, 12), 339 => to_unsigned(2803, 12), 340 => to_unsigned(2866, 12), 341 => to_unsigned(2203, 12), 342 => to_unsigned(2711, 12), 343 => to_unsigned(2758, 12), 344 => to_unsigned(1244, 12), 345 => to_unsigned(2056, 12), 346 => to_unsigned(204, 12), 347 => to_unsigned(3699, 12), 348 => to_unsigned(3990, 12), 349 => to_unsigned(3540, 12), 350 => to_unsigned(549, 12), 351 => to_unsigned(4063, 12), 352 => to_unsigned(2039, 12), 353 => to_unsigned(2401, 12), 354 => to_unsigned(3845, 12), 355 => to_unsigned(1183, 12), 356 => to_unsigned(3809, 12), 357 => to_unsigned(1288, 12), 358 => to_unsigned(2875, 12), 359 => to_unsigned(416, 12), 360 => to_unsigned(1974, 12), 361 => to_unsigned(1982, 12), 362 => to_unsigned(1729, 12), 363 => to_unsigned(1978, 12), 364 => to_unsigned(1554, 12), 365 => to_unsigned(1245, 12), 366 => to_unsigned(3694, 12), 367 => to_unsigned(1373, 12), 368 => to_unsigned(1498, 12), 369 => to_unsigned(621, 12), 370 => to_unsigned(581, 12), 371 => to_unsigned(1477, 12), 372 => to_unsigned(1697, 12), 373 => to_unsigned(1208, 12), 374 => to_unsigned(2086, 12), 375 => to_unsigned(3072, 12), 376 => to_unsigned(622, 12), 377 => to_unsigned(3476, 12), 378 => to_unsigned(3183, 12), 379 => to_unsigned(939, 12), 380 => to_unsigned(1761, 12), 381 => to_unsigned(2446, 12), 382 => to_unsigned(2471, 12), 383 => to_unsigned(4022, 12), 384 => to_unsigned(450, 12), 385 => to_unsigned(109, 12), 386 => to_unsigned(2843, 12), 387 => to_unsigned(648, 12), 388 => to_unsigned(1189, 12), 389 => to_unsigned(19, 12), 390 => to_unsigned(2882, 12), 391 => to_unsigned(3719, 12), 392 => to_unsigned(547, 12), 393 => to_unsigned(3693, 12), 394 => to_unsigned(818, 12), 395 => to_unsigned(871, 12), 396 => to_unsigned(782, 12), 397 => to_unsigned(2081, 12), 398 => to_unsigned(967, 12), 399 => to_unsigned(183, 12), 400 => to_unsigned(1715, 12), 401 => to_unsigned(3701, 12), 402 => to_unsigned(2421, 12), 403 => to_unsigned(2192, 12), 404 => to_unsigned(24, 12), 405 => to_unsigned(2974, 12), 406 => to_unsigned(1510, 12), 407 => to_unsigned(1580, 12), 408 => to_unsigned(3463, 12), 409 => to_unsigned(2223, 12), 410 => to_unsigned(101, 12), 411 => to_unsigned(745, 12), 412 => to_unsigned(1004, 12), 413 => to_unsigned(211, 12), 414 => to_unsigned(399, 12), 415 => to_unsigned(3931, 12), 416 => to_unsigned(2378, 12), 417 => to_unsigned(3409, 12), 418 => to_unsigned(95, 12), 419 => to_unsigned(60, 12), 420 => to_unsigned(2720, 12), 421 => to_unsigned(1910, 12), 422 => to_unsigned(2485, 12), 423 => to_unsigned(92, 12), 424 => to_unsigned(1535, 12), 425 => to_unsigned(490, 12), 426 => to_unsigned(2821, 12), 427 => to_unsigned(1498, 12), 428 => to_unsigned(3233, 12), 429 => to_unsigned(2805, 12), 430 => to_unsigned(126, 12), 431 => to_unsigned(3195, 12), 432 => to_unsigned(3507, 12), 433 => to_unsigned(933, 12), 434 => to_unsigned(1994, 12), 435 => to_unsigned(2743, 12), 436 => to_unsigned(3184, 12), 437 => to_unsigned(1030, 12), 438 => to_unsigned(1381, 12), 439 => to_unsigned(3295, 12), 440 => to_unsigned(2845, 12), 441 => to_unsigned(1623, 12), 442 => to_unsigned(557, 12), 443 => to_unsigned(3860, 12), 444 => to_unsigned(1149, 12), 445 => to_unsigned(3534, 12), 446 => to_unsigned(1986, 12), 447 => to_unsigned(3846, 12), 448 => to_unsigned(3732, 12), 449 => to_unsigned(1431, 12), 450 => to_unsigned(1902, 12), 451 => to_unsigned(1424, 12), 452 => to_unsigned(3412, 12), 453 => to_unsigned(2453, 12), 454 => to_unsigned(2605, 12), 455 => to_unsigned(3088, 12), 456 => to_unsigned(317, 12), 457 => to_unsigned(1282, 12), 458 => to_unsigned(3107, 12), 459 => to_unsigned(678, 12), 460 => to_unsigned(1735, 12), 461 => to_unsigned(2785, 12), 462 => to_unsigned(3029, 12), 463 => to_unsigned(305, 12), 464 => to_unsigned(1775, 12), 465 => to_unsigned(1866, 12), 466 => to_unsigned(622, 12), 467 => to_unsigned(443, 12), 468 => to_unsigned(1221, 12), 469 => to_unsigned(1301, 12), 470 => to_unsigned(2756, 12), 471 => to_unsigned(679, 12), 472 => to_unsigned(3381, 12), 473 => to_unsigned(2813, 12), 474 => to_unsigned(461, 12), 475 => to_unsigned(3536, 12), 476 => to_unsigned(3948, 12), 477 => to_unsigned(2524, 12), 478 => to_unsigned(1066, 12), 479 => to_unsigned(3469, 12), 480 => to_unsigned(3981, 12), 481 => to_unsigned(1139, 12), 482 => to_unsigned(1431, 12), 483 => to_unsigned(3012, 12), 484 => to_unsigned(2231, 12), 485 => to_unsigned(1727, 12), 486 => to_unsigned(2065, 12), 487 => to_unsigned(990, 12), 488 => to_unsigned(1995, 12), 489 => to_unsigned(401, 12), 490 => to_unsigned(1160, 12), 491 => to_unsigned(1081, 12), 492 => to_unsigned(3007, 12), 493 => to_unsigned(16, 12), 494 => to_unsigned(681, 12), 495 => to_unsigned(1200, 12), 496 => to_unsigned(3354, 12), 497 => to_unsigned(4066, 12), 498 => to_unsigned(1401, 12), 499 => to_unsigned(1124, 12), 500 => to_unsigned(699, 12), 501 => to_unsigned(448, 12), 502 => to_unsigned(941, 12), 503 => to_unsigned(1265, 12), 504 => to_unsigned(1160, 12), 505 => to_unsigned(3199, 12), 506 => to_unsigned(2427, 12), 507 => to_unsigned(3619, 12), 508 => to_unsigned(13, 12), 509 => to_unsigned(3540, 12), 510 => to_unsigned(865, 12), 511 => to_unsigned(849, 12), 512 => to_unsigned(1978, 12), 513 => to_unsigned(1094, 12), 514 => to_unsigned(1388, 12), 515 => to_unsigned(2321, 12), 516 => to_unsigned(2653, 12), 517 => to_unsigned(930, 12), 518 => to_unsigned(1439, 12), 519 => to_unsigned(84, 12), 520 => to_unsigned(3159, 12), 521 => to_unsigned(3560, 12), 522 => to_unsigned(4056, 12), 523 => to_unsigned(3531, 12), 524 => to_unsigned(1833, 12), 525 => to_unsigned(2514, 12), 526 => to_unsigned(2121, 12), 527 => to_unsigned(4041, 12), 528 => to_unsigned(625, 12), 529 => to_unsigned(2684, 12), 530 => to_unsigned(3357, 12), 531 => to_unsigned(2017, 12), 532 => to_unsigned(3310, 12), 533 => to_unsigned(1659, 12), 534 => to_unsigned(3295, 12), 535 => to_unsigned(4054, 12), 536 => to_unsigned(89, 12), 537 => to_unsigned(2750, 12), 538 => to_unsigned(5, 12), 539 => to_unsigned(3709, 12), 540 => to_unsigned(3368, 12), 541 => to_unsigned(1571, 12), 542 => to_unsigned(3885, 12), 543 => to_unsigned(1298, 12), 544 => to_unsigned(2262, 12), 545 => to_unsigned(1889, 12), 546 => to_unsigned(4046, 12), 547 => to_unsigned(2785, 12), 548 => to_unsigned(3943, 12), 549 => to_unsigned(678, 12), 550 => to_unsigned(389, 12), 551 => to_unsigned(1793, 12), 552 => to_unsigned(3077, 12), 553 => to_unsigned(486, 12), 554 => to_unsigned(1823, 12), 555 => to_unsigned(1505, 12), 556 => to_unsigned(168, 12), 557 => to_unsigned(1388, 12), 558 => to_unsigned(129, 12), 559 => to_unsigned(1492, 12), 560 => to_unsigned(3942, 12), 561 => to_unsigned(3183, 12), 562 => to_unsigned(2471, 12), 563 => to_unsigned(724, 12), 564 => to_unsigned(2829, 12), 565 => to_unsigned(427, 12), 566 => to_unsigned(1107, 12), 567 => to_unsigned(2539, 12), 568 => to_unsigned(1433, 12), 569 => to_unsigned(2360, 12), 570 => to_unsigned(3956, 12), 571 => to_unsigned(3644, 12), 572 => to_unsigned(316, 12), 573 => to_unsigned(3329, 12), 574 => to_unsigned(2796, 12), 575 => to_unsigned(2053, 12), 576 => to_unsigned(5, 12), 577 => to_unsigned(472, 12), 578 => to_unsigned(858, 12), 579 => to_unsigned(2169, 12), 580 => to_unsigned(3676, 12), 581 => to_unsigned(3362, 12), 582 => to_unsigned(756, 12), 583 => to_unsigned(3096, 12), 584 => to_unsigned(2388, 12), 585 => to_unsigned(2030, 12), 586 => to_unsigned(3025, 12), 587 => to_unsigned(823, 12), 588 => to_unsigned(2032, 12), 589 => to_unsigned(1595, 12), 590 => to_unsigned(3712, 12), 591 => to_unsigned(3362, 12), 592 => to_unsigned(2526, 12), 593 => to_unsigned(3827, 12), 594 => to_unsigned(2950, 12), 595 => to_unsigned(4024, 12), 596 => to_unsigned(1262, 12), 597 => to_unsigned(2116, 12), 598 => to_unsigned(1288, 12), 599 => to_unsigned(2323, 12), 600 => to_unsigned(2371, 12), 601 => to_unsigned(3488, 12), 602 => to_unsigned(1407, 12), 603 => to_unsigned(3651, 12), 604 => to_unsigned(615, 12), 605 => to_unsigned(3133, 12), 606 => to_unsigned(2970, 12), 607 => to_unsigned(2195, 12), 608 => to_unsigned(1228, 12), 609 => to_unsigned(896, 12), 610 => to_unsigned(981, 12), 611 => to_unsigned(3028, 12), 612 => to_unsigned(2865, 12), 613 => to_unsigned(2427, 12), 614 => to_unsigned(2154, 12), 615 => to_unsigned(3650, 12), 616 => to_unsigned(3328, 12), 617 => to_unsigned(3473, 12), 618 => to_unsigned(3616, 12), 619 => to_unsigned(3248, 12), 620 => to_unsigned(2850, 12), 621 => to_unsigned(2153, 12), 622 => to_unsigned(1925, 12), 623 => to_unsigned(3494, 12), 624 => to_unsigned(2354, 12), 625 => to_unsigned(1554, 12), 626 => to_unsigned(1720, 12), 627 => to_unsigned(1874, 12), 628 => to_unsigned(1248, 12), 629 => to_unsigned(2214, 12), 630 => to_unsigned(1752, 12), 631 => to_unsigned(960, 12), 632 => to_unsigned(3464, 12), 633 => to_unsigned(3425, 12), 634 => to_unsigned(1923, 12), 635 => to_unsigned(2732, 12), 636 => to_unsigned(2476, 12), 637 => to_unsigned(434, 12), 638 => to_unsigned(1595, 12), 639 => to_unsigned(2300, 12), 640 => to_unsigned(459, 12), 641 => to_unsigned(3640, 12), 642 => to_unsigned(2561, 12), 643 => to_unsigned(2601, 12), 644 => to_unsigned(1050, 12), 645 => to_unsigned(2904, 12), 646 => to_unsigned(1012, 12), 647 => to_unsigned(2491, 12), 648 => to_unsigned(3197, 12), 649 => to_unsigned(2454, 12), 650 => to_unsigned(3711, 12), 651 => to_unsigned(2029, 12), 652 => to_unsigned(2543, 12), 653 => to_unsigned(1476, 12), 654 => to_unsigned(397, 12), 655 => to_unsigned(1014, 12), 656 => to_unsigned(2356, 12), 657 => to_unsigned(3172, 12), 658 => to_unsigned(1746, 12), 659 => to_unsigned(1725, 12), 660 => to_unsigned(1834, 12), 661 => to_unsigned(2905, 12), 662 => to_unsigned(3968, 12), 663 => to_unsigned(513, 12), 664 => to_unsigned(3100, 12), 665 => to_unsigned(2835, 12), 666 => to_unsigned(3231, 12), 667 => to_unsigned(1556, 12), 668 => to_unsigned(3827, 12), 669 => to_unsigned(2732, 12), 670 => to_unsigned(1803, 12), 671 => to_unsigned(3987, 12), 672 => to_unsigned(2216, 12), 673 => to_unsigned(4063, 12), 674 => to_unsigned(4025, 12), 675 => to_unsigned(3465, 12), 676 => to_unsigned(249, 12), 677 => to_unsigned(847, 12), 678 => to_unsigned(1953, 12), 679 => to_unsigned(2420, 12), 680 => to_unsigned(660, 12), 681 => to_unsigned(776, 12), 682 => to_unsigned(2501, 12), 683 => to_unsigned(1231, 12), 684 => to_unsigned(1746, 12), 685 => to_unsigned(777, 12), 686 => to_unsigned(3772, 12), 687 => to_unsigned(2054, 12), 688 => to_unsigned(2483, 12), 689 => to_unsigned(3202, 12), 690 => to_unsigned(1805, 12), 691 => to_unsigned(2582, 12), 692 => to_unsigned(895, 12), 693 => to_unsigned(950, 12), 694 => to_unsigned(2946, 12), 695 => to_unsigned(3639, 12), 696 => to_unsigned(377, 12), 697 => to_unsigned(1368, 12), 698 => to_unsigned(2351, 12), 699 => to_unsigned(2225, 12), 700 => to_unsigned(476, 12), 701 => to_unsigned(1833, 12), 702 => to_unsigned(2473, 12), 703 => to_unsigned(1462, 12), 704 => to_unsigned(28, 12), 705 => to_unsigned(3540, 12), 706 => to_unsigned(3928, 12), 707 => to_unsigned(2247, 12), 708 => to_unsigned(1293, 12), 709 => to_unsigned(2925, 12), 710 => to_unsigned(2290, 12), 711 => to_unsigned(1135, 12), 712 => to_unsigned(3642, 12), 713 => to_unsigned(243, 12), 714 => to_unsigned(3061, 12), 715 => to_unsigned(342, 12), 716 => to_unsigned(2670, 12), 717 => to_unsigned(2774, 12), 718 => to_unsigned(3877, 12), 719 => to_unsigned(2257, 12), 720 => to_unsigned(3327, 12), 721 => to_unsigned(149, 12), 722 => to_unsigned(532, 12), 723 => to_unsigned(2998, 12), 724 => to_unsigned(3138, 12), 725 => to_unsigned(1645, 12), 726 => to_unsigned(2381, 12), 727 => to_unsigned(3119, 12), 728 => to_unsigned(2826, 12), 729 => to_unsigned(770, 12), 730 => to_unsigned(1787, 12), 731 => to_unsigned(3718, 12), 732 => to_unsigned(2383, 12), 733 => to_unsigned(325, 12), 734 => to_unsigned(3216, 12), 735 => to_unsigned(2766, 12), 736 => to_unsigned(2602, 12), 737 => to_unsigned(1819, 12), 738 => to_unsigned(3976, 12), 739 => to_unsigned(2157, 12), 740 => to_unsigned(2988, 12), 741 => to_unsigned(1093, 12), 742 => to_unsigned(1980, 12), 743 => to_unsigned(1353, 12), 744 => to_unsigned(2431, 12), 745 => to_unsigned(2355, 12), 746 => to_unsigned(931, 12), 747 => to_unsigned(1736, 12), 748 => to_unsigned(2597, 12), 749 => to_unsigned(690, 12), 750 => to_unsigned(3460, 12), 751 => to_unsigned(3063, 12), 752 => to_unsigned(1732, 12), 753 => to_unsigned(2919, 12), 754 => to_unsigned(3005, 12), 755 => to_unsigned(557, 12), 756 => to_unsigned(302, 12), 757 => to_unsigned(820, 12), 758 => to_unsigned(2232, 12), 759 => to_unsigned(587, 12), 760 => to_unsigned(660, 12), 761 => to_unsigned(3464, 12), 762 => to_unsigned(3449, 12), 763 => to_unsigned(2784, 12), 764 => to_unsigned(2466, 12), 765 => to_unsigned(3947, 12), 766 => to_unsigned(1637, 12), 767 => to_unsigned(1556, 12), 768 => to_unsigned(51, 12), 769 => to_unsigned(2899, 12), 770 => to_unsigned(1087, 12), 771 => to_unsigned(3716, 12), 772 => to_unsigned(2090, 12), 773 => to_unsigned(3373, 12), 774 => to_unsigned(2977, 12), 775 => to_unsigned(2673, 12), 776 => to_unsigned(975, 12), 777 => to_unsigned(1265, 12), 778 => to_unsigned(996, 12), 779 => to_unsigned(823, 12), 780 => to_unsigned(3160, 12), 781 => to_unsigned(36, 12), 782 => to_unsigned(3287, 12), 783 => to_unsigned(2400, 12), 784 => to_unsigned(55, 12), 785 => to_unsigned(1005, 12), 786 => to_unsigned(3548, 12), 787 => to_unsigned(3202, 12), 788 => to_unsigned(134, 12), 789 => to_unsigned(3138, 12), 790 => to_unsigned(555, 12), 791 => to_unsigned(919, 12), 792 => to_unsigned(1743, 12), 793 => to_unsigned(1710, 12), 794 => to_unsigned(3035, 12), 795 => to_unsigned(1518, 12), 796 => to_unsigned(1331, 12), 797 => to_unsigned(963, 12), 798 => to_unsigned(2475, 12), 799 => to_unsigned(2013, 12), 800 => to_unsigned(620, 12), 801 => to_unsigned(1142, 12), 802 => to_unsigned(2793, 12), 803 => to_unsigned(1597, 12), 804 => to_unsigned(2178, 12), 805 => to_unsigned(2902, 12), 806 => to_unsigned(320, 12), 807 => to_unsigned(948, 12), 808 => to_unsigned(447, 12), 809 => to_unsigned(3255, 12), 810 => to_unsigned(3385, 12), 811 => to_unsigned(1196, 12), 812 => to_unsigned(241, 12), 813 => to_unsigned(4082, 12), 814 => to_unsigned(1856, 12), 815 => to_unsigned(993, 12), 816 => to_unsigned(1487, 12), 817 => to_unsigned(314, 12), 818 => to_unsigned(2694, 12), 819 => to_unsigned(3570, 12), 820 => to_unsigned(3521, 12), 821 => to_unsigned(0, 12), 822 => to_unsigned(85, 12), 823 => to_unsigned(3440, 12), 824 => to_unsigned(3857, 12), 825 => to_unsigned(1018, 12), 826 => to_unsigned(2822, 12), 827 => to_unsigned(62, 12), 828 => to_unsigned(3256, 12), 829 => to_unsigned(2636, 12), 830 => to_unsigned(3081, 12), 831 => to_unsigned(3086, 12), 832 => to_unsigned(4038, 12), 833 => to_unsigned(506, 12), 834 => to_unsigned(1650, 12), 835 => to_unsigned(2527, 12), 836 => to_unsigned(1729, 12), 837 => to_unsigned(1502, 12), 838 => to_unsigned(820, 12), 839 => to_unsigned(2400, 12), 840 => to_unsigned(2200, 12), 841 => to_unsigned(1763, 12), 842 => to_unsigned(3019, 12), 843 => to_unsigned(1300, 12), 844 => to_unsigned(3650, 12), 845 => to_unsigned(2290, 12), 846 => to_unsigned(1720, 12), 847 => to_unsigned(2892, 12), 848 => to_unsigned(2288, 12), 849 => to_unsigned(3857, 12), 850 => to_unsigned(20, 12), 851 => to_unsigned(1135, 12), 852 => to_unsigned(1248, 12), 853 => to_unsigned(1601, 12), 854 => to_unsigned(3137, 12), 855 => to_unsigned(3682, 12), 856 => to_unsigned(711, 12), 857 => to_unsigned(3378, 12), 858 => to_unsigned(3517, 12), 859 => to_unsigned(407, 12), 860 => to_unsigned(2407, 12), 861 => to_unsigned(2369, 12), 862 => to_unsigned(1384, 12), 863 => to_unsigned(1713, 12), 864 => to_unsigned(1878, 12), 865 => to_unsigned(653, 12), 866 => to_unsigned(3112, 12), 867 => to_unsigned(3978, 12), 868 => to_unsigned(3173, 12), 869 => to_unsigned(2242, 12), 870 => to_unsigned(815, 12), 871 => to_unsigned(2661, 12), 872 => to_unsigned(834, 12), 873 => to_unsigned(1311, 12), 874 => to_unsigned(2096, 12), 875 => to_unsigned(675, 12), 876 => to_unsigned(2715, 12), 877 => to_unsigned(1241, 12), 878 => to_unsigned(1290, 12), 879 => to_unsigned(1382, 12), 880 => to_unsigned(3814, 12), 881 => to_unsigned(2602, 12), 882 => to_unsigned(2520, 12), 883 => to_unsigned(1310, 12), 884 => to_unsigned(121, 12), 885 => to_unsigned(1338, 12), 886 => to_unsigned(1802, 12), 887 => to_unsigned(1069, 12), 888 => to_unsigned(874, 12), 889 => to_unsigned(2042, 12), 890 => to_unsigned(1411, 12), 891 => to_unsigned(1926, 12), 892 => to_unsigned(3385, 12), 893 => to_unsigned(3081, 12), 894 => to_unsigned(299, 12), 895 => to_unsigned(3457, 12), 896 => to_unsigned(1609, 12), 897 => to_unsigned(2609, 12), 898 => to_unsigned(3929, 12), 899 => to_unsigned(1488, 12), 900 => to_unsigned(3847, 12), 901 => to_unsigned(2280, 12), 902 => to_unsigned(235, 12), 903 => to_unsigned(1921, 12), 904 => to_unsigned(59, 12), 905 => to_unsigned(3648, 12), 906 => to_unsigned(1367, 12), 907 => to_unsigned(115, 12), 908 => to_unsigned(47, 12), 909 => to_unsigned(3246, 12), 910 => to_unsigned(2074, 12), 911 => to_unsigned(2610, 12), 912 => to_unsigned(1330, 12), 913 => to_unsigned(2260, 12), 914 => to_unsigned(3115, 12), 915 => to_unsigned(408, 12), 916 => to_unsigned(682, 12), 917 => to_unsigned(1222, 12), 918 => to_unsigned(2644, 12), 919 => to_unsigned(2095, 12), 920 => to_unsigned(1393, 12), 921 => to_unsigned(1145, 12), 922 => to_unsigned(3947, 12), 923 => to_unsigned(3556, 12), 924 => to_unsigned(389, 12), 925 => to_unsigned(1262, 12), 926 => to_unsigned(3380, 12), 927 => to_unsigned(327, 12), 928 => to_unsigned(3100, 12), 929 => to_unsigned(54, 12), 930 => to_unsigned(3976, 12), 931 => to_unsigned(2671, 12), 932 => to_unsigned(3815, 12), 933 => to_unsigned(3574, 12), 934 => to_unsigned(1824, 12), 935 => to_unsigned(526, 12), 936 => to_unsigned(2769, 12), 937 => to_unsigned(1436, 12), 938 => to_unsigned(2885, 12), 939 => to_unsigned(2550, 12), 940 => to_unsigned(861, 12), 941 => to_unsigned(1581, 12), 942 => to_unsigned(3245, 12), 943 => to_unsigned(1640, 12), 944 => to_unsigned(3603, 12), 945 => to_unsigned(4046, 12), 946 => to_unsigned(2093, 12), 947 => to_unsigned(1112, 12), 948 => to_unsigned(2503, 12), 949 => to_unsigned(1914, 12), 950 => to_unsigned(760, 12), 951 => to_unsigned(1135, 12), 952 => to_unsigned(1102, 12), 953 => to_unsigned(1882, 12), 954 => to_unsigned(1439, 12), 955 => to_unsigned(2445, 12), 956 => to_unsigned(478, 12), 957 => to_unsigned(646, 12), 958 => to_unsigned(1340, 12), 959 => to_unsigned(437, 12), 960 => to_unsigned(2685, 12), 961 => to_unsigned(3042, 12), 962 => to_unsigned(4070, 12), 963 => to_unsigned(2284, 12), 964 => to_unsigned(642, 12), 965 => to_unsigned(1573, 12), 966 => to_unsigned(1767, 12), 967 => to_unsigned(1409, 12), 968 => to_unsigned(2938, 12), 969 => to_unsigned(385, 12), 970 => to_unsigned(3862, 12), 971 => to_unsigned(3888, 12), 972 => to_unsigned(3754, 12), 973 => to_unsigned(891, 12), 974 => to_unsigned(494, 12), 975 => to_unsigned(878, 12), 976 => to_unsigned(2803, 12), 977 => to_unsigned(1145, 12), 978 => to_unsigned(522, 12), 979 => to_unsigned(2510, 12), 980 => to_unsigned(2292, 12), 981 => to_unsigned(1557, 12), 982 => to_unsigned(4021, 12), 983 => to_unsigned(3751, 12), 984 => to_unsigned(987, 12), 985 => to_unsigned(2903, 12), 986 => to_unsigned(2750, 12), 987 => to_unsigned(116, 12), 988 => to_unsigned(1598, 12), 989 => to_unsigned(2560, 12), 990 => to_unsigned(1381, 12), 991 => to_unsigned(263, 12), 992 => to_unsigned(779, 12), 993 => to_unsigned(503, 12), 994 => to_unsigned(879, 12), 995 => to_unsigned(1411, 12), 996 => to_unsigned(1363, 12), 997 => to_unsigned(3488, 12), 998 => to_unsigned(3693, 12), 999 => to_unsigned(3048, 12), 1000 => to_unsigned(4080, 12), 1001 => to_unsigned(51, 12), 1002 => to_unsigned(1351, 12), 1003 => to_unsigned(2919, 12), 1004 => to_unsigned(2440, 12), 1005 => to_unsigned(3338, 12), 1006 => to_unsigned(1877, 12), 1007 => to_unsigned(2788, 12), 1008 => to_unsigned(3789, 12), 1009 => to_unsigned(3038, 12), 1010 => to_unsigned(3933, 12), 1011 => to_unsigned(1904, 12), 1012 => to_unsigned(2842, 12), 1013 => to_unsigned(1150, 12), 1014 => to_unsigned(2568, 12), 1015 => to_unsigned(979, 12), 1016 => to_unsigned(4030, 12), 1017 => to_unsigned(3862, 12), 1018 => to_unsigned(559, 12), 1019 => to_unsigned(298, 12), 1020 => to_unsigned(1514, 12), 1021 => to_unsigned(3082, 12), 1022 => to_unsigned(1562, 12), 1023 => to_unsigned(538, 12), 1024 => to_unsigned(1049, 12), 1025 => to_unsigned(1732, 12), 1026 => to_unsigned(1509, 12), 1027 => to_unsigned(422, 12), 1028 => to_unsigned(1810, 12), 1029 => to_unsigned(370, 12), 1030 => to_unsigned(991, 12), 1031 => to_unsigned(1660, 12), 1032 => to_unsigned(3000, 12), 1033 => to_unsigned(2127, 12), 1034 => to_unsigned(3244, 12), 1035 => to_unsigned(2798, 12), 1036 => to_unsigned(3034, 12), 1037 => to_unsigned(699, 12), 1038 => to_unsigned(514, 12), 1039 => to_unsigned(25, 12), 1040 => to_unsigned(3489, 12), 1041 => to_unsigned(3585, 12), 1042 => to_unsigned(3509, 12), 1043 => to_unsigned(2956, 12), 1044 => to_unsigned(3777, 12), 1045 => to_unsigned(2173, 12), 1046 => to_unsigned(331, 12), 1047 => to_unsigned(257, 12), 1048 => to_unsigned(1347, 12), 1049 => to_unsigned(2194, 12), 1050 => to_unsigned(1055, 12), 1051 => to_unsigned(1655, 12), 1052 => to_unsigned(3210, 12), 1053 => to_unsigned(639, 12), 1054 => to_unsigned(1217, 12), 1055 => to_unsigned(63, 12), 1056 => to_unsigned(512, 12), 1057 => to_unsigned(140, 12), 1058 => to_unsigned(340, 12), 1059 => to_unsigned(1306, 12), 1060 => to_unsigned(2394, 12), 1061 => to_unsigned(2369, 12), 1062 => to_unsigned(3767, 12), 1063 => to_unsigned(184, 12), 1064 => to_unsigned(118, 12), 1065 => to_unsigned(2724, 12), 1066 => to_unsigned(3836, 12), 1067 => to_unsigned(1447, 12), 1068 => to_unsigned(2867, 12), 1069 => to_unsigned(2358, 12), 1070 => to_unsigned(2832, 12), 1071 => to_unsigned(1468, 12), 1072 => to_unsigned(693, 12), 1073 => to_unsigned(993, 12), 1074 => to_unsigned(3997, 12), 1075 => to_unsigned(2622, 12), 1076 => to_unsigned(2033, 12), 1077 => to_unsigned(2660, 12), 1078 => to_unsigned(3412, 12), 1079 => to_unsigned(1534, 12), 1080 => to_unsigned(425, 12), 1081 => to_unsigned(3930, 12), 1082 => to_unsigned(2375, 12), 1083 => to_unsigned(2608, 12), 1084 => to_unsigned(1913, 12), 1085 => to_unsigned(1821, 12), 1086 => to_unsigned(814, 12), 1087 => to_unsigned(4040, 12), 1088 => to_unsigned(1949, 12), 1089 => to_unsigned(2639, 12), 1090 => to_unsigned(3132, 12), 1091 => to_unsigned(3280, 12), 1092 => to_unsigned(734, 12), 1093 => to_unsigned(1289, 12), 1094 => to_unsigned(1117, 12), 1095 => to_unsigned(2459, 12), 1096 => to_unsigned(3167, 12), 1097 => to_unsigned(1029, 12), 1098 => to_unsigned(3029, 12), 1099 => to_unsigned(1164, 12), 1100 => to_unsigned(2640, 12), 1101 => to_unsigned(2316, 12), 1102 => to_unsigned(3256, 12), 1103 => to_unsigned(3961, 12), 1104 => to_unsigned(2799, 12), 1105 => to_unsigned(284, 12), 1106 => to_unsigned(329, 12), 1107 => to_unsigned(3225, 12), 1108 => to_unsigned(1896, 12), 1109 => to_unsigned(2596, 12), 1110 => to_unsigned(2724, 12), 1111 => to_unsigned(3620, 12), 1112 => to_unsigned(2862, 12), 1113 => to_unsigned(811, 12), 1114 => to_unsigned(3132, 12), 1115 => to_unsigned(3061, 12), 1116 => to_unsigned(3793, 12), 1117 => to_unsigned(2072, 12), 1118 => to_unsigned(1879, 12), 1119 => to_unsigned(3828, 12), 1120 => to_unsigned(659, 12), 1121 => to_unsigned(2510, 12), 1122 => to_unsigned(923, 12), 1123 => to_unsigned(3927, 12), 1124 => to_unsigned(270, 12), 1125 => to_unsigned(2217, 12), 1126 => to_unsigned(2283, 12), 1127 => to_unsigned(3472, 12), 1128 => to_unsigned(3421, 12), 1129 => to_unsigned(2076, 12), 1130 => to_unsigned(2799, 12), 1131 => to_unsigned(332, 12), 1132 => to_unsigned(576, 12), 1133 => to_unsigned(4075, 12), 1134 => to_unsigned(551, 12), 1135 => to_unsigned(1883, 12), 1136 => to_unsigned(3156, 12), 1137 => to_unsigned(3667, 12), 1138 => to_unsigned(392, 12), 1139 => to_unsigned(3781, 12), 1140 => to_unsigned(1031, 12), 1141 => to_unsigned(3550, 12), 1142 => to_unsigned(3458, 12), 1143 => to_unsigned(3299, 12), 1144 => to_unsigned(2632, 12), 1145 => to_unsigned(2192, 12), 1146 => to_unsigned(3728, 12), 1147 => to_unsigned(2151, 12), 1148 => to_unsigned(3079, 12), 1149 => to_unsigned(3816, 12), 1150 => to_unsigned(3691, 12), 1151 => to_unsigned(1210, 12), 1152 => to_unsigned(1600, 12), 1153 => to_unsigned(726, 12), 1154 => to_unsigned(3684, 12), 1155 => to_unsigned(305, 12), 1156 => to_unsigned(2676, 12), 1157 => to_unsigned(2033, 12), 1158 => to_unsigned(2725, 12), 1159 => to_unsigned(3129, 12), 1160 => to_unsigned(57, 12), 1161 => to_unsigned(1017, 12), 1162 => to_unsigned(2893, 12), 1163 => to_unsigned(2938, 12), 1164 => to_unsigned(554, 12), 1165 => to_unsigned(1863, 12), 1166 => to_unsigned(1977, 12), 1167 => to_unsigned(2693, 12), 1168 => to_unsigned(2085, 12), 1169 => to_unsigned(1963, 12), 1170 => to_unsigned(3085, 12), 1171 => to_unsigned(3198, 12), 1172 => to_unsigned(1059, 12), 1173 => to_unsigned(2455, 12), 1174 => to_unsigned(570, 12), 1175 => to_unsigned(782, 12), 1176 => to_unsigned(2345, 12), 1177 => to_unsigned(3775, 12), 1178 => to_unsigned(2815, 12), 1179 => to_unsigned(3013, 12), 1180 => to_unsigned(405, 12), 1181 => to_unsigned(1133, 12), 1182 => to_unsigned(922, 12), 1183 => to_unsigned(2522, 12), 1184 => to_unsigned(2669, 12), 1185 => to_unsigned(2058, 12), 1186 => to_unsigned(1452, 12), 1187 => to_unsigned(871, 12), 1188 => to_unsigned(1433, 12), 1189 => to_unsigned(7, 12), 1190 => to_unsigned(2111, 12), 1191 => to_unsigned(954, 12), 1192 => to_unsigned(3890, 12), 1193 => to_unsigned(853, 12), 1194 => to_unsigned(938, 12), 1195 => to_unsigned(3529, 12), 1196 => to_unsigned(1388, 12), 1197 => to_unsigned(3676, 12), 1198 => to_unsigned(3725, 12), 1199 => to_unsigned(2553, 12), 1200 => to_unsigned(1855, 12), 1201 => to_unsigned(2799, 12), 1202 => to_unsigned(3303, 12), 1203 => to_unsigned(1904, 12), 1204 => to_unsigned(2444, 12), 1205 => to_unsigned(591, 12), 1206 => to_unsigned(3131, 12), 1207 => to_unsigned(2468, 12), 1208 => to_unsigned(1085, 12), 1209 => to_unsigned(73, 12), 1210 => to_unsigned(1734, 12), 1211 => to_unsigned(3372, 12), 1212 => to_unsigned(3508, 12), 1213 => to_unsigned(1493, 12), 1214 => to_unsigned(551, 12), 1215 => to_unsigned(790, 12), 1216 => to_unsigned(2252, 12), 1217 => to_unsigned(420, 12), 1218 => to_unsigned(730, 12), 1219 => to_unsigned(1955, 12), 1220 => to_unsigned(3059, 12), 1221 => to_unsigned(984, 12), 1222 => to_unsigned(136, 12), 1223 => to_unsigned(1537, 12), 1224 => to_unsigned(1711, 12), 1225 => to_unsigned(407, 12), 1226 => to_unsigned(1454, 12), 1227 => to_unsigned(1004, 12), 1228 => to_unsigned(3102, 12), 1229 => to_unsigned(3974, 12), 1230 => to_unsigned(2442, 12), 1231 => to_unsigned(325, 12), 1232 => to_unsigned(2005, 12), 1233 => to_unsigned(2219, 12), 1234 => to_unsigned(2884, 12), 1235 => to_unsigned(1345, 12), 1236 => to_unsigned(2807, 12), 1237 => to_unsigned(3496, 12), 1238 => to_unsigned(430, 12), 1239 => to_unsigned(4028, 12), 1240 => to_unsigned(4018, 12), 1241 => to_unsigned(1100, 12), 1242 => to_unsigned(1778, 12), 1243 => to_unsigned(707, 12), 1244 => to_unsigned(630, 12), 1245 => to_unsigned(3028, 12), 1246 => to_unsigned(2408, 12), 1247 => to_unsigned(2743, 12), 1248 => to_unsigned(526, 12), 1249 => to_unsigned(3531, 12), 1250 => to_unsigned(3912, 12), 1251 => to_unsigned(1037, 12), 1252 => to_unsigned(226, 12), 1253 => to_unsigned(3747, 12), 1254 => to_unsigned(3846, 12), 1255 => to_unsigned(1657, 12), 1256 => to_unsigned(328, 12), 1257 => to_unsigned(1870, 12), 1258 => to_unsigned(3168, 12), 1259 => to_unsigned(2929, 12), 1260 => to_unsigned(721, 12), 1261 => to_unsigned(4001, 12), 1262 => to_unsigned(3443, 12), 1263 => to_unsigned(1018, 12), 1264 => to_unsigned(1873, 12), 1265 => to_unsigned(2908, 12), 1266 => to_unsigned(1234, 12), 1267 => to_unsigned(20, 12), 1268 => to_unsigned(1000, 12), 1269 => to_unsigned(1029, 12), 1270 => to_unsigned(3673, 12), 1271 => to_unsigned(1886, 12), 1272 => to_unsigned(3105, 12), 1273 => to_unsigned(994, 12), 1274 => to_unsigned(1454, 12), 1275 => to_unsigned(799, 12), 1276 => to_unsigned(3341, 12), 1277 => to_unsigned(3663, 12), 1278 => to_unsigned(3769, 12), 1279 => to_unsigned(324, 12), 1280 => to_unsigned(3765, 12), 1281 => to_unsigned(2557, 12), 1282 => to_unsigned(1914, 12), 1283 => to_unsigned(3033, 12), 1284 => to_unsigned(3102, 12), 1285 => to_unsigned(2639, 12), 1286 => to_unsigned(2686, 12), 1287 => to_unsigned(1901, 12), 1288 => to_unsigned(2970, 12), 1289 => to_unsigned(1268, 12), 1290 => to_unsigned(1230, 12), 1291 => to_unsigned(3053, 12), 1292 => to_unsigned(1981, 12), 1293 => to_unsigned(68, 12), 1294 => to_unsigned(1886, 12), 1295 => to_unsigned(407, 12), 1296 => to_unsigned(1646, 12), 1297 => to_unsigned(3636, 12), 1298 => to_unsigned(622, 12), 1299 => to_unsigned(2592, 12), 1300 => to_unsigned(2548, 12), 1301 => to_unsigned(1722, 12), 1302 => to_unsigned(986, 12), 1303 => to_unsigned(1607, 12), 1304 => to_unsigned(716, 12), 1305 => to_unsigned(1072, 12), 1306 => to_unsigned(2531, 12), 1307 => to_unsigned(1383, 12), 1308 => to_unsigned(2700, 12), 1309 => to_unsigned(1509, 12), 1310 => to_unsigned(2273, 12), 1311 => to_unsigned(3409, 12), 1312 => to_unsigned(3502, 12), 1313 => to_unsigned(1544, 12), 1314 => to_unsigned(3123, 12), 1315 => to_unsigned(3269, 12), 1316 => to_unsigned(3836, 12), 1317 => to_unsigned(797, 12), 1318 => to_unsigned(851, 12), 1319 => to_unsigned(336, 12), 1320 => to_unsigned(11, 12), 1321 => to_unsigned(2788, 12), 1322 => to_unsigned(1173, 12), 1323 => to_unsigned(2666, 12), 1324 => to_unsigned(3421, 12), 1325 => to_unsigned(3720, 12), 1326 => to_unsigned(2504, 12), 1327 => to_unsigned(4021, 12), 1328 => to_unsigned(3655, 12), 1329 => to_unsigned(329, 12), 1330 => to_unsigned(3502, 12), 1331 => to_unsigned(1137, 12), 1332 => to_unsigned(1160, 12), 1333 => to_unsigned(3365, 12), 1334 => to_unsigned(492, 12), 1335 => to_unsigned(3921, 12), 1336 => to_unsigned(2048, 12), 1337 => to_unsigned(1501, 12), 1338 => to_unsigned(239, 12), 1339 => to_unsigned(1145, 12), 1340 => to_unsigned(241, 12), 1341 => to_unsigned(1451, 12), 1342 => to_unsigned(1955, 12), 1343 => to_unsigned(2043, 12), 1344 => to_unsigned(2905, 12), 1345 => to_unsigned(663, 12), 1346 => to_unsigned(752, 12), 1347 => to_unsigned(1722, 12), 1348 => to_unsigned(159, 12), 1349 => to_unsigned(3326, 12), 1350 => to_unsigned(838, 12), 1351 => to_unsigned(1692, 12), 1352 => to_unsigned(2173, 12), 1353 => to_unsigned(1604, 12), 1354 => to_unsigned(1204, 12), 1355 => to_unsigned(2763, 12), 1356 => to_unsigned(3281, 12), 1357 => to_unsigned(1921, 12), 1358 => to_unsigned(2631, 12), 1359 => to_unsigned(1462, 12), 1360 => to_unsigned(2728, 12), 1361 => to_unsigned(1367, 12), 1362 => to_unsigned(790, 12), 1363 => to_unsigned(664, 12), 1364 => to_unsigned(2019, 12), 1365 => to_unsigned(1334, 12), 1366 => to_unsigned(1255, 12), 1367 => to_unsigned(1411, 12), 1368 => to_unsigned(498, 12), 1369 => to_unsigned(2227, 12), 1370 => to_unsigned(2021, 12), 1371 => to_unsigned(3258, 12), 1372 => to_unsigned(951, 12), 1373 => to_unsigned(1591, 12), 1374 => to_unsigned(1248, 12), 1375 => to_unsigned(3711, 12), 1376 => to_unsigned(3424, 12), 1377 => to_unsigned(3394, 12), 1378 => to_unsigned(1820, 12), 1379 => to_unsigned(1004, 12), 1380 => to_unsigned(3147, 12), 1381 => to_unsigned(509, 12), 1382 => to_unsigned(714, 12), 1383 => to_unsigned(3247, 12), 1384 => to_unsigned(3630, 12), 1385 => to_unsigned(55, 12), 1386 => to_unsigned(1917, 12), 1387 => to_unsigned(1875, 12), 1388 => to_unsigned(1016, 12), 1389 => to_unsigned(3212, 12), 1390 => to_unsigned(471, 12), 1391 => to_unsigned(2353, 12), 1392 => to_unsigned(3369, 12), 1393 => to_unsigned(2609, 12), 1394 => to_unsigned(3395, 12), 1395 => to_unsigned(3442, 12), 1396 => to_unsigned(3171, 12), 1397 => to_unsigned(3895, 12), 1398 => to_unsigned(2103, 12), 1399 => to_unsigned(1111, 12), 1400 => to_unsigned(1529, 12), 1401 => to_unsigned(1218, 12), 1402 => to_unsigned(2367, 12), 1403 => to_unsigned(1394, 12), 1404 => to_unsigned(213, 12), 1405 => to_unsigned(386, 12), 1406 => to_unsigned(3611, 12), 1407 => to_unsigned(2550, 12), 1408 => to_unsigned(3133, 12), 1409 => to_unsigned(2563, 12), 1410 => to_unsigned(197, 12), 1411 => to_unsigned(3650, 12), 1412 => to_unsigned(846, 12), 1413 => to_unsigned(1551, 12), 1414 => to_unsigned(3488, 12), 1415 => to_unsigned(2828, 12), 1416 => to_unsigned(944, 12), 1417 => to_unsigned(60, 12), 1418 => to_unsigned(4026, 12), 1419 => to_unsigned(520, 12), 1420 => to_unsigned(3015, 12), 1421 => to_unsigned(2731, 12), 1422 => to_unsigned(894, 12), 1423 => to_unsigned(4083, 12), 1424 => to_unsigned(2402, 12), 1425 => to_unsigned(205, 12), 1426 => to_unsigned(2795, 12), 1427 => to_unsigned(3896, 12), 1428 => to_unsigned(3571, 12), 1429 => to_unsigned(3660, 12), 1430 => to_unsigned(1717, 12), 1431 => to_unsigned(2853, 12), 1432 => to_unsigned(1889, 12), 1433 => to_unsigned(3183, 12), 1434 => to_unsigned(2936, 12), 1435 => to_unsigned(2536, 12), 1436 => to_unsigned(476, 12), 1437 => to_unsigned(3660, 12), 1438 => to_unsigned(2158, 12), 1439 => to_unsigned(497, 12), 1440 => to_unsigned(3767, 12), 1441 => to_unsigned(33, 12), 1442 => to_unsigned(49, 12), 1443 => to_unsigned(2019, 12), 1444 => to_unsigned(2913, 12), 1445 => to_unsigned(3932, 12), 1446 => to_unsigned(1026, 12), 1447 => to_unsigned(2974, 12), 1448 => to_unsigned(4015, 12), 1449 => to_unsigned(132, 12), 1450 => to_unsigned(2519, 12), 1451 => to_unsigned(2958, 12), 1452 => to_unsigned(2212, 12), 1453 => to_unsigned(1860, 12), 1454 => to_unsigned(229, 12), 1455 => to_unsigned(3832, 12), 1456 => to_unsigned(1490, 12), 1457 => to_unsigned(2131, 12), 1458 => to_unsigned(382, 12), 1459 => to_unsigned(3635, 12), 1460 => to_unsigned(230, 12), 1461 => to_unsigned(1617, 12), 1462 => to_unsigned(2538, 12), 1463 => to_unsigned(3827, 12), 1464 => to_unsigned(2456, 12), 1465 => to_unsigned(1334, 12), 1466 => to_unsigned(1153, 12), 1467 => to_unsigned(1126, 12), 1468 => to_unsigned(3006, 12), 1469 => to_unsigned(1845, 12), 1470 => to_unsigned(160, 12), 1471 => to_unsigned(4034, 12), 1472 => to_unsigned(805, 12), 1473 => to_unsigned(1353, 12), 1474 => to_unsigned(3855, 12), 1475 => to_unsigned(1029, 12), 1476 => to_unsigned(1414, 12), 1477 => to_unsigned(2076, 12), 1478 => to_unsigned(2851, 12), 1479 => to_unsigned(292, 12), 1480 => to_unsigned(3517, 12), 1481 => to_unsigned(712, 12), 1482 => to_unsigned(1207, 12), 1483 => to_unsigned(3378, 12), 1484 => to_unsigned(2881, 12), 1485 => to_unsigned(3398, 12), 1486 => to_unsigned(2383, 12), 1487 => to_unsigned(3519, 12), 1488 => to_unsigned(775, 12), 1489 => to_unsigned(2741, 12), 1490 => to_unsigned(2057, 12), 1491 => to_unsigned(752, 12), 1492 => to_unsigned(3306, 12), 1493 => to_unsigned(592, 12), 1494 => to_unsigned(1387, 12), 1495 => to_unsigned(2002, 12), 1496 => to_unsigned(1291, 12), 1497 => to_unsigned(1621, 12), 1498 => to_unsigned(3040, 12), 1499 => to_unsigned(2293, 12), 1500 => to_unsigned(3345, 12), 1501 => to_unsigned(1289, 12), 1502 => to_unsigned(2577, 12), 1503 => to_unsigned(3835, 12), 1504 => to_unsigned(1544, 12), 1505 => to_unsigned(2276, 12), 1506 => to_unsigned(4011, 12), 1507 => to_unsigned(283, 12), 1508 => to_unsigned(849, 12), 1509 => to_unsigned(2601, 12), 1510 => to_unsigned(1857, 12), 1511 => to_unsigned(2413, 12), 1512 => to_unsigned(3420, 12), 1513 => to_unsigned(726, 12), 1514 => to_unsigned(916, 12), 1515 => to_unsigned(3427, 12), 1516 => to_unsigned(169, 12), 1517 => to_unsigned(401, 12), 1518 => to_unsigned(3051, 12), 1519 => to_unsigned(3337, 12), 1520 => to_unsigned(1695, 12), 1521 => to_unsigned(752, 12), 1522 => to_unsigned(1056, 12), 1523 => to_unsigned(2463, 12), 1524 => to_unsigned(139, 12), 1525 => to_unsigned(543, 12), 1526 => to_unsigned(1782, 12), 1527 => to_unsigned(3471, 12), 1528 => to_unsigned(952, 12), 1529 => to_unsigned(339, 12), 1530 => to_unsigned(3741, 12), 1531 => to_unsigned(3731, 12), 1532 => to_unsigned(793, 12), 1533 => to_unsigned(171, 12), 1534 => to_unsigned(1621, 12), 1535 => to_unsigned(858, 12), 1536 => to_unsigned(3392, 12), 1537 => to_unsigned(337, 12), 1538 => to_unsigned(128, 12), 1539 => to_unsigned(2537, 12), 1540 => to_unsigned(3193, 12), 1541 => to_unsigned(1407, 12), 1542 => to_unsigned(4041, 12), 1543 => to_unsigned(3190, 12), 1544 => to_unsigned(2217, 12), 1545 => to_unsigned(1550, 12), 1546 => to_unsigned(171, 12), 1547 => to_unsigned(2888, 12), 1548 => to_unsigned(2276, 12), 1549 => to_unsigned(1259, 12), 1550 => to_unsigned(2038, 12), 1551 => to_unsigned(1636, 12), 1552 => to_unsigned(4012, 12), 1553 => to_unsigned(971, 12), 1554 => to_unsigned(685, 12), 1555 => to_unsigned(1747, 12), 1556 => to_unsigned(789, 12), 1557 => to_unsigned(140, 12), 1558 => to_unsigned(1154, 12), 1559 => to_unsigned(1015, 12), 1560 => to_unsigned(1282, 12), 1561 => to_unsigned(2948, 12), 1562 => to_unsigned(201, 12), 1563 => to_unsigned(2156, 12), 1564 => to_unsigned(1068, 12), 1565 => to_unsigned(1556, 12), 1566 => to_unsigned(1236, 12), 1567 => to_unsigned(1983, 12), 1568 => to_unsigned(3132, 12), 1569 => to_unsigned(1710, 12), 1570 => to_unsigned(3285, 12), 1571 => to_unsigned(3746, 12), 1572 => to_unsigned(1719, 12), 1573 => to_unsigned(1112, 12), 1574 => to_unsigned(2045, 12), 1575 => to_unsigned(1702, 12), 1576 => to_unsigned(1072, 12), 1577 => to_unsigned(2976, 12), 1578 => to_unsigned(228, 12), 1579 => to_unsigned(422, 12), 1580 => to_unsigned(148, 12), 1581 => to_unsigned(1256, 12), 1582 => to_unsigned(275, 12), 1583 => to_unsigned(3086, 12), 1584 => to_unsigned(1217, 12), 1585 => to_unsigned(3070, 12), 1586 => to_unsigned(410, 12), 1587 => to_unsigned(1521, 12), 1588 => to_unsigned(777, 12), 1589 => to_unsigned(2796, 12), 1590 => to_unsigned(1000, 12), 1591 => to_unsigned(2919, 12), 1592 => to_unsigned(716, 12), 1593 => to_unsigned(3444, 12), 1594 => to_unsigned(1208, 12), 1595 => to_unsigned(796, 12), 1596 => to_unsigned(940, 12), 1597 => to_unsigned(3204, 12), 1598 => to_unsigned(857, 12), 1599 => to_unsigned(800, 12), 1600 => to_unsigned(1216, 12), 1601 => to_unsigned(2407, 12), 1602 => to_unsigned(1410, 12), 1603 => to_unsigned(2923, 12), 1604 => to_unsigned(1718, 12), 1605 => to_unsigned(3121, 12), 1606 => to_unsigned(2164, 12), 1607 => to_unsigned(3836, 12), 1608 => to_unsigned(4045, 12), 1609 => to_unsigned(2210, 12), 1610 => to_unsigned(2991, 12), 1611 => to_unsigned(1382, 12), 1612 => to_unsigned(4050, 12), 1613 => to_unsigned(932, 12), 1614 => to_unsigned(3472, 12), 1615 => to_unsigned(4024, 12), 1616 => to_unsigned(3637, 12), 1617 => to_unsigned(1955, 12), 1618 => to_unsigned(1149, 12), 1619 => to_unsigned(1072, 12), 1620 => to_unsigned(1128, 12), 1621 => to_unsigned(1961, 12), 1622 => to_unsigned(3223, 12), 1623 => to_unsigned(1505, 12), 1624 => to_unsigned(3646, 12), 1625 => to_unsigned(2754, 12), 1626 => to_unsigned(4054, 12), 1627 => to_unsigned(1886, 12), 1628 => to_unsigned(2909, 12), 1629 => to_unsigned(3848, 12), 1630 => to_unsigned(210, 12), 1631 => to_unsigned(1660, 12), 1632 => to_unsigned(3682, 12), 1633 => to_unsigned(2919, 12), 1634 => to_unsigned(3984, 12), 1635 => to_unsigned(1848, 12), 1636 => to_unsigned(225, 12), 1637 => to_unsigned(3094, 12), 1638 => to_unsigned(3615, 12), 1639 => to_unsigned(4019, 12), 1640 => to_unsigned(1883, 12), 1641 => to_unsigned(2298, 12), 1642 => to_unsigned(1540, 12), 1643 => to_unsigned(66, 12), 1644 => to_unsigned(1881, 12), 1645 => to_unsigned(794, 12), 1646 => to_unsigned(3955, 12), 1647 => to_unsigned(1535, 12), 1648 => to_unsigned(2645, 12), 1649 => to_unsigned(3811, 12), 1650 => to_unsigned(1517, 12), 1651 => to_unsigned(2921, 12), 1652 => to_unsigned(3224, 12), 1653 => to_unsigned(1605, 12), 1654 => to_unsigned(3840, 12), 1655 => to_unsigned(3898, 12), 1656 => to_unsigned(3939, 12), 1657 => to_unsigned(2365, 12), 1658 => to_unsigned(770, 12), 1659 => to_unsigned(2708, 12), 1660 => to_unsigned(2520, 12), 1661 => to_unsigned(781, 12), 1662 => to_unsigned(424, 12), 1663 => to_unsigned(3786, 12), 1664 => to_unsigned(3959, 12), 1665 => to_unsigned(1253, 12), 1666 => to_unsigned(2782, 12), 1667 => to_unsigned(2771, 12), 1668 => to_unsigned(3914, 12), 1669 => to_unsigned(2451, 12), 1670 => to_unsigned(1334, 12), 1671 => to_unsigned(3771, 12), 1672 => to_unsigned(2751, 12), 1673 => to_unsigned(2587, 12), 1674 => to_unsigned(1058, 12), 1675 => to_unsigned(2209, 12), 1676 => to_unsigned(2700, 12), 1677 => to_unsigned(218, 12), 1678 => to_unsigned(3875, 12), 1679 => to_unsigned(375, 12), 1680 => to_unsigned(247, 12), 1681 => to_unsigned(333, 12), 1682 => to_unsigned(290, 12), 1683 => to_unsigned(748, 12), 1684 => to_unsigned(122, 12), 1685 => to_unsigned(1328, 12), 1686 => to_unsigned(2657, 12), 1687 => to_unsigned(2504, 12), 1688 => to_unsigned(1208, 12), 1689 => to_unsigned(666, 12), 1690 => to_unsigned(796, 12), 1691 => to_unsigned(3484, 12), 1692 => to_unsigned(1971, 12), 1693 => to_unsigned(3792, 12), 1694 => to_unsigned(329, 12), 1695 => to_unsigned(3752, 12), 1696 => to_unsigned(3944, 12), 1697 => to_unsigned(324, 12), 1698 => to_unsigned(1285, 12), 1699 => to_unsigned(453, 12), 1700 => to_unsigned(787, 12), 1701 => to_unsigned(1380, 12), 1702 => to_unsigned(1218, 12), 1703 => to_unsigned(1250, 12), 1704 => to_unsigned(1267, 12), 1705 => to_unsigned(373, 12), 1706 => to_unsigned(160, 12), 1707 => to_unsigned(2515, 12), 1708 => to_unsigned(3254, 12), 1709 => to_unsigned(293, 12), 1710 => to_unsigned(1456, 12), 1711 => to_unsigned(1732, 12), 1712 => to_unsigned(3831, 12), 1713 => to_unsigned(3076, 12), 1714 => to_unsigned(2994, 12), 1715 => to_unsigned(1784, 12), 1716 => to_unsigned(4041, 12), 1717 => to_unsigned(754, 12), 1718 => to_unsigned(4085, 12), 1719 => to_unsigned(1095, 12), 1720 => to_unsigned(1152, 12), 1721 => to_unsigned(450, 12), 1722 => to_unsigned(3069, 12), 1723 => to_unsigned(1283, 12), 1724 => to_unsigned(3656, 12), 1725 => to_unsigned(2666, 12), 1726 => to_unsigned(3078, 12), 1727 => to_unsigned(1763, 12), 1728 => to_unsigned(2078, 12), 1729 => to_unsigned(3284, 12), 1730 => to_unsigned(1783, 12), 1731 => to_unsigned(3242, 12), 1732 => to_unsigned(2354, 12), 1733 => to_unsigned(3674, 12), 1734 => to_unsigned(170, 12), 1735 => to_unsigned(2026, 12), 1736 => to_unsigned(2085, 12), 1737 => to_unsigned(1318, 12), 1738 => to_unsigned(3044, 12), 1739 => to_unsigned(975, 12), 1740 => to_unsigned(242, 12), 1741 => to_unsigned(3330, 12), 1742 => to_unsigned(2105, 12), 1743 => to_unsigned(1685, 12), 1744 => to_unsigned(428, 12), 1745 => to_unsigned(176, 12), 1746 => to_unsigned(908, 12), 1747 => to_unsigned(143, 12), 1748 => to_unsigned(2187, 12), 1749 => to_unsigned(2453, 12), 1750 => to_unsigned(1409, 12), 1751 => to_unsigned(1101, 12), 1752 => to_unsigned(1553, 12), 1753 => to_unsigned(2169, 12), 1754 => to_unsigned(1189, 12), 1755 => to_unsigned(1957, 12), 1756 => to_unsigned(3801, 12), 1757 => to_unsigned(3956, 12), 1758 => to_unsigned(377, 12), 1759 => to_unsigned(4044, 12), 1760 => to_unsigned(909, 12), 1761 => to_unsigned(2999, 12), 1762 => to_unsigned(1761, 12), 1763 => to_unsigned(1923, 12), 1764 => to_unsigned(2352, 12), 1765 => to_unsigned(1200, 12), 1766 => to_unsigned(3876, 12), 1767 => to_unsigned(4095, 12), 1768 => to_unsigned(1445, 12), 1769 => to_unsigned(4071, 12), 1770 => to_unsigned(418, 12), 1771 => to_unsigned(3493, 12), 1772 => to_unsigned(2442, 12), 1773 => to_unsigned(3618, 12), 1774 => to_unsigned(861, 12), 1775 => to_unsigned(737, 12), 1776 => to_unsigned(3868, 12), 1777 => to_unsigned(3118, 12), 1778 => to_unsigned(2037, 12), 1779 => to_unsigned(1053, 12), 1780 => to_unsigned(2486, 12), 1781 => to_unsigned(2033, 12), 1782 => to_unsigned(734, 12), 1783 => to_unsigned(38, 12), 1784 => to_unsigned(2752, 12), 1785 => to_unsigned(2397, 12), 1786 => to_unsigned(3648, 12), 1787 => to_unsigned(1231, 12), 1788 => to_unsigned(1472, 12), 1789 => to_unsigned(486, 12), 1790 => to_unsigned(1423, 12), 1791 => to_unsigned(1030, 12), 1792 => to_unsigned(2566, 12), 1793 => to_unsigned(1672, 12), 1794 => to_unsigned(672, 12), 1795 => to_unsigned(3630, 12), 1796 => to_unsigned(2342, 12), 1797 => to_unsigned(366, 12), 1798 => to_unsigned(3307, 12), 1799 => to_unsigned(3234, 12), 1800 => to_unsigned(501, 12), 1801 => to_unsigned(896, 12), 1802 => to_unsigned(2736, 12), 1803 => to_unsigned(3939, 12), 1804 => to_unsigned(3988, 12), 1805 => to_unsigned(973, 12), 1806 => to_unsigned(435, 12), 1807 => to_unsigned(2231, 12), 1808 => to_unsigned(3799, 12), 1809 => to_unsigned(485, 12), 1810 => to_unsigned(12, 12), 1811 => to_unsigned(1562, 12), 1812 => to_unsigned(2718, 12), 1813 => to_unsigned(669, 12), 1814 => to_unsigned(633, 12), 1815 => to_unsigned(559, 12), 1816 => to_unsigned(1239, 12), 1817 => to_unsigned(3791, 12), 1818 => to_unsigned(2349, 12), 1819 => to_unsigned(2823, 12), 1820 => to_unsigned(757, 12), 1821 => to_unsigned(568, 12), 1822 => to_unsigned(916, 12), 1823 => to_unsigned(1259, 12), 1824 => to_unsigned(1272, 12), 1825 => to_unsigned(2819, 12), 1826 => to_unsigned(3551, 12), 1827 => to_unsigned(375, 12), 1828 => to_unsigned(314, 12), 1829 => to_unsigned(768, 12), 1830 => to_unsigned(2468, 12), 1831 => to_unsigned(3836, 12), 1832 => to_unsigned(2311, 12), 1833 => to_unsigned(1661, 12), 1834 => to_unsigned(2331, 12), 1835 => to_unsigned(1554, 12), 1836 => to_unsigned(3291, 12), 1837 => to_unsigned(942, 12), 1838 => to_unsigned(3874, 12), 1839 => to_unsigned(2386, 12), 1840 => to_unsigned(3311, 12), 1841 => to_unsigned(2418, 12), 1842 => to_unsigned(2560, 12), 1843 => to_unsigned(1629, 12), 1844 => to_unsigned(1017, 12), 1845 => to_unsigned(2422, 12), 1846 => to_unsigned(2525, 12), 1847 => to_unsigned(2039, 12), 1848 => to_unsigned(2844, 12), 1849 => to_unsigned(143, 12), 1850 => to_unsigned(2044, 12), 1851 => to_unsigned(4011, 12), 1852 => to_unsigned(1218, 12), 1853 => to_unsigned(2097, 12), 1854 => to_unsigned(3911, 12), 1855 => to_unsigned(774, 12), 1856 => to_unsigned(3268, 12), 1857 => to_unsigned(624, 12), 1858 => to_unsigned(2669, 12), 1859 => to_unsigned(2713, 12), 1860 => to_unsigned(2990, 12), 1861 => to_unsigned(1488, 12), 1862 => to_unsigned(3836, 12), 1863 => to_unsigned(75, 12), 1864 => to_unsigned(489, 12), 1865 => to_unsigned(836, 12), 1866 => to_unsigned(2334, 12), 1867 => to_unsigned(3834, 12), 1868 => to_unsigned(1432, 12), 1869 => to_unsigned(372, 12), 1870 => to_unsigned(774, 12), 1871 => to_unsigned(1206, 12), 1872 => to_unsigned(311, 12), 1873 => to_unsigned(1650, 12), 1874 => to_unsigned(480, 12), 1875 => to_unsigned(4055, 12), 1876 => to_unsigned(3155, 12), 1877 => to_unsigned(1381, 12), 1878 => to_unsigned(2214, 12), 1879 => to_unsigned(2598, 12), 1880 => to_unsigned(3898, 12), 1881 => to_unsigned(2884, 12), 1882 => to_unsigned(204, 12), 1883 => to_unsigned(3537, 12), 1884 => to_unsigned(702, 12), 1885 => to_unsigned(1672, 12), 1886 => to_unsigned(1569, 12), 1887 => to_unsigned(1225, 12), 1888 => to_unsigned(3623, 12), 1889 => to_unsigned(1060, 12), 1890 => to_unsigned(2002, 12), 1891 => to_unsigned(2560, 12), 1892 => to_unsigned(1656, 12), 1893 => to_unsigned(528, 12), 1894 => to_unsigned(619, 12), 1895 => to_unsigned(1351, 12), 1896 => to_unsigned(3890, 12), 1897 => to_unsigned(2487, 12), 1898 => to_unsigned(2353, 12), 1899 => to_unsigned(1458, 12), 1900 => to_unsigned(1767, 12), 1901 => to_unsigned(210, 12), 1902 => to_unsigned(3460, 12), 1903 => to_unsigned(153, 12), 1904 => to_unsigned(1802, 12), 1905 => to_unsigned(1120, 12), 1906 => to_unsigned(3117, 12), 1907 => to_unsigned(341, 12), 1908 => to_unsigned(3426, 12), 1909 => to_unsigned(3508, 12), 1910 => to_unsigned(3342, 12), 1911 => to_unsigned(1310, 12), 1912 => to_unsigned(74, 12), 1913 => to_unsigned(327, 12), 1914 => to_unsigned(3152, 12), 1915 => to_unsigned(4076, 12), 1916 => to_unsigned(27, 12), 1917 => to_unsigned(1900, 12), 1918 => to_unsigned(1076, 12), 1919 => to_unsigned(416, 12), 1920 => to_unsigned(3495, 12), 1921 => to_unsigned(631, 12), 1922 => to_unsigned(3512, 12), 1923 => to_unsigned(2045, 12), 1924 => to_unsigned(3607, 12), 1925 => to_unsigned(242, 12), 1926 => to_unsigned(829, 12), 1927 => to_unsigned(2886, 12), 1928 => to_unsigned(1164, 12), 1929 => to_unsigned(627, 12), 1930 => to_unsigned(3460, 12), 1931 => to_unsigned(1938, 12), 1932 => to_unsigned(590, 12), 1933 => to_unsigned(2836, 12), 1934 => to_unsigned(3941, 12), 1935 => to_unsigned(1208, 12), 1936 => to_unsigned(1827, 12), 1937 => to_unsigned(1350, 12), 1938 => to_unsigned(1260, 12), 1939 => to_unsigned(29, 12), 1940 => to_unsigned(3195, 12), 1941 => to_unsigned(3210, 12), 1942 => to_unsigned(3290, 12), 1943 => to_unsigned(386, 12), 1944 => to_unsigned(2518, 12), 1945 => to_unsigned(613, 12), 1946 => to_unsigned(2449, 12), 1947 => to_unsigned(2094, 12), 1948 => to_unsigned(2785, 12), 1949 => to_unsigned(2332, 12), 1950 => to_unsigned(1202, 12), 1951 => to_unsigned(3010, 12), 1952 => to_unsigned(41, 12), 1953 => to_unsigned(3528, 12), 1954 => to_unsigned(1426, 12), 1955 => to_unsigned(2444, 12), 1956 => to_unsigned(3281, 12), 1957 => to_unsigned(1517, 12), 1958 => to_unsigned(1717, 12), 1959 => to_unsigned(284, 12), 1960 => to_unsigned(360, 12), 1961 => to_unsigned(249, 12), 1962 => to_unsigned(274, 12), 1963 => to_unsigned(591, 12), 1964 => to_unsigned(3900, 12), 1965 => to_unsigned(3456, 12), 1966 => to_unsigned(2678, 12), 1967 => to_unsigned(2988, 12), 1968 => to_unsigned(1668, 12), 1969 => to_unsigned(3533, 12), 1970 => to_unsigned(1454, 12), 1971 => to_unsigned(2797, 12), 1972 => to_unsigned(1227, 12), 1973 => to_unsigned(2715, 12), 1974 => to_unsigned(2795, 12), 1975 => to_unsigned(4027, 12), 1976 => to_unsigned(903, 12), 1977 => to_unsigned(693, 12), 1978 => to_unsigned(664, 12), 1979 => to_unsigned(11, 12), 1980 => to_unsigned(2842, 12), 1981 => to_unsigned(1123, 12), 1982 => to_unsigned(959, 12), 1983 => to_unsigned(2703, 12), 1984 => to_unsigned(2252, 12), 1985 => to_unsigned(718, 12), 1986 => to_unsigned(2758, 12), 1987 => to_unsigned(1298, 12), 1988 => to_unsigned(1395, 12), 1989 => to_unsigned(508, 12), 1990 => to_unsigned(1640, 12), 1991 => to_unsigned(2063, 12), 1992 => to_unsigned(2990, 12), 1993 => to_unsigned(3028, 12), 1994 => to_unsigned(3921, 12), 1995 => to_unsigned(3016, 12), 1996 => to_unsigned(1884, 12), 1997 => to_unsigned(1934, 12), 1998 => to_unsigned(2209, 12), 1999 => to_unsigned(2357, 12), 2000 => to_unsigned(95, 12), 2001 => to_unsigned(1675, 12), 2002 => to_unsigned(309, 12), 2003 => to_unsigned(1033, 12), 2004 => to_unsigned(108, 12), 2005 => to_unsigned(1312, 12), 2006 => to_unsigned(751, 12), 2007 => to_unsigned(1128, 12), 2008 => to_unsigned(341, 12), 2009 => to_unsigned(1639, 12), 2010 => to_unsigned(2698, 12), 2011 => to_unsigned(1249, 12), 2012 => to_unsigned(2441, 12), 2013 => to_unsigned(540, 12), 2014 => to_unsigned(1154, 12), 2015 => to_unsigned(3962, 12), 2016 => to_unsigned(3725, 12), 2017 => to_unsigned(1274, 12), 2018 => to_unsigned(234, 12), 2019 => to_unsigned(1803, 12), 2020 => to_unsigned(3918, 12), 2021 => to_unsigned(109, 12), 2022 => to_unsigned(985, 12), 2023 => to_unsigned(1024, 12), 2024 => to_unsigned(2008, 12), 2025 => to_unsigned(747, 12), 2026 => to_unsigned(2503, 12), 2027 => to_unsigned(2066, 12), 2028 => to_unsigned(2739, 12), 2029 => to_unsigned(897, 12), 2030 => to_unsigned(1727, 12), 2031 => to_unsigned(2052, 12), 2032 => to_unsigned(2854, 12), 2033 => to_unsigned(2725, 12), 2034 => to_unsigned(1657, 12), 2035 => to_unsigned(3452, 12), 2036 => to_unsigned(1362, 12), 2037 => to_unsigned(3301, 12), 2038 => to_unsigned(1208, 12), 2039 => to_unsigned(1289, 12), 2040 => to_unsigned(721, 12), 2041 => to_unsigned(104, 12), 2042 => to_unsigned(3174, 12), 2043 => to_unsigned(852, 12), 2044 => to_unsigned(2829, 12), 2045 => to_unsigned(559, 12), 2046 => to_unsigned(282, 12), 2047 => to_unsigned(825, 12)),
            5 => (0 => to_unsigned(1731, 12), 1 => to_unsigned(2321, 12), 2 => to_unsigned(3872, 12), 3 => to_unsigned(3854, 12), 4 => to_unsigned(971, 12), 5 => to_unsigned(359, 12), 6 => to_unsigned(1193, 12), 7 => to_unsigned(1434, 12), 8 => to_unsigned(568, 12), 9 => to_unsigned(851, 12), 10 => to_unsigned(2051, 12), 11 => to_unsigned(2706, 12), 12 => to_unsigned(46, 12), 13 => to_unsigned(32, 12), 14 => to_unsigned(2417, 12), 15 => to_unsigned(2488, 12), 16 => to_unsigned(1810, 12), 17 => to_unsigned(4084, 12), 18 => to_unsigned(3522, 12), 19 => to_unsigned(2360, 12), 20 => to_unsigned(3039, 12), 21 => to_unsigned(1020, 12), 22 => to_unsigned(3140, 12), 23 => to_unsigned(3396, 12), 24 => to_unsigned(3846, 12), 25 => to_unsigned(1523, 12), 26 => to_unsigned(2502, 12), 27 => to_unsigned(1153, 12), 28 => to_unsigned(3661, 12), 29 => to_unsigned(514, 12), 30 => to_unsigned(1461, 12), 31 => to_unsigned(848, 12), 32 => to_unsigned(2639, 12), 33 => to_unsigned(1038, 12), 34 => to_unsigned(114, 12), 35 => to_unsigned(3335, 12), 36 => to_unsigned(3531, 12), 37 => to_unsigned(594, 12), 38 => to_unsigned(2467, 12), 39 => to_unsigned(2679, 12), 40 => to_unsigned(131, 12), 41 => to_unsigned(3968, 12), 42 => to_unsigned(3245, 12), 43 => to_unsigned(1716, 12), 44 => to_unsigned(3219, 12), 45 => to_unsigned(2791, 12), 46 => to_unsigned(2805, 12), 47 => to_unsigned(1746, 12), 48 => to_unsigned(368, 12), 49 => to_unsigned(266, 12), 50 => to_unsigned(2285, 12), 51 => to_unsigned(3117, 12), 52 => to_unsigned(1249, 12), 53 => to_unsigned(1623, 12), 54 => to_unsigned(1048, 12), 55 => to_unsigned(2006, 12), 56 => to_unsigned(2637, 12), 57 => to_unsigned(1503, 12), 58 => to_unsigned(3583, 12), 59 => to_unsigned(2571, 12), 60 => to_unsigned(3205, 12), 61 => to_unsigned(309, 12), 62 => to_unsigned(1906, 12), 63 => to_unsigned(546, 12), 64 => to_unsigned(2168, 12), 65 => to_unsigned(843, 12), 66 => to_unsigned(929, 12), 67 => to_unsigned(2438, 12), 68 => to_unsigned(408, 12), 69 => to_unsigned(3136, 12), 70 => to_unsigned(1541, 12), 71 => to_unsigned(3503, 12), 72 => to_unsigned(866, 12), 73 => to_unsigned(1055, 12), 74 => to_unsigned(3419, 12), 75 => to_unsigned(3854, 12), 76 => to_unsigned(3720, 12), 77 => to_unsigned(254, 12), 78 => to_unsigned(3731, 12), 79 => to_unsigned(1780, 12), 80 => to_unsigned(2391, 12), 81 => to_unsigned(2023, 12), 82 => to_unsigned(2934, 12), 83 => to_unsigned(1796, 12), 84 => to_unsigned(3736, 12), 85 => to_unsigned(396, 12), 86 => to_unsigned(841, 12), 87 => to_unsigned(77, 12), 88 => to_unsigned(3219, 12), 89 => to_unsigned(2047, 12), 90 => to_unsigned(3819, 12), 91 => to_unsigned(2085, 12), 92 => to_unsigned(343, 12), 93 => to_unsigned(3213, 12), 94 => to_unsigned(2194, 12), 95 => to_unsigned(3647, 12), 96 => to_unsigned(1516, 12), 97 => to_unsigned(1229, 12), 98 => to_unsigned(369, 12), 99 => to_unsigned(314, 12), 100 => to_unsigned(2958, 12), 101 => to_unsigned(4010, 12), 102 => to_unsigned(3087, 12), 103 => to_unsigned(1409, 12), 104 => to_unsigned(3510, 12), 105 => to_unsigned(3277, 12), 106 => to_unsigned(2095, 12), 107 => to_unsigned(435, 12), 108 => to_unsigned(2595, 12), 109 => to_unsigned(1720, 12), 110 => to_unsigned(193, 12), 111 => to_unsigned(3982, 12), 112 => to_unsigned(2183, 12), 113 => to_unsigned(2572, 12), 114 => to_unsigned(286, 12), 115 => to_unsigned(3572, 12), 116 => to_unsigned(3359, 12), 117 => to_unsigned(3581, 12), 118 => to_unsigned(1040, 12), 119 => to_unsigned(1221, 12), 120 => to_unsigned(491, 12), 121 => to_unsigned(425, 12), 122 => to_unsigned(2437, 12), 123 => to_unsigned(1816, 12), 124 => to_unsigned(800, 12), 125 => to_unsigned(651, 12), 126 => to_unsigned(52, 12), 127 => to_unsigned(892, 12), 128 => to_unsigned(3237, 12), 129 => to_unsigned(3431, 12), 130 => to_unsigned(1521, 12), 131 => to_unsigned(1884, 12), 132 => to_unsigned(4002, 12), 133 => to_unsigned(2205, 12), 134 => to_unsigned(3957, 12), 135 => to_unsigned(1223, 12), 136 => to_unsigned(3132, 12), 137 => to_unsigned(3551, 12), 138 => to_unsigned(2467, 12), 139 => to_unsigned(2476, 12), 140 => to_unsigned(70, 12), 141 => to_unsigned(3714, 12), 142 => to_unsigned(524, 12), 143 => to_unsigned(2812, 12), 144 => to_unsigned(3987, 12), 145 => to_unsigned(3956, 12), 146 => to_unsigned(3040, 12), 147 => to_unsigned(3941, 12), 148 => to_unsigned(3176, 12), 149 => to_unsigned(1363, 12), 150 => to_unsigned(1864, 12), 151 => to_unsigned(951, 12), 152 => to_unsigned(2064, 12), 153 => to_unsigned(613, 12), 154 => to_unsigned(98, 12), 155 => to_unsigned(2641, 12), 156 => to_unsigned(2105, 12), 157 => to_unsigned(125, 12), 158 => to_unsigned(1645, 12), 159 => to_unsigned(1890, 12), 160 => to_unsigned(1257, 12), 161 => to_unsigned(1608, 12), 162 => to_unsigned(2213, 12), 163 => to_unsigned(2783, 12), 164 => to_unsigned(307, 12), 165 => to_unsigned(323, 12), 166 => to_unsigned(817, 12), 167 => to_unsigned(1432, 12), 168 => to_unsigned(457, 12), 169 => to_unsigned(1757, 12), 170 => to_unsigned(262, 12), 171 => to_unsigned(59, 12), 172 => to_unsigned(1005, 12), 173 => to_unsigned(2467, 12), 174 => to_unsigned(2829, 12), 175 => to_unsigned(2321, 12), 176 => to_unsigned(2974, 12), 177 => to_unsigned(1234, 12), 178 => to_unsigned(1617, 12), 179 => to_unsigned(3992, 12), 180 => to_unsigned(1707, 12), 181 => to_unsigned(2836, 12), 182 => to_unsigned(2639, 12), 183 => to_unsigned(3684, 12), 184 => to_unsigned(978, 12), 185 => to_unsigned(261, 12), 186 => to_unsigned(2133, 12), 187 => to_unsigned(3839, 12), 188 => to_unsigned(2545, 12), 189 => to_unsigned(437, 12), 190 => to_unsigned(479, 12), 191 => to_unsigned(721, 12), 192 => to_unsigned(2690, 12), 193 => to_unsigned(1404, 12), 194 => to_unsigned(1193, 12), 195 => to_unsigned(2998, 12), 196 => to_unsigned(281, 12), 197 => to_unsigned(2323, 12), 198 => to_unsigned(2253, 12), 199 => to_unsigned(3292, 12), 200 => to_unsigned(3793, 12), 201 => to_unsigned(1009, 12), 202 => to_unsigned(3797, 12), 203 => to_unsigned(837, 12), 204 => to_unsigned(1424, 12), 205 => to_unsigned(2745, 12), 206 => to_unsigned(1991, 12), 207 => to_unsigned(2129, 12), 208 => to_unsigned(3299, 12), 209 => to_unsigned(3375, 12), 210 => to_unsigned(730, 12), 211 => to_unsigned(1613, 12), 212 => to_unsigned(3477, 12), 213 => to_unsigned(1414, 12), 214 => to_unsigned(1030, 12), 215 => to_unsigned(3386, 12), 216 => to_unsigned(2452, 12), 217 => to_unsigned(3010, 12), 218 => to_unsigned(195, 12), 219 => to_unsigned(1905, 12), 220 => to_unsigned(832, 12), 221 => to_unsigned(1021, 12), 222 => to_unsigned(930, 12), 223 => to_unsigned(2916, 12), 224 => to_unsigned(3493, 12), 225 => to_unsigned(1967, 12), 226 => to_unsigned(2441, 12), 227 => to_unsigned(2236, 12), 228 => to_unsigned(654, 12), 229 => to_unsigned(3005, 12), 230 => to_unsigned(60, 12), 231 => to_unsigned(782, 12), 232 => to_unsigned(1144, 12), 233 => to_unsigned(620, 12), 234 => to_unsigned(3897, 12), 235 => to_unsigned(2784, 12), 236 => to_unsigned(3100, 12), 237 => to_unsigned(2719, 12), 238 => to_unsigned(3677, 12), 239 => to_unsigned(2366, 12), 240 => to_unsigned(3311, 12), 241 => to_unsigned(480, 12), 242 => to_unsigned(2674, 12), 243 => to_unsigned(3042, 12), 244 => to_unsigned(849, 12), 245 => to_unsigned(272, 12), 246 => to_unsigned(1437, 12), 247 => to_unsigned(95, 12), 248 => to_unsigned(2904, 12), 249 => to_unsigned(1099, 12), 250 => to_unsigned(3956, 12), 251 => to_unsigned(3244, 12), 252 => to_unsigned(1333, 12), 253 => to_unsigned(2838, 12), 254 => to_unsigned(645, 12), 255 => to_unsigned(1461, 12), 256 => to_unsigned(1033, 12), 257 => to_unsigned(616, 12), 258 => to_unsigned(3284, 12), 259 => to_unsigned(1913, 12), 260 => to_unsigned(1239, 12), 261 => to_unsigned(1983, 12), 262 => to_unsigned(2101, 12), 263 => to_unsigned(1144, 12), 264 => to_unsigned(2883, 12), 265 => to_unsigned(3495, 12), 266 => to_unsigned(1470, 12), 267 => to_unsigned(405, 12), 268 => to_unsigned(2803, 12), 269 => to_unsigned(3130, 12), 270 => to_unsigned(504, 12), 271 => to_unsigned(1291, 12), 272 => to_unsigned(804, 12), 273 => to_unsigned(2186, 12), 274 => to_unsigned(440, 12), 275 => to_unsigned(710, 12), 276 => to_unsigned(635, 12), 277 => to_unsigned(1524, 12), 278 => to_unsigned(3818, 12), 279 => to_unsigned(2870, 12), 280 => to_unsigned(3769, 12), 281 => to_unsigned(2469, 12), 282 => to_unsigned(967, 12), 283 => to_unsigned(2696, 12), 284 => to_unsigned(1632, 12), 285 => to_unsigned(3985, 12), 286 => to_unsigned(2092, 12), 287 => to_unsigned(4008, 12), 288 => to_unsigned(121, 12), 289 => to_unsigned(2108, 12), 290 => to_unsigned(346, 12), 291 => to_unsigned(2016, 12), 292 => to_unsigned(1332, 12), 293 => to_unsigned(1158, 12), 294 => to_unsigned(3477, 12), 295 => to_unsigned(889, 12), 296 => to_unsigned(3568, 12), 297 => to_unsigned(1737, 12), 298 => to_unsigned(99, 12), 299 => to_unsigned(1162, 12), 300 => to_unsigned(743, 12), 301 => to_unsigned(1959, 12), 302 => to_unsigned(2537, 12), 303 => to_unsigned(2611, 12), 304 => to_unsigned(1202, 12), 305 => to_unsigned(2526, 12), 306 => to_unsigned(3670, 12), 307 => to_unsigned(2260, 12), 308 => to_unsigned(1933, 12), 309 => to_unsigned(1672, 12), 310 => to_unsigned(1450, 12), 311 => to_unsigned(3020, 12), 312 => to_unsigned(1242, 12), 313 => to_unsigned(3097, 12), 314 => to_unsigned(857, 12), 315 => to_unsigned(756, 12), 316 => to_unsigned(3126, 12), 317 => to_unsigned(1496, 12), 318 => to_unsigned(51, 12), 319 => to_unsigned(2266, 12), 320 => to_unsigned(3981, 12), 321 => to_unsigned(1319, 12), 322 => to_unsigned(1394, 12), 323 => to_unsigned(1594, 12), 324 => to_unsigned(975, 12), 325 => to_unsigned(3873, 12), 326 => to_unsigned(3845, 12), 327 => to_unsigned(3954, 12), 328 => to_unsigned(2969, 12), 329 => to_unsigned(3878, 12), 330 => to_unsigned(3062, 12), 331 => to_unsigned(729, 12), 332 => to_unsigned(2743, 12), 333 => to_unsigned(3393, 12), 334 => to_unsigned(337, 12), 335 => to_unsigned(1932, 12), 336 => to_unsigned(3627, 12), 337 => to_unsigned(733, 12), 338 => to_unsigned(3360, 12), 339 => to_unsigned(851, 12), 340 => to_unsigned(2453, 12), 341 => to_unsigned(268, 12), 342 => to_unsigned(749, 12), 343 => to_unsigned(3392, 12), 344 => to_unsigned(401, 12), 345 => to_unsigned(517, 12), 346 => to_unsigned(3721, 12), 347 => to_unsigned(1150, 12), 348 => to_unsigned(2148, 12), 349 => to_unsigned(394, 12), 350 => to_unsigned(3650, 12), 351 => to_unsigned(1096, 12), 352 => to_unsigned(1119, 12), 353 => to_unsigned(2071, 12), 354 => to_unsigned(3266, 12), 355 => to_unsigned(253, 12), 356 => to_unsigned(2690, 12), 357 => to_unsigned(2538, 12), 358 => to_unsigned(2265, 12), 359 => to_unsigned(3885, 12), 360 => to_unsigned(2461, 12), 361 => to_unsigned(935, 12), 362 => to_unsigned(2621, 12), 363 => to_unsigned(318, 12), 364 => to_unsigned(1104, 12), 365 => to_unsigned(852, 12), 366 => to_unsigned(3223, 12), 367 => to_unsigned(2537, 12), 368 => to_unsigned(293, 12), 369 => to_unsigned(4065, 12), 370 => to_unsigned(3044, 12), 371 => to_unsigned(477, 12), 372 => to_unsigned(82, 12), 373 => to_unsigned(1243, 12), 374 => to_unsigned(3680, 12), 375 => to_unsigned(3443, 12), 376 => to_unsigned(3154, 12), 377 => to_unsigned(3728, 12), 378 => to_unsigned(0, 12), 379 => to_unsigned(907, 12), 380 => to_unsigned(2335, 12), 381 => to_unsigned(192, 12), 382 => to_unsigned(2730, 12), 383 => to_unsigned(1287, 12), 384 => to_unsigned(468, 12), 385 => to_unsigned(2290, 12), 386 => to_unsigned(514, 12), 387 => to_unsigned(1661, 12), 388 => to_unsigned(1261, 12), 389 => to_unsigned(2099, 12), 390 => to_unsigned(695, 12), 391 => to_unsigned(3226, 12), 392 => to_unsigned(3879, 12), 393 => to_unsigned(1262, 12), 394 => to_unsigned(360, 12), 395 => to_unsigned(2046, 12), 396 => to_unsigned(925, 12), 397 => to_unsigned(3538, 12), 398 => to_unsigned(2217, 12), 399 => to_unsigned(2585, 12), 400 => to_unsigned(2988, 12), 401 => to_unsigned(770, 12), 402 => to_unsigned(334, 12), 403 => to_unsigned(2474, 12), 404 => to_unsigned(1922, 12), 405 => to_unsigned(1122, 12), 406 => to_unsigned(915, 12), 407 => to_unsigned(502, 12), 408 => to_unsigned(811, 12), 409 => to_unsigned(2825, 12), 410 => to_unsigned(844, 12), 411 => to_unsigned(2154, 12), 412 => to_unsigned(1153, 12), 413 => to_unsigned(2458, 12), 414 => to_unsigned(2240, 12), 415 => to_unsigned(153, 12), 416 => to_unsigned(3453, 12), 417 => to_unsigned(2756, 12), 418 => to_unsigned(3921, 12), 419 => to_unsigned(40, 12), 420 => to_unsigned(3590, 12), 421 => to_unsigned(3335, 12), 422 => to_unsigned(3513, 12), 423 => to_unsigned(3628, 12), 424 => to_unsigned(3505, 12), 425 => to_unsigned(1610, 12), 426 => to_unsigned(2699, 12), 427 => to_unsigned(743, 12), 428 => to_unsigned(337, 12), 429 => to_unsigned(1943, 12), 430 => to_unsigned(3102, 12), 431 => to_unsigned(1065, 12), 432 => to_unsigned(3901, 12), 433 => to_unsigned(3208, 12), 434 => to_unsigned(2386, 12), 435 => to_unsigned(1241, 12), 436 => to_unsigned(925, 12), 437 => to_unsigned(121, 12), 438 => to_unsigned(3873, 12), 439 => to_unsigned(3267, 12), 440 => to_unsigned(3864, 12), 441 => to_unsigned(1664, 12), 442 => to_unsigned(4013, 12), 443 => to_unsigned(3401, 12), 444 => to_unsigned(2760, 12), 445 => to_unsigned(29, 12), 446 => to_unsigned(1294, 12), 447 => to_unsigned(2595, 12), 448 => to_unsigned(598, 12), 449 => to_unsigned(3202, 12), 450 => to_unsigned(3347, 12), 451 => to_unsigned(1563, 12), 452 => to_unsigned(2714, 12), 453 => to_unsigned(1429, 12), 454 => to_unsigned(3519, 12), 455 => to_unsigned(3378, 12), 456 => to_unsigned(8, 12), 457 => to_unsigned(1214, 12), 458 => to_unsigned(3421, 12), 459 => to_unsigned(2791, 12), 460 => to_unsigned(1873, 12), 461 => to_unsigned(3146, 12), 462 => to_unsigned(3624, 12), 463 => to_unsigned(2957, 12), 464 => to_unsigned(3217, 12), 465 => to_unsigned(2681, 12), 466 => to_unsigned(3151, 12), 467 => to_unsigned(2615, 12), 468 => to_unsigned(1236, 12), 469 => to_unsigned(2274, 12), 470 => to_unsigned(2780, 12), 471 => to_unsigned(419, 12), 472 => to_unsigned(3338, 12), 473 => to_unsigned(2942, 12), 474 => to_unsigned(199, 12), 475 => to_unsigned(3119, 12), 476 => to_unsigned(589, 12), 477 => to_unsigned(3705, 12), 478 => to_unsigned(3640, 12), 479 => to_unsigned(3189, 12), 480 => to_unsigned(3842, 12), 481 => to_unsigned(3271, 12), 482 => to_unsigned(2809, 12), 483 => to_unsigned(983, 12), 484 => to_unsigned(1719, 12), 485 => to_unsigned(665, 12), 486 => to_unsigned(1309, 12), 487 => to_unsigned(3294, 12), 488 => to_unsigned(607, 12), 489 => to_unsigned(2267, 12), 490 => to_unsigned(3297, 12), 491 => to_unsigned(3477, 12), 492 => to_unsigned(321, 12), 493 => to_unsigned(257, 12), 494 => to_unsigned(3449, 12), 495 => to_unsigned(3211, 12), 496 => to_unsigned(2543, 12), 497 => to_unsigned(2635, 12), 498 => to_unsigned(874, 12), 499 => to_unsigned(1176, 12), 500 => to_unsigned(1345, 12), 501 => to_unsigned(3309, 12), 502 => to_unsigned(1981, 12), 503 => to_unsigned(1168, 12), 504 => to_unsigned(3854, 12), 505 => to_unsigned(2501, 12), 506 => to_unsigned(2003, 12), 507 => to_unsigned(2573, 12), 508 => to_unsigned(785, 12), 509 => to_unsigned(3493, 12), 510 => to_unsigned(1643, 12), 511 => to_unsigned(2843, 12), 512 => to_unsigned(3885, 12), 513 => to_unsigned(3145, 12), 514 => to_unsigned(305, 12), 515 => to_unsigned(165, 12), 516 => to_unsigned(1085, 12), 517 => to_unsigned(3856, 12), 518 => to_unsigned(3505, 12), 519 => to_unsigned(458, 12), 520 => to_unsigned(1945, 12), 521 => to_unsigned(1660, 12), 522 => to_unsigned(664, 12), 523 => to_unsigned(1125, 12), 524 => to_unsigned(3461, 12), 525 => to_unsigned(2106, 12), 526 => to_unsigned(2176, 12), 527 => to_unsigned(2890, 12), 528 => to_unsigned(3501, 12), 529 => to_unsigned(1575, 12), 530 => to_unsigned(2994, 12), 531 => to_unsigned(1932, 12), 532 => to_unsigned(1494, 12), 533 => to_unsigned(1302, 12), 534 => to_unsigned(313, 12), 535 => to_unsigned(1472, 12), 536 => to_unsigned(3554, 12), 537 => to_unsigned(1669, 12), 538 => to_unsigned(897, 12), 539 => to_unsigned(3011, 12), 540 => to_unsigned(2382, 12), 541 => to_unsigned(2430, 12), 542 => to_unsigned(1880, 12), 543 => to_unsigned(2354, 12), 544 => to_unsigned(301, 12), 545 => to_unsigned(3939, 12), 546 => to_unsigned(3786, 12), 547 => to_unsigned(3932, 12), 548 => to_unsigned(3668, 12), 549 => to_unsigned(2671, 12), 550 => to_unsigned(829, 12), 551 => to_unsigned(947, 12), 552 => to_unsigned(3344, 12), 553 => to_unsigned(3610, 12), 554 => to_unsigned(2309, 12), 555 => to_unsigned(1437, 12), 556 => to_unsigned(596, 12), 557 => to_unsigned(4007, 12), 558 => to_unsigned(2678, 12), 559 => to_unsigned(1915, 12), 560 => to_unsigned(231, 12), 561 => to_unsigned(1360, 12), 562 => to_unsigned(2484, 12), 563 => to_unsigned(20, 12), 564 => to_unsigned(3385, 12), 565 => to_unsigned(1275, 12), 566 => to_unsigned(3018, 12), 567 => to_unsigned(3255, 12), 568 => to_unsigned(276, 12), 569 => to_unsigned(459, 12), 570 => to_unsigned(1164, 12), 571 => to_unsigned(1649, 12), 572 => to_unsigned(725, 12), 573 => to_unsigned(145, 12), 574 => to_unsigned(61, 12), 575 => to_unsigned(833, 12), 576 => to_unsigned(1103, 12), 577 => to_unsigned(2000, 12), 578 => to_unsigned(2021, 12), 579 => to_unsigned(1436, 12), 580 => to_unsigned(2672, 12), 581 => to_unsigned(3682, 12), 582 => to_unsigned(3163, 12), 583 => to_unsigned(682, 12), 584 => to_unsigned(216, 12), 585 => to_unsigned(2927, 12), 586 => to_unsigned(723, 12), 587 => to_unsigned(2766, 12), 588 => to_unsigned(2679, 12), 589 => to_unsigned(2628, 12), 590 => to_unsigned(1265, 12), 591 => to_unsigned(2998, 12), 592 => to_unsigned(1326, 12), 593 => to_unsigned(451, 12), 594 => to_unsigned(2902, 12), 595 => to_unsigned(3408, 12), 596 => to_unsigned(1102, 12), 597 => to_unsigned(3441, 12), 598 => to_unsigned(2627, 12), 599 => to_unsigned(2735, 12), 600 => to_unsigned(3409, 12), 601 => to_unsigned(1750, 12), 602 => to_unsigned(1829, 12), 603 => to_unsigned(3662, 12), 604 => to_unsigned(3241, 12), 605 => to_unsigned(3159, 12), 606 => to_unsigned(632, 12), 607 => to_unsigned(624, 12), 608 => to_unsigned(2401, 12), 609 => to_unsigned(499, 12), 610 => to_unsigned(1668, 12), 611 => to_unsigned(1795, 12), 612 => to_unsigned(1962, 12), 613 => to_unsigned(3490, 12), 614 => to_unsigned(2424, 12), 615 => to_unsigned(3428, 12), 616 => to_unsigned(2908, 12), 617 => to_unsigned(1719, 12), 618 => to_unsigned(1420, 12), 619 => to_unsigned(487, 12), 620 => to_unsigned(3276, 12), 621 => to_unsigned(3526, 12), 622 => to_unsigned(221, 12), 623 => to_unsigned(456, 12), 624 => to_unsigned(3097, 12), 625 => to_unsigned(2585, 12), 626 => to_unsigned(1302, 12), 627 => to_unsigned(5, 12), 628 => to_unsigned(371, 12), 629 => to_unsigned(819, 12), 630 => to_unsigned(3208, 12), 631 => to_unsigned(1405, 12), 632 => to_unsigned(1750, 12), 633 => to_unsigned(2876, 12), 634 => to_unsigned(1396, 12), 635 => to_unsigned(3722, 12), 636 => to_unsigned(23, 12), 637 => to_unsigned(1621, 12), 638 => to_unsigned(507, 12), 639 => to_unsigned(2359, 12), 640 => to_unsigned(881, 12), 641 => to_unsigned(1451, 12), 642 => to_unsigned(2326, 12), 643 => to_unsigned(812, 12), 644 => to_unsigned(492, 12), 645 => to_unsigned(264, 12), 646 => to_unsigned(81, 12), 647 => to_unsigned(367, 12), 648 => to_unsigned(2971, 12), 649 => to_unsigned(2899, 12), 650 => to_unsigned(2649, 12), 651 => to_unsigned(2225, 12), 652 => to_unsigned(2025, 12), 653 => to_unsigned(1646, 12), 654 => to_unsigned(3454, 12), 655 => to_unsigned(443, 12), 656 => to_unsigned(2644, 12), 657 => to_unsigned(779, 12), 658 => to_unsigned(3424, 12), 659 => to_unsigned(2561, 12), 660 => to_unsigned(3534, 12), 661 => to_unsigned(641, 12), 662 => to_unsigned(101, 12), 663 => to_unsigned(3173, 12), 664 => to_unsigned(2665, 12), 665 => to_unsigned(2227, 12), 666 => to_unsigned(1402, 12), 667 => to_unsigned(1577, 12), 668 => to_unsigned(2672, 12), 669 => to_unsigned(3634, 12), 670 => to_unsigned(3993, 12), 671 => to_unsigned(1898, 12), 672 => to_unsigned(125, 12), 673 => to_unsigned(3680, 12), 674 => to_unsigned(2683, 12), 675 => to_unsigned(1238, 12), 676 => to_unsigned(2935, 12), 677 => to_unsigned(80, 12), 678 => to_unsigned(403, 12), 679 => to_unsigned(3393, 12), 680 => to_unsigned(1548, 12), 681 => to_unsigned(1283, 12), 682 => to_unsigned(1205, 12), 683 => to_unsigned(3866, 12), 684 => to_unsigned(3568, 12), 685 => to_unsigned(2698, 12), 686 => to_unsigned(3248, 12), 687 => to_unsigned(2277, 12), 688 => to_unsigned(2227, 12), 689 => to_unsigned(2761, 12), 690 => to_unsigned(4046, 12), 691 => to_unsigned(3830, 12), 692 => to_unsigned(2528, 12), 693 => to_unsigned(1279, 12), 694 => to_unsigned(2768, 12), 695 => to_unsigned(2288, 12), 696 => to_unsigned(1543, 12), 697 => to_unsigned(3756, 12), 698 => to_unsigned(3505, 12), 699 => to_unsigned(2218, 12), 700 => to_unsigned(3227, 12), 701 => to_unsigned(3233, 12), 702 => to_unsigned(349, 12), 703 => to_unsigned(2963, 12), 704 => to_unsigned(1568, 12), 705 => to_unsigned(1037, 12), 706 => to_unsigned(3102, 12), 707 => to_unsigned(712, 12), 708 => to_unsigned(2362, 12), 709 => to_unsigned(2567, 12), 710 => to_unsigned(1602, 12), 711 => to_unsigned(1455, 12), 712 => to_unsigned(731, 12), 713 => to_unsigned(663, 12), 714 => to_unsigned(2776, 12), 715 => to_unsigned(2547, 12), 716 => to_unsigned(3063, 12), 717 => to_unsigned(311, 12), 718 => to_unsigned(1182, 12), 719 => to_unsigned(1308, 12), 720 => to_unsigned(324, 12), 721 => to_unsigned(676, 12), 722 => to_unsigned(423, 12), 723 => to_unsigned(3676, 12), 724 => to_unsigned(2216, 12), 725 => to_unsigned(3583, 12), 726 => to_unsigned(892, 12), 727 => to_unsigned(1074, 12), 728 => to_unsigned(3898, 12), 729 => to_unsigned(1755, 12), 730 => to_unsigned(810, 12), 731 => to_unsigned(946, 12), 732 => to_unsigned(1079, 12), 733 => to_unsigned(3225, 12), 734 => to_unsigned(2114, 12), 735 => to_unsigned(2777, 12), 736 => to_unsigned(1299, 12), 737 => to_unsigned(201, 12), 738 => to_unsigned(81, 12), 739 => to_unsigned(2987, 12), 740 => to_unsigned(272, 12), 741 => to_unsigned(3061, 12), 742 => to_unsigned(4057, 12), 743 => to_unsigned(3858, 12), 744 => to_unsigned(2870, 12), 745 => to_unsigned(1542, 12), 746 => to_unsigned(3259, 12), 747 => to_unsigned(1357, 12), 748 => to_unsigned(1792, 12), 749 => to_unsigned(2848, 12), 750 => to_unsigned(3327, 12), 751 => to_unsigned(190, 12), 752 => to_unsigned(2411, 12), 753 => to_unsigned(312, 12), 754 => to_unsigned(3323, 12), 755 => to_unsigned(629, 12), 756 => to_unsigned(2814, 12), 757 => to_unsigned(3509, 12), 758 => to_unsigned(2289, 12), 759 => to_unsigned(1573, 12), 760 => to_unsigned(2006, 12), 761 => to_unsigned(2555, 12), 762 => to_unsigned(2152, 12), 763 => to_unsigned(3367, 12), 764 => to_unsigned(3844, 12), 765 => to_unsigned(2498, 12), 766 => to_unsigned(503, 12), 767 => to_unsigned(393, 12), 768 => to_unsigned(1612, 12), 769 => to_unsigned(2140, 12), 770 => to_unsigned(3109, 12), 771 => to_unsigned(3523, 12), 772 => to_unsigned(3154, 12), 773 => to_unsigned(3219, 12), 774 => to_unsigned(3805, 12), 775 => to_unsigned(2241, 12), 776 => to_unsigned(2933, 12), 777 => to_unsigned(944, 12), 778 => to_unsigned(1161, 12), 779 => to_unsigned(463, 12), 780 => to_unsigned(1996, 12), 781 => to_unsigned(3521, 12), 782 => to_unsigned(3626, 12), 783 => to_unsigned(3431, 12), 784 => to_unsigned(3123, 12), 785 => to_unsigned(1300, 12), 786 => to_unsigned(1040, 12), 787 => to_unsigned(1126, 12), 788 => to_unsigned(2950, 12), 789 => to_unsigned(2000, 12), 790 => to_unsigned(2000, 12), 791 => to_unsigned(2602, 12), 792 => to_unsigned(1121, 12), 793 => to_unsigned(2054, 12), 794 => to_unsigned(3738, 12), 795 => to_unsigned(3544, 12), 796 => to_unsigned(186, 12), 797 => to_unsigned(2394, 12), 798 => to_unsigned(2521, 12), 799 => to_unsigned(2961, 12), 800 => to_unsigned(3779, 12), 801 => to_unsigned(1466, 12), 802 => to_unsigned(817, 12), 803 => to_unsigned(158, 12), 804 => to_unsigned(2187, 12), 805 => to_unsigned(3092, 12), 806 => to_unsigned(1957, 12), 807 => to_unsigned(3047, 12), 808 => to_unsigned(826, 12), 809 => to_unsigned(2705, 12), 810 => to_unsigned(3323, 12), 811 => to_unsigned(4070, 12), 812 => to_unsigned(3159, 12), 813 => to_unsigned(730, 12), 814 => to_unsigned(3441, 12), 815 => to_unsigned(895, 12), 816 => to_unsigned(3591, 12), 817 => to_unsigned(4032, 12), 818 => to_unsigned(766, 12), 819 => to_unsigned(1933, 12), 820 => to_unsigned(3020, 12), 821 => to_unsigned(2604, 12), 822 => to_unsigned(533, 12), 823 => to_unsigned(1892, 12), 824 => to_unsigned(664, 12), 825 => to_unsigned(380, 12), 826 => to_unsigned(3373, 12), 827 => to_unsigned(1277, 12), 828 => to_unsigned(324, 12), 829 => to_unsigned(4028, 12), 830 => to_unsigned(3492, 12), 831 => to_unsigned(3497, 12), 832 => to_unsigned(1008, 12), 833 => to_unsigned(826, 12), 834 => to_unsigned(3866, 12), 835 => to_unsigned(929, 12), 836 => to_unsigned(368, 12), 837 => to_unsigned(2507, 12), 838 => to_unsigned(1078, 12), 839 => to_unsigned(2960, 12), 840 => to_unsigned(1255, 12), 841 => to_unsigned(2123, 12), 842 => to_unsigned(1898, 12), 843 => to_unsigned(3949, 12), 844 => to_unsigned(2311, 12), 845 => to_unsigned(861, 12), 846 => to_unsigned(1931, 12), 847 => to_unsigned(160, 12), 848 => to_unsigned(2360, 12), 849 => to_unsigned(60, 12), 850 => to_unsigned(3712, 12), 851 => to_unsigned(3480, 12), 852 => to_unsigned(1508, 12), 853 => to_unsigned(815, 12), 854 => to_unsigned(350, 12), 855 => to_unsigned(378, 12), 856 => to_unsigned(2508, 12), 857 => to_unsigned(3420, 12), 858 => to_unsigned(1638, 12), 859 => to_unsigned(1210, 12), 860 => to_unsigned(1650, 12), 861 => to_unsigned(1887, 12), 862 => to_unsigned(3459, 12), 863 => to_unsigned(2890, 12), 864 => to_unsigned(1992, 12), 865 => to_unsigned(1436, 12), 866 => to_unsigned(4057, 12), 867 => to_unsigned(3182, 12), 868 => to_unsigned(75, 12), 869 => to_unsigned(3002, 12), 870 => to_unsigned(2426, 12), 871 => to_unsigned(68, 12), 872 => to_unsigned(221, 12), 873 => to_unsigned(1819, 12), 874 => to_unsigned(2960, 12), 875 => to_unsigned(3110, 12), 876 => to_unsigned(7, 12), 877 => to_unsigned(1306, 12), 878 => to_unsigned(2225, 12), 879 => to_unsigned(2651, 12), 880 => to_unsigned(4026, 12), 881 => to_unsigned(1073, 12), 882 => to_unsigned(2652, 12), 883 => to_unsigned(3023, 12), 884 => to_unsigned(466, 12), 885 => to_unsigned(1182, 12), 886 => to_unsigned(1075, 12), 887 => to_unsigned(1107, 12), 888 => to_unsigned(2528, 12), 889 => to_unsigned(1593, 12), 890 => to_unsigned(1435, 12), 891 => to_unsigned(3447, 12), 892 => to_unsigned(509, 12), 893 => to_unsigned(3454, 12), 894 => to_unsigned(72, 12), 895 => to_unsigned(388, 12), 896 => to_unsigned(411, 12), 897 => to_unsigned(1575, 12), 898 => to_unsigned(2753, 12), 899 => to_unsigned(3985, 12), 900 => to_unsigned(841, 12), 901 => to_unsigned(437, 12), 902 => to_unsigned(1250, 12), 903 => to_unsigned(726, 12), 904 => to_unsigned(2676, 12), 905 => to_unsigned(2112, 12), 906 => to_unsigned(1756, 12), 907 => to_unsigned(4064, 12), 908 => to_unsigned(3619, 12), 909 => to_unsigned(1058, 12), 910 => to_unsigned(1891, 12), 911 => to_unsigned(1871, 12), 912 => to_unsigned(2097, 12), 913 => to_unsigned(2520, 12), 914 => to_unsigned(3932, 12), 915 => to_unsigned(1910, 12), 916 => to_unsigned(3718, 12), 917 => to_unsigned(1168, 12), 918 => to_unsigned(1480, 12), 919 => to_unsigned(721, 12), 920 => to_unsigned(2489, 12), 921 => to_unsigned(3234, 12), 922 => to_unsigned(1090, 12), 923 => to_unsigned(1800, 12), 924 => to_unsigned(1611, 12), 925 => to_unsigned(104, 12), 926 => to_unsigned(3632, 12), 927 => to_unsigned(1592, 12), 928 => to_unsigned(199, 12), 929 => to_unsigned(1241, 12), 930 => to_unsigned(311, 12), 931 => to_unsigned(724, 12), 932 => to_unsigned(619, 12), 933 => to_unsigned(3238, 12), 934 => to_unsigned(3248, 12), 935 => to_unsigned(1777, 12), 936 => to_unsigned(2297, 12), 937 => to_unsigned(727, 12), 938 => to_unsigned(1122, 12), 939 => to_unsigned(2684, 12), 940 => to_unsigned(996, 12), 941 => to_unsigned(641, 12), 942 => to_unsigned(3184, 12), 943 => to_unsigned(1013, 12), 944 => to_unsigned(2903, 12), 945 => to_unsigned(2033, 12), 946 => to_unsigned(1134, 12), 947 => to_unsigned(3770, 12), 948 => to_unsigned(3972, 12), 949 => to_unsigned(3497, 12), 950 => to_unsigned(1516, 12), 951 => to_unsigned(3597, 12), 952 => to_unsigned(2220, 12), 953 => to_unsigned(2958, 12), 954 => to_unsigned(2786, 12), 955 => to_unsigned(2080, 12), 956 => to_unsigned(1267, 12), 957 => to_unsigned(2736, 12), 958 => to_unsigned(2360, 12), 959 => to_unsigned(1505, 12), 960 => to_unsigned(1808, 12), 961 => to_unsigned(1154, 12), 962 => to_unsigned(3782, 12), 963 => to_unsigned(2452, 12), 964 => to_unsigned(935, 12), 965 => to_unsigned(4095, 12), 966 => to_unsigned(550, 12), 967 => to_unsigned(2690, 12), 968 => to_unsigned(434, 12), 969 => to_unsigned(1417, 12), 970 => to_unsigned(2138, 12), 971 => to_unsigned(3184, 12), 972 => to_unsigned(1598, 12), 973 => to_unsigned(233, 12), 974 => to_unsigned(121, 12), 975 => to_unsigned(1635, 12), 976 => to_unsigned(3239, 12), 977 => to_unsigned(659, 12), 978 => to_unsigned(115, 12), 979 => to_unsigned(1251, 12), 980 => to_unsigned(1996, 12), 981 => to_unsigned(1537, 12), 982 => to_unsigned(1176, 12), 983 => to_unsigned(2011, 12), 984 => to_unsigned(2368, 12), 985 => to_unsigned(3082, 12), 986 => to_unsigned(3619, 12), 987 => to_unsigned(2755, 12), 988 => to_unsigned(1305, 12), 989 => to_unsigned(3227, 12), 990 => to_unsigned(2230, 12), 991 => to_unsigned(1113, 12), 992 => to_unsigned(761, 12), 993 => to_unsigned(1291, 12), 994 => to_unsigned(1232, 12), 995 => to_unsigned(342, 12), 996 => to_unsigned(1727, 12), 997 => to_unsigned(520, 12), 998 => to_unsigned(4066, 12), 999 => to_unsigned(1044, 12), 1000 => to_unsigned(3384, 12), 1001 => to_unsigned(832, 12), 1002 => to_unsigned(477, 12), 1003 => to_unsigned(443, 12), 1004 => to_unsigned(3807, 12), 1005 => to_unsigned(3685, 12), 1006 => to_unsigned(2587, 12), 1007 => to_unsigned(166, 12), 1008 => to_unsigned(1995, 12), 1009 => to_unsigned(1326, 12), 1010 => to_unsigned(3976, 12), 1011 => to_unsigned(2344, 12), 1012 => to_unsigned(3490, 12), 1013 => to_unsigned(3065, 12), 1014 => to_unsigned(1672, 12), 1015 => to_unsigned(3960, 12), 1016 => to_unsigned(1075, 12), 1017 => to_unsigned(3869, 12), 1018 => to_unsigned(99, 12), 1019 => to_unsigned(2749, 12), 1020 => to_unsigned(1239, 12), 1021 => to_unsigned(92, 12), 1022 => to_unsigned(292, 12), 1023 => to_unsigned(1199, 12), 1024 => to_unsigned(2901, 12), 1025 => to_unsigned(1431, 12), 1026 => to_unsigned(1387, 12), 1027 => to_unsigned(926, 12), 1028 => to_unsigned(2597, 12), 1029 => to_unsigned(25, 12), 1030 => to_unsigned(3884, 12), 1031 => to_unsigned(2308, 12), 1032 => to_unsigned(2452, 12), 1033 => to_unsigned(3324, 12), 1034 => to_unsigned(1403, 12), 1035 => to_unsigned(2140, 12), 1036 => to_unsigned(793, 12), 1037 => to_unsigned(836, 12), 1038 => to_unsigned(3279, 12), 1039 => to_unsigned(3970, 12), 1040 => to_unsigned(839, 12), 1041 => to_unsigned(304, 12), 1042 => to_unsigned(450, 12), 1043 => to_unsigned(1247, 12), 1044 => to_unsigned(1690, 12), 1045 => to_unsigned(959, 12), 1046 => to_unsigned(895, 12), 1047 => to_unsigned(774, 12), 1048 => to_unsigned(2050, 12), 1049 => to_unsigned(2923, 12), 1050 => to_unsigned(3437, 12), 1051 => to_unsigned(985, 12), 1052 => to_unsigned(2107, 12), 1053 => to_unsigned(3686, 12), 1054 => to_unsigned(1423, 12), 1055 => to_unsigned(1403, 12), 1056 => to_unsigned(1947, 12), 1057 => to_unsigned(1691, 12), 1058 => to_unsigned(3292, 12), 1059 => to_unsigned(1753, 12), 1060 => to_unsigned(192, 12), 1061 => to_unsigned(1318, 12), 1062 => to_unsigned(1211, 12), 1063 => to_unsigned(3467, 12), 1064 => to_unsigned(277, 12), 1065 => to_unsigned(2822, 12), 1066 => to_unsigned(47, 12), 1067 => to_unsigned(1177, 12), 1068 => to_unsigned(2039, 12), 1069 => to_unsigned(915, 12), 1070 => to_unsigned(3378, 12), 1071 => to_unsigned(259, 12), 1072 => to_unsigned(608, 12), 1073 => to_unsigned(1426, 12), 1074 => to_unsigned(1693, 12), 1075 => to_unsigned(890, 12), 1076 => to_unsigned(1088, 12), 1077 => to_unsigned(2188, 12), 1078 => to_unsigned(44, 12), 1079 => to_unsigned(2275, 12), 1080 => to_unsigned(3816, 12), 1081 => to_unsigned(1336, 12), 1082 => to_unsigned(2123, 12), 1083 => to_unsigned(771, 12), 1084 => to_unsigned(1709, 12), 1085 => to_unsigned(1593, 12), 1086 => to_unsigned(157, 12), 1087 => to_unsigned(3482, 12), 1088 => to_unsigned(2696, 12), 1089 => to_unsigned(3521, 12), 1090 => to_unsigned(961, 12), 1091 => to_unsigned(3060, 12), 1092 => to_unsigned(1606, 12), 1093 => to_unsigned(511, 12), 1094 => to_unsigned(472, 12), 1095 => to_unsigned(3000, 12), 1096 => to_unsigned(2895, 12), 1097 => to_unsigned(1098, 12), 1098 => to_unsigned(1810, 12), 1099 => to_unsigned(628, 12), 1100 => to_unsigned(214, 12), 1101 => to_unsigned(2729, 12), 1102 => to_unsigned(2889, 12), 1103 => to_unsigned(3143, 12), 1104 => to_unsigned(321, 12), 1105 => to_unsigned(1989, 12), 1106 => to_unsigned(3465, 12), 1107 => to_unsigned(1157, 12), 1108 => to_unsigned(1647, 12), 1109 => to_unsigned(687, 12), 1110 => to_unsigned(1780, 12), 1111 => to_unsigned(2100, 12), 1112 => to_unsigned(2239, 12), 1113 => to_unsigned(1966, 12), 1114 => to_unsigned(2003, 12), 1115 => to_unsigned(4011, 12), 1116 => to_unsigned(3164, 12), 1117 => to_unsigned(1960, 12), 1118 => to_unsigned(3693, 12), 1119 => to_unsigned(1234, 12), 1120 => to_unsigned(1611, 12), 1121 => to_unsigned(1222, 12), 1122 => to_unsigned(1202, 12), 1123 => to_unsigned(531, 12), 1124 => to_unsigned(2294, 12), 1125 => to_unsigned(3401, 12), 1126 => to_unsigned(4019, 12), 1127 => to_unsigned(3899, 12), 1128 => to_unsigned(2401, 12), 1129 => to_unsigned(3348, 12), 1130 => to_unsigned(482, 12), 1131 => to_unsigned(4088, 12), 1132 => to_unsigned(332, 12), 1133 => to_unsigned(573, 12), 1134 => to_unsigned(2505, 12), 1135 => to_unsigned(860, 12), 1136 => to_unsigned(3907, 12), 1137 => to_unsigned(2000, 12), 1138 => to_unsigned(2350, 12), 1139 => to_unsigned(3853, 12), 1140 => to_unsigned(2608, 12), 1141 => to_unsigned(3444, 12), 1142 => to_unsigned(1333, 12), 1143 => to_unsigned(3391, 12), 1144 => to_unsigned(174, 12), 1145 => to_unsigned(181, 12), 1146 => to_unsigned(2771, 12), 1147 => to_unsigned(1267, 12), 1148 => to_unsigned(2977, 12), 1149 => to_unsigned(1680, 12), 1150 => to_unsigned(296, 12), 1151 => to_unsigned(1538, 12), 1152 => to_unsigned(3645, 12), 1153 => to_unsigned(399, 12), 1154 => to_unsigned(848, 12), 1155 => to_unsigned(3828, 12), 1156 => to_unsigned(3952, 12), 1157 => to_unsigned(3253, 12), 1158 => to_unsigned(907, 12), 1159 => to_unsigned(133, 12), 1160 => to_unsigned(2239, 12), 1161 => to_unsigned(2516, 12), 1162 => to_unsigned(463, 12), 1163 => to_unsigned(1085, 12), 1164 => to_unsigned(2701, 12), 1165 => to_unsigned(3099, 12), 1166 => to_unsigned(3222, 12), 1167 => to_unsigned(3198, 12), 1168 => to_unsigned(3834, 12), 1169 => to_unsigned(3414, 12), 1170 => to_unsigned(1735, 12), 1171 => to_unsigned(1066, 12), 1172 => to_unsigned(3735, 12), 1173 => to_unsigned(1496, 12), 1174 => to_unsigned(3937, 12), 1175 => to_unsigned(854, 12), 1176 => to_unsigned(2278, 12), 1177 => to_unsigned(900, 12), 1178 => to_unsigned(3939, 12), 1179 => to_unsigned(2085, 12), 1180 => to_unsigned(2660, 12), 1181 => to_unsigned(673, 12), 1182 => to_unsigned(3702, 12), 1183 => to_unsigned(1140, 12), 1184 => to_unsigned(2989, 12), 1185 => to_unsigned(3624, 12), 1186 => to_unsigned(2084, 12), 1187 => to_unsigned(1557, 12), 1188 => to_unsigned(2908, 12), 1189 => to_unsigned(1064, 12), 1190 => to_unsigned(2108, 12), 1191 => to_unsigned(3034, 12), 1192 => to_unsigned(1157, 12), 1193 => to_unsigned(465, 12), 1194 => to_unsigned(1227, 12), 1195 => to_unsigned(773, 12), 1196 => to_unsigned(4055, 12), 1197 => to_unsigned(2991, 12), 1198 => to_unsigned(1379, 12), 1199 => to_unsigned(1653, 12), 1200 => to_unsigned(797, 12), 1201 => to_unsigned(513, 12), 1202 => to_unsigned(2228, 12), 1203 => to_unsigned(665, 12), 1204 => to_unsigned(55, 12), 1205 => to_unsigned(2212, 12), 1206 => to_unsigned(1751, 12), 1207 => to_unsigned(3418, 12), 1208 => to_unsigned(1794, 12), 1209 => to_unsigned(3097, 12), 1210 => to_unsigned(2124, 12), 1211 => to_unsigned(1978, 12), 1212 => to_unsigned(1972, 12), 1213 => to_unsigned(2682, 12), 1214 => to_unsigned(52, 12), 1215 => to_unsigned(3606, 12), 1216 => to_unsigned(331, 12), 1217 => to_unsigned(3447, 12), 1218 => to_unsigned(2913, 12), 1219 => to_unsigned(2615, 12), 1220 => to_unsigned(2069, 12), 1221 => to_unsigned(1466, 12), 1222 => to_unsigned(3489, 12), 1223 => to_unsigned(3174, 12), 1224 => to_unsigned(951, 12), 1225 => to_unsigned(1722, 12), 1226 => to_unsigned(2904, 12), 1227 => to_unsigned(3490, 12), 1228 => to_unsigned(2312, 12), 1229 => to_unsigned(3134, 12), 1230 => to_unsigned(3976, 12), 1231 => to_unsigned(4006, 12), 1232 => to_unsigned(96, 12), 1233 => to_unsigned(2765, 12), 1234 => to_unsigned(1315, 12), 1235 => to_unsigned(1182, 12), 1236 => to_unsigned(127, 12), 1237 => to_unsigned(359, 12), 1238 => to_unsigned(1662, 12), 1239 => to_unsigned(1008, 12), 1240 => to_unsigned(4041, 12), 1241 => to_unsigned(1405, 12), 1242 => to_unsigned(2413, 12), 1243 => to_unsigned(1428, 12), 1244 => to_unsigned(720, 12), 1245 => to_unsigned(271, 12), 1246 => to_unsigned(1893, 12), 1247 => to_unsigned(3160, 12), 1248 => to_unsigned(179, 12), 1249 => to_unsigned(477, 12), 1250 => to_unsigned(1515, 12), 1251 => to_unsigned(464, 12), 1252 => to_unsigned(1290, 12), 1253 => to_unsigned(2116, 12), 1254 => to_unsigned(3220, 12), 1255 => to_unsigned(3544, 12), 1256 => to_unsigned(1751, 12), 1257 => to_unsigned(1581, 12), 1258 => to_unsigned(2660, 12), 1259 => to_unsigned(2165, 12), 1260 => to_unsigned(510, 12), 1261 => to_unsigned(1437, 12), 1262 => to_unsigned(811, 12), 1263 => to_unsigned(179, 12), 1264 => to_unsigned(3477, 12), 1265 => to_unsigned(2890, 12), 1266 => to_unsigned(106, 12), 1267 => to_unsigned(1913, 12), 1268 => to_unsigned(642, 12), 1269 => to_unsigned(2373, 12), 1270 => to_unsigned(3565, 12), 1271 => to_unsigned(3784, 12), 1272 => to_unsigned(3222, 12), 1273 => to_unsigned(1250, 12), 1274 => to_unsigned(228, 12), 1275 => to_unsigned(2605, 12), 1276 => to_unsigned(3296, 12), 1277 => to_unsigned(1067, 12), 1278 => to_unsigned(3194, 12), 1279 => to_unsigned(1731, 12), 1280 => to_unsigned(30, 12), 1281 => to_unsigned(3114, 12), 1282 => to_unsigned(1964, 12), 1283 => to_unsigned(1654, 12), 1284 => to_unsigned(2465, 12), 1285 => to_unsigned(2351, 12), 1286 => to_unsigned(2787, 12), 1287 => to_unsigned(49, 12), 1288 => to_unsigned(289, 12), 1289 => to_unsigned(356, 12), 1290 => to_unsigned(3624, 12), 1291 => to_unsigned(1929, 12), 1292 => to_unsigned(1025, 12), 1293 => to_unsigned(1405, 12), 1294 => to_unsigned(3119, 12), 1295 => to_unsigned(3604, 12), 1296 => to_unsigned(902, 12), 1297 => to_unsigned(2763, 12), 1298 => to_unsigned(2811, 12), 1299 => to_unsigned(419, 12), 1300 => to_unsigned(292, 12), 1301 => to_unsigned(3457, 12), 1302 => to_unsigned(4011, 12), 1303 => to_unsigned(1093, 12), 1304 => to_unsigned(2807, 12), 1305 => to_unsigned(190, 12), 1306 => to_unsigned(2131, 12), 1307 => to_unsigned(3813, 12), 1308 => to_unsigned(1883, 12), 1309 => to_unsigned(2918, 12), 1310 => to_unsigned(1531, 12), 1311 => to_unsigned(770, 12), 1312 => to_unsigned(1177, 12), 1313 => to_unsigned(3777, 12), 1314 => to_unsigned(961, 12), 1315 => to_unsigned(1912, 12), 1316 => to_unsigned(3597, 12), 1317 => to_unsigned(588, 12), 1318 => to_unsigned(2359, 12), 1319 => to_unsigned(633, 12), 1320 => to_unsigned(3211, 12), 1321 => to_unsigned(3219, 12), 1322 => to_unsigned(2771, 12), 1323 => to_unsigned(1792, 12), 1324 => to_unsigned(3326, 12), 1325 => to_unsigned(3889, 12), 1326 => to_unsigned(1195, 12), 1327 => to_unsigned(1680, 12), 1328 => to_unsigned(161, 12), 1329 => to_unsigned(3817, 12), 1330 => to_unsigned(467, 12), 1331 => to_unsigned(281, 12), 1332 => to_unsigned(2499, 12), 1333 => to_unsigned(1986, 12), 1334 => to_unsigned(2950, 12), 1335 => to_unsigned(3507, 12), 1336 => to_unsigned(3657, 12), 1337 => to_unsigned(1664, 12), 1338 => to_unsigned(975, 12), 1339 => to_unsigned(2031, 12), 1340 => to_unsigned(2151, 12), 1341 => to_unsigned(1222, 12), 1342 => to_unsigned(542, 12), 1343 => to_unsigned(787, 12), 1344 => to_unsigned(1298, 12), 1345 => to_unsigned(1510, 12), 1346 => to_unsigned(2369, 12), 1347 => to_unsigned(3797, 12), 1348 => to_unsigned(1182, 12), 1349 => to_unsigned(3688, 12), 1350 => to_unsigned(674, 12), 1351 => to_unsigned(785, 12), 1352 => to_unsigned(2152, 12), 1353 => to_unsigned(1664, 12), 1354 => to_unsigned(981, 12), 1355 => to_unsigned(413, 12), 1356 => to_unsigned(2226, 12), 1357 => to_unsigned(512, 12), 1358 => to_unsigned(157, 12), 1359 => to_unsigned(2915, 12), 1360 => to_unsigned(1152, 12), 1361 => to_unsigned(1981, 12), 1362 => to_unsigned(2685, 12), 1363 => to_unsigned(2150, 12), 1364 => to_unsigned(462, 12), 1365 => to_unsigned(248, 12), 1366 => to_unsigned(483, 12), 1367 => to_unsigned(1972, 12), 1368 => to_unsigned(86, 12), 1369 => to_unsigned(2836, 12), 1370 => to_unsigned(3504, 12), 1371 => to_unsigned(2845, 12), 1372 => to_unsigned(3964, 12), 1373 => to_unsigned(3470, 12), 1374 => to_unsigned(818, 12), 1375 => to_unsigned(2279, 12), 1376 => to_unsigned(724, 12), 1377 => to_unsigned(2327, 12), 1378 => to_unsigned(419, 12), 1379 => to_unsigned(1228, 12), 1380 => to_unsigned(2219, 12), 1381 => to_unsigned(2665, 12), 1382 => to_unsigned(2741, 12), 1383 => to_unsigned(3229, 12), 1384 => to_unsigned(258, 12), 1385 => to_unsigned(2737, 12), 1386 => to_unsigned(326, 12), 1387 => to_unsigned(56, 12), 1388 => to_unsigned(3121, 12), 1389 => to_unsigned(2047, 12), 1390 => to_unsigned(2534, 12), 1391 => to_unsigned(1469, 12), 1392 => to_unsigned(1325, 12), 1393 => to_unsigned(819, 12), 1394 => to_unsigned(116, 12), 1395 => to_unsigned(30, 12), 1396 => to_unsigned(3379, 12), 1397 => to_unsigned(1401, 12), 1398 => to_unsigned(2214, 12), 1399 => to_unsigned(2308, 12), 1400 => to_unsigned(2849, 12), 1401 => to_unsigned(2684, 12), 1402 => to_unsigned(383, 12), 1403 => to_unsigned(623, 12), 1404 => to_unsigned(2076, 12), 1405 => to_unsigned(4030, 12), 1406 => to_unsigned(4056, 12), 1407 => to_unsigned(3113, 12), 1408 => to_unsigned(1591, 12), 1409 => to_unsigned(3056, 12), 1410 => to_unsigned(1475, 12), 1411 => to_unsigned(1681, 12), 1412 => to_unsigned(3757, 12), 1413 => to_unsigned(1797, 12), 1414 => to_unsigned(2017, 12), 1415 => to_unsigned(458, 12), 1416 => to_unsigned(1024, 12), 1417 => to_unsigned(545, 12), 1418 => to_unsigned(338, 12), 1419 => to_unsigned(834, 12), 1420 => to_unsigned(3181, 12), 1421 => to_unsigned(2051, 12), 1422 => to_unsigned(2559, 12), 1423 => to_unsigned(3219, 12), 1424 => to_unsigned(1115, 12), 1425 => to_unsigned(3954, 12), 1426 => to_unsigned(1386, 12), 1427 => to_unsigned(2578, 12), 1428 => to_unsigned(680, 12), 1429 => to_unsigned(2267, 12), 1430 => to_unsigned(954, 12), 1431 => to_unsigned(1785, 12), 1432 => to_unsigned(1412, 12), 1433 => to_unsigned(3340, 12), 1434 => to_unsigned(3729, 12), 1435 => to_unsigned(3093, 12), 1436 => to_unsigned(3507, 12), 1437 => to_unsigned(1502, 12), 1438 => to_unsigned(1142, 12), 1439 => to_unsigned(2662, 12), 1440 => to_unsigned(4073, 12), 1441 => to_unsigned(2058, 12), 1442 => to_unsigned(3171, 12), 1443 => to_unsigned(2617, 12), 1444 => to_unsigned(3497, 12), 1445 => to_unsigned(1212, 12), 1446 => to_unsigned(2964, 12), 1447 => to_unsigned(2645, 12), 1448 => to_unsigned(840, 12), 1449 => to_unsigned(2994, 12), 1450 => to_unsigned(1273, 12), 1451 => to_unsigned(2449, 12), 1452 => to_unsigned(3333, 12), 1453 => to_unsigned(526, 12), 1454 => to_unsigned(3236, 12), 1455 => to_unsigned(2257, 12), 1456 => to_unsigned(485, 12), 1457 => to_unsigned(3607, 12), 1458 => to_unsigned(3511, 12), 1459 => to_unsigned(662, 12), 1460 => to_unsigned(2397, 12), 1461 => to_unsigned(3345, 12), 1462 => to_unsigned(2515, 12), 1463 => to_unsigned(3847, 12), 1464 => to_unsigned(641, 12), 1465 => to_unsigned(3631, 12), 1466 => to_unsigned(2646, 12), 1467 => to_unsigned(649, 12), 1468 => to_unsigned(2824, 12), 1469 => to_unsigned(339, 12), 1470 => to_unsigned(1343, 12), 1471 => to_unsigned(2796, 12), 1472 => to_unsigned(3993, 12), 1473 => to_unsigned(2867, 12), 1474 => to_unsigned(1493, 12), 1475 => to_unsigned(3354, 12), 1476 => to_unsigned(3455, 12), 1477 => to_unsigned(3723, 12), 1478 => to_unsigned(3561, 12), 1479 => to_unsigned(1038, 12), 1480 => to_unsigned(1053, 12), 1481 => to_unsigned(1586, 12), 1482 => to_unsigned(1657, 12), 1483 => to_unsigned(246, 12), 1484 => to_unsigned(1068, 12), 1485 => to_unsigned(3194, 12), 1486 => to_unsigned(2130, 12), 1487 => to_unsigned(3550, 12), 1488 => to_unsigned(3303, 12), 1489 => to_unsigned(3553, 12), 1490 => to_unsigned(2068, 12), 1491 => to_unsigned(2082, 12), 1492 => to_unsigned(2850, 12), 1493 => to_unsigned(374, 12), 1494 => to_unsigned(3230, 12), 1495 => to_unsigned(559, 12), 1496 => to_unsigned(2493, 12), 1497 => to_unsigned(2163, 12), 1498 => to_unsigned(3834, 12), 1499 => to_unsigned(3541, 12), 1500 => to_unsigned(2020, 12), 1501 => to_unsigned(3973, 12), 1502 => to_unsigned(3655, 12), 1503 => to_unsigned(3008, 12), 1504 => to_unsigned(225, 12), 1505 => to_unsigned(1068, 12), 1506 => to_unsigned(1288, 12), 1507 => to_unsigned(3908, 12), 1508 => to_unsigned(3497, 12), 1509 => to_unsigned(1557, 12), 1510 => to_unsigned(3090, 12), 1511 => to_unsigned(765, 12), 1512 => to_unsigned(2795, 12), 1513 => to_unsigned(3681, 12), 1514 => to_unsigned(1955, 12), 1515 => to_unsigned(919, 12), 1516 => to_unsigned(2783, 12), 1517 => to_unsigned(3925, 12), 1518 => to_unsigned(3626, 12), 1519 => to_unsigned(3066, 12), 1520 => to_unsigned(301, 12), 1521 => to_unsigned(2256, 12), 1522 => to_unsigned(3644, 12), 1523 => to_unsigned(1752, 12), 1524 => to_unsigned(3294, 12), 1525 => to_unsigned(3255, 12), 1526 => to_unsigned(972, 12), 1527 => to_unsigned(2610, 12), 1528 => to_unsigned(2628, 12), 1529 => to_unsigned(2676, 12), 1530 => to_unsigned(2457, 12), 1531 => to_unsigned(3607, 12), 1532 => to_unsigned(525, 12), 1533 => to_unsigned(1284, 12), 1534 => to_unsigned(987, 12), 1535 => to_unsigned(3888, 12), 1536 => to_unsigned(1718, 12), 1537 => to_unsigned(2479, 12), 1538 => to_unsigned(1450, 12), 1539 => to_unsigned(3891, 12), 1540 => to_unsigned(434, 12), 1541 => to_unsigned(884, 12), 1542 => to_unsigned(2879, 12), 1543 => to_unsigned(2613, 12), 1544 => to_unsigned(1865, 12), 1545 => to_unsigned(1432, 12), 1546 => to_unsigned(684, 12), 1547 => to_unsigned(2215, 12), 1548 => to_unsigned(2119, 12), 1549 => to_unsigned(2169, 12), 1550 => to_unsigned(2038, 12), 1551 => to_unsigned(167, 12), 1552 => to_unsigned(3202, 12), 1553 => to_unsigned(3094, 12), 1554 => to_unsigned(2963, 12), 1555 => to_unsigned(1109, 12), 1556 => to_unsigned(3156, 12), 1557 => to_unsigned(1232, 12), 1558 => to_unsigned(655, 12), 1559 => to_unsigned(3938, 12), 1560 => to_unsigned(2242, 12), 1561 => to_unsigned(2149, 12), 1562 => to_unsigned(204, 12), 1563 => to_unsigned(58, 12), 1564 => to_unsigned(663, 12), 1565 => to_unsigned(3596, 12), 1566 => to_unsigned(3491, 12), 1567 => to_unsigned(2023, 12), 1568 => to_unsigned(493, 12), 1569 => to_unsigned(1086, 12), 1570 => to_unsigned(460, 12), 1571 => to_unsigned(3491, 12), 1572 => to_unsigned(554, 12), 1573 => to_unsigned(827, 12), 1574 => to_unsigned(757, 12), 1575 => to_unsigned(475, 12), 1576 => to_unsigned(3747, 12), 1577 => to_unsigned(2873, 12), 1578 => to_unsigned(3028, 12), 1579 => to_unsigned(562, 12), 1580 => to_unsigned(3882, 12), 1581 => to_unsigned(2223, 12), 1582 => to_unsigned(2396, 12), 1583 => to_unsigned(364, 12), 1584 => to_unsigned(3657, 12), 1585 => to_unsigned(3244, 12), 1586 => to_unsigned(2972, 12), 1587 => to_unsigned(1323, 12), 1588 => to_unsigned(2362, 12), 1589 => to_unsigned(1501, 12), 1590 => to_unsigned(172, 12), 1591 => to_unsigned(86, 12), 1592 => to_unsigned(1628, 12), 1593 => to_unsigned(1708, 12), 1594 => to_unsigned(4071, 12), 1595 => to_unsigned(2611, 12), 1596 => to_unsigned(924, 12), 1597 => to_unsigned(3747, 12), 1598 => to_unsigned(1286, 12), 1599 => to_unsigned(106, 12), 1600 => to_unsigned(614, 12), 1601 => to_unsigned(297, 12), 1602 => to_unsigned(2982, 12), 1603 => to_unsigned(2539, 12), 1604 => to_unsigned(44, 12), 1605 => to_unsigned(242, 12), 1606 => to_unsigned(691, 12), 1607 => to_unsigned(3108, 12), 1608 => to_unsigned(1408, 12), 1609 => to_unsigned(1088, 12), 1610 => to_unsigned(111, 12), 1611 => to_unsigned(697, 12), 1612 => to_unsigned(783, 12), 1613 => to_unsigned(3972, 12), 1614 => to_unsigned(303, 12), 1615 => to_unsigned(3130, 12), 1616 => to_unsigned(734, 12), 1617 => to_unsigned(109, 12), 1618 => to_unsigned(1823, 12), 1619 => to_unsigned(2451, 12), 1620 => to_unsigned(1458, 12), 1621 => to_unsigned(2273, 12), 1622 => to_unsigned(211, 12), 1623 => to_unsigned(3989, 12), 1624 => to_unsigned(121, 12), 1625 => to_unsigned(4062, 12), 1626 => to_unsigned(3421, 12), 1627 => to_unsigned(2046, 12), 1628 => to_unsigned(2266, 12), 1629 => to_unsigned(1504, 12), 1630 => to_unsigned(2896, 12), 1631 => to_unsigned(1167, 12), 1632 => to_unsigned(2404, 12), 1633 => to_unsigned(1295, 12), 1634 => to_unsigned(1542, 12), 1635 => to_unsigned(798, 12), 1636 => to_unsigned(1211, 12), 1637 => to_unsigned(1529, 12), 1638 => to_unsigned(1199, 12), 1639 => to_unsigned(2068, 12), 1640 => to_unsigned(3293, 12), 1641 => to_unsigned(2408, 12), 1642 => to_unsigned(533, 12), 1643 => to_unsigned(316, 12), 1644 => to_unsigned(1695, 12), 1645 => to_unsigned(323, 12), 1646 => to_unsigned(1411, 12), 1647 => to_unsigned(2045, 12), 1648 => to_unsigned(772, 12), 1649 => to_unsigned(3309, 12), 1650 => to_unsigned(660, 12), 1651 => to_unsigned(1853, 12), 1652 => to_unsigned(3522, 12), 1653 => to_unsigned(395, 12), 1654 => to_unsigned(524, 12), 1655 => to_unsigned(4005, 12), 1656 => to_unsigned(3848, 12), 1657 => to_unsigned(3030, 12), 1658 => to_unsigned(1963, 12), 1659 => to_unsigned(1192, 12), 1660 => to_unsigned(3383, 12), 1661 => to_unsigned(2700, 12), 1662 => to_unsigned(3711, 12), 1663 => to_unsigned(4058, 12), 1664 => to_unsigned(346, 12), 1665 => to_unsigned(116, 12), 1666 => to_unsigned(3025, 12), 1667 => to_unsigned(2983, 12), 1668 => to_unsigned(2743, 12), 1669 => to_unsigned(3198, 12), 1670 => to_unsigned(3843, 12), 1671 => to_unsigned(2181, 12), 1672 => to_unsigned(2839, 12), 1673 => to_unsigned(304, 12), 1674 => to_unsigned(2221, 12), 1675 => to_unsigned(3047, 12), 1676 => to_unsigned(4009, 12), 1677 => to_unsigned(1962, 12), 1678 => to_unsigned(691, 12), 1679 => to_unsigned(814, 12), 1680 => to_unsigned(1717, 12), 1681 => to_unsigned(612, 12), 1682 => to_unsigned(74, 12), 1683 => to_unsigned(372, 12), 1684 => to_unsigned(3780, 12), 1685 => to_unsigned(1239, 12), 1686 => to_unsigned(3920, 12), 1687 => to_unsigned(2806, 12), 1688 => to_unsigned(1213, 12), 1689 => to_unsigned(3725, 12), 1690 => to_unsigned(3756, 12), 1691 => to_unsigned(2351, 12), 1692 => to_unsigned(2051, 12), 1693 => to_unsigned(1498, 12), 1694 => to_unsigned(674, 12), 1695 => to_unsigned(368, 12), 1696 => to_unsigned(1395, 12), 1697 => to_unsigned(3690, 12), 1698 => to_unsigned(684, 12), 1699 => to_unsigned(2818, 12), 1700 => to_unsigned(77, 12), 1701 => to_unsigned(2262, 12), 1702 => to_unsigned(2828, 12), 1703 => to_unsigned(521, 12), 1704 => to_unsigned(3664, 12), 1705 => to_unsigned(643, 12), 1706 => to_unsigned(3264, 12), 1707 => to_unsigned(313, 12), 1708 => to_unsigned(524, 12), 1709 => to_unsigned(4002, 12), 1710 => to_unsigned(1340, 12), 1711 => to_unsigned(640, 12), 1712 => to_unsigned(2069, 12), 1713 => to_unsigned(924, 12), 1714 => to_unsigned(503, 12), 1715 => to_unsigned(1217, 12), 1716 => to_unsigned(2458, 12), 1717 => to_unsigned(2496, 12), 1718 => to_unsigned(1749, 12), 1719 => to_unsigned(2582, 12), 1720 => to_unsigned(115, 12), 1721 => to_unsigned(1442, 12), 1722 => to_unsigned(3050, 12), 1723 => to_unsigned(1505, 12), 1724 => to_unsigned(345, 12), 1725 => to_unsigned(1863, 12), 1726 => to_unsigned(2315, 12), 1727 => to_unsigned(2285, 12), 1728 => to_unsigned(1749, 12), 1729 => to_unsigned(1014, 12), 1730 => to_unsigned(598, 12), 1731 => to_unsigned(3975, 12), 1732 => to_unsigned(417, 12), 1733 => to_unsigned(2203, 12), 1734 => to_unsigned(953, 12), 1735 => to_unsigned(1479, 12), 1736 => to_unsigned(3558, 12), 1737 => to_unsigned(454, 12), 1738 => to_unsigned(1512, 12), 1739 => to_unsigned(3993, 12), 1740 => to_unsigned(1283, 12), 1741 => to_unsigned(3976, 12), 1742 => to_unsigned(2477, 12), 1743 => to_unsigned(3662, 12), 1744 => to_unsigned(3026, 12), 1745 => to_unsigned(2619, 12), 1746 => to_unsigned(3911, 12), 1747 => to_unsigned(2623, 12), 1748 => to_unsigned(658, 12), 1749 => to_unsigned(1299, 12), 1750 => to_unsigned(2470, 12), 1751 => to_unsigned(3709, 12), 1752 => to_unsigned(414, 12), 1753 => to_unsigned(2190, 12), 1754 => to_unsigned(247, 12), 1755 => to_unsigned(2447, 12), 1756 => to_unsigned(2372, 12), 1757 => to_unsigned(2782, 12), 1758 => to_unsigned(2786, 12), 1759 => to_unsigned(2416, 12), 1760 => to_unsigned(139, 12), 1761 => to_unsigned(2129, 12), 1762 => to_unsigned(3439, 12), 1763 => to_unsigned(1269, 12), 1764 => to_unsigned(585, 12), 1765 => to_unsigned(2277, 12), 1766 => to_unsigned(1441, 12), 1767 => to_unsigned(3277, 12), 1768 => to_unsigned(2469, 12), 1769 => to_unsigned(2001, 12), 1770 => to_unsigned(3236, 12), 1771 => to_unsigned(285, 12), 1772 => to_unsigned(1074, 12), 1773 => to_unsigned(171, 12), 1774 => to_unsigned(2558, 12), 1775 => to_unsigned(3480, 12), 1776 => to_unsigned(3958, 12), 1777 => to_unsigned(1722, 12), 1778 => to_unsigned(1511, 12), 1779 => to_unsigned(3713, 12), 1780 => to_unsigned(499, 12), 1781 => to_unsigned(611, 12), 1782 => to_unsigned(1382, 12), 1783 => to_unsigned(183, 12), 1784 => to_unsigned(1724, 12), 1785 => to_unsigned(1905, 12), 1786 => to_unsigned(511, 12), 1787 => to_unsigned(2480, 12), 1788 => to_unsigned(3499, 12), 1789 => to_unsigned(618, 12), 1790 => to_unsigned(818, 12), 1791 => to_unsigned(3169, 12), 1792 => to_unsigned(2850, 12), 1793 => to_unsigned(486, 12), 1794 => to_unsigned(863, 12), 1795 => to_unsigned(2555, 12), 1796 => to_unsigned(2758, 12), 1797 => to_unsigned(92, 12), 1798 => to_unsigned(1196, 12), 1799 => to_unsigned(3315, 12), 1800 => to_unsigned(2381, 12), 1801 => to_unsigned(3060, 12), 1802 => to_unsigned(1197, 12), 1803 => to_unsigned(104, 12), 1804 => to_unsigned(1621, 12), 1805 => to_unsigned(4025, 12), 1806 => to_unsigned(3796, 12), 1807 => to_unsigned(594, 12), 1808 => to_unsigned(2239, 12), 1809 => to_unsigned(3415, 12), 1810 => to_unsigned(4, 12), 1811 => to_unsigned(2651, 12), 1812 => to_unsigned(280, 12), 1813 => to_unsigned(1804, 12), 1814 => to_unsigned(1949, 12), 1815 => to_unsigned(3036, 12), 1816 => to_unsigned(3734, 12), 1817 => to_unsigned(3017, 12), 1818 => to_unsigned(101, 12), 1819 => to_unsigned(402, 12), 1820 => to_unsigned(34, 12), 1821 => to_unsigned(1551, 12), 1822 => to_unsigned(3930, 12), 1823 => to_unsigned(2059, 12), 1824 => to_unsigned(1041, 12), 1825 => to_unsigned(3740, 12), 1826 => to_unsigned(3117, 12), 1827 => to_unsigned(2451, 12), 1828 => to_unsigned(1360, 12), 1829 => to_unsigned(1682, 12), 1830 => to_unsigned(884, 12), 1831 => to_unsigned(3571, 12), 1832 => to_unsigned(3576, 12), 1833 => to_unsigned(2520, 12), 1834 => to_unsigned(5, 12), 1835 => to_unsigned(3258, 12), 1836 => to_unsigned(2129, 12), 1837 => to_unsigned(58, 12), 1838 => to_unsigned(1838, 12), 1839 => to_unsigned(1149, 12), 1840 => to_unsigned(3483, 12), 1841 => to_unsigned(1616, 12), 1842 => to_unsigned(725, 12), 1843 => to_unsigned(1118, 12), 1844 => to_unsigned(1911, 12), 1845 => to_unsigned(3900, 12), 1846 => to_unsigned(1900, 12), 1847 => to_unsigned(897, 12), 1848 => to_unsigned(2691, 12), 1849 => to_unsigned(3304, 12), 1850 => to_unsigned(2992, 12), 1851 => to_unsigned(2239, 12), 1852 => to_unsigned(4040, 12), 1853 => to_unsigned(1372, 12), 1854 => to_unsigned(526, 12), 1855 => to_unsigned(750, 12), 1856 => to_unsigned(3429, 12), 1857 => to_unsigned(3408, 12), 1858 => to_unsigned(3721, 12), 1859 => to_unsigned(182, 12), 1860 => to_unsigned(1281, 12), 1861 => to_unsigned(1493, 12), 1862 => to_unsigned(3079, 12), 1863 => to_unsigned(776, 12), 1864 => to_unsigned(1974, 12), 1865 => to_unsigned(537, 12), 1866 => to_unsigned(3801, 12), 1867 => to_unsigned(930, 12), 1868 => to_unsigned(1865, 12), 1869 => to_unsigned(2363, 12), 1870 => to_unsigned(739, 12), 1871 => to_unsigned(280, 12), 1872 => to_unsigned(1006, 12), 1873 => to_unsigned(1689, 12), 1874 => to_unsigned(61, 12), 1875 => to_unsigned(1345, 12), 1876 => to_unsigned(902, 12), 1877 => to_unsigned(1489, 12), 1878 => to_unsigned(740, 12), 1879 => to_unsigned(474, 12), 1880 => to_unsigned(3046, 12), 1881 => to_unsigned(1660, 12), 1882 => to_unsigned(816, 12), 1883 => to_unsigned(203, 12), 1884 => to_unsigned(2502, 12), 1885 => to_unsigned(2434, 12), 1886 => to_unsigned(3595, 12), 1887 => to_unsigned(867, 12), 1888 => to_unsigned(533, 12), 1889 => to_unsigned(365, 12), 1890 => to_unsigned(2636, 12), 1891 => to_unsigned(2033, 12), 1892 => to_unsigned(722, 12), 1893 => to_unsigned(4012, 12), 1894 => to_unsigned(2878, 12), 1895 => to_unsigned(3287, 12), 1896 => to_unsigned(2728, 12), 1897 => to_unsigned(3781, 12), 1898 => to_unsigned(3799, 12), 1899 => to_unsigned(4042, 12), 1900 => to_unsigned(1986, 12), 1901 => to_unsigned(813, 12), 1902 => to_unsigned(392, 12), 1903 => to_unsigned(3898, 12), 1904 => to_unsigned(3550, 12), 1905 => to_unsigned(3279, 12), 1906 => to_unsigned(3902, 12), 1907 => to_unsigned(1387, 12), 1908 => to_unsigned(1383, 12), 1909 => to_unsigned(2230, 12), 1910 => to_unsigned(956, 12), 1911 => to_unsigned(2776, 12), 1912 => to_unsigned(1984, 12), 1913 => to_unsigned(3379, 12), 1914 => to_unsigned(1121, 12), 1915 => to_unsigned(213, 12), 1916 => to_unsigned(3502, 12), 1917 => to_unsigned(1072, 12), 1918 => to_unsigned(1712, 12), 1919 => to_unsigned(2026, 12), 1920 => to_unsigned(1269, 12), 1921 => to_unsigned(1642, 12), 1922 => to_unsigned(1703, 12), 1923 => to_unsigned(2339, 12), 1924 => to_unsigned(1373, 12), 1925 => to_unsigned(358, 12), 1926 => to_unsigned(1516, 12), 1927 => to_unsigned(469, 12), 1928 => to_unsigned(2713, 12), 1929 => to_unsigned(1317, 12), 1930 => to_unsigned(2828, 12), 1931 => to_unsigned(1337, 12), 1932 => to_unsigned(1301, 12), 1933 => to_unsigned(3096, 12), 1934 => to_unsigned(2839, 12), 1935 => to_unsigned(34, 12), 1936 => to_unsigned(3829, 12), 1937 => to_unsigned(1581, 12), 1938 => to_unsigned(1887, 12), 1939 => to_unsigned(4076, 12), 1940 => to_unsigned(2558, 12), 1941 => to_unsigned(3061, 12), 1942 => to_unsigned(324, 12), 1943 => to_unsigned(3391, 12), 1944 => to_unsigned(1021, 12), 1945 => to_unsigned(2785, 12), 1946 => to_unsigned(3014, 12), 1947 => to_unsigned(1774, 12), 1948 => to_unsigned(2207, 12), 1949 => to_unsigned(3738, 12), 1950 => to_unsigned(2616, 12), 1951 => to_unsigned(1788, 12), 1952 => to_unsigned(3028, 12), 1953 => to_unsigned(2016, 12), 1954 => to_unsigned(2118, 12), 1955 => to_unsigned(1923, 12), 1956 => to_unsigned(336, 12), 1957 => to_unsigned(946, 12), 1958 => to_unsigned(750, 12), 1959 => to_unsigned(3704, 12), 1960 => to_unsigned(254, 12), 1961 => to_unsigned(2430, 12), 1962 => to_unsigned(2111, 12), 1963 => to_unsigned(3320, 12), 1964 => to_unsigned(2136, 12), 1965 => to_unsigned(646, 12), 1966 => to_unsigned(2078, 12), 1967 => to_unsigned(3969, 12), 1968 => to_unsigned(1761, 12), 1969 => to_unsigned(4075, 12), 1970 => to_unsigned(383, 12), 1971 => to_unsigned(696, 12), 1972 => to_unsigned(1030, 12), 1973 => to_unsigned(1560, 12), 1974 => to_unsigned(160, 12), 1975 => to_unsigned(1607, 12), 1976 => to_unsigned(3178, 12), 1977 => to_unsigned(3970, 12), 1978 => to_unsigned(970, 12), 1979 => to_unsigned(305, 12), 1980 => to_unsigned(3905, 12), 1981 => to_unsigned(98, 12), 1982 => to_unsigned(66, 12), 1983 => to_unsigned(2015, 12), 1984 => to_unsigned(1694, 12), 1985 => to_unsigned(2619, 12), 1986 => to_unsigned(2338, 12), 1987 => to_unsigned(2990, 12), 1988 => to_unsigned(861, 12), 1989 => to_unsigned(3530, 12), 1990 => to_unsigned(61, 12), 1991 => to_unsigned(1100, 12), 1992 => to_unsigned(3993, 12), 1993 => to_unsigned(2132, 12), 1994 => to_unsigned(2998, 12), 1995 => to_unsigned(3720, 12), 1996 => to_unsigned(2760, 12), 1997 => to_unsigned(1694, 12), 1998 => to_unsigned(507, 12), 1999 => to_unsigned(2790, 12), 2000 => to_unsigned(2633, 12), 2001 => to_unsigned(1381, 12), 2002 => to_unsigned(504, 12), 2003 => to_unsigned(2003, 12), 2004 => to_unsigned(1039, 12), 2005 => to_unsigned(1108, 12), 2006 => to_unsigned(1871, 12), 2007 => to_unsigned(1401, 12), 2008 => to_unsigned(3854, 12), 2009 => to_unsigned(2815, 12), 2010 => to_unsigned(242, 12), 2011 => to_unsigned(915, 12), 2012 => to_unsigned(4077, 12), 2013 => to_unsigned(626, 12), 2014 => to_unsigned(3250, 12), 2015 => to_unsigned(3096, 12), 2016 => to_unsigned(2048, 12), 2017 => to_unsigned(2041, 12), 2018 => to_unsigned(1111, 12), 2019 => to_unsigned(2984, 12), 2020 => to_unsigned(761, 12), 2021 => to_unsigned(3124, 12), 2022 => to_unsigned(1178, 12), 2023 => to_unsigned(731, 12), 2024 => to_unsigned(682, 12), 2025 => to_unsigned(3432, 12), 2026 => to_unsigned(2915, 12), 2027 => to_unsigned(2852, 12), 2028 => to_unsigned(455, 12), 2029 => to_unsigned(3519, 12), 2030 => to_unsigned(3275, 12), 2031 => to_unsigned(1595, 12), 2032 => to_unsigned(4068, 12), 2033 => to_unsigned(29, 12), 2034 => to_unsigned(442, 12), 2035 => to_unsigned(3413, 12), 2036 => to_unsigned(1936, 12), 2037 => to_unsigned(107, 12), 2038 => to_unsigned(70, 12), 2039 => to_unsigned(3732, 12), 2040 => to_unsigned(2802, 12), 2041 => to_unsigned(1944, 12), 2042 => to_unsigned(291, 12), 2043 => to_unsigned(1521, 12), 2044 => to_unsigned(1104, 12), 2045 => to_unsigned(1450, 12), 2046 => to_unsigned(2712, 12), 2047 => to_unsigned(1839, 12)),
            6 => (0 => to_unsigned(3099, 12), 1 => to_unsigned(2053, 12), 2 => to_unsigned(2527, 12), 3 => to_unsigned(1433, 12), 4 => to_unsigned(1223, 12), 5 => to_unsigned(2016, 12), 6 => to_unsigned(2687, 12), 7 => to_unsigned(1260, 12), 8 => to_unsigned(537, 12), 9 => to_unsigned(406, 12), 10 => to_unsigned(3983, 12), 11 => to_unsigned(1764, 12), 12 => to_unsigned(943, 12), 13 => to_unsigned(3087, 12), 14 => to_unsigned(2549, 12), 15 => to_unsigned(431, 12), 16 => to_unsigned(2986, 12), 17 => to_unsigned(1970, 12), 18 => to_unsigned(3947, 12), 19 => to_unsigned(2008, 12), 20 => to_unsigned(3566, 12), 21 => to_unsigned(653, 12), 22 => to_unsigned(2583, 12), 23 => to_unsigned(2025, 12), 24 => to_unsigned(4025, 12), 25 => to_unsigned(3121, 12), 26 => to_unsigned(3052, 12), 27 => to_unsigned(1076, 12), 28 => to_unsigned(1642, 12), 29 => to_unsigned(1746, 12), 30 => to_unsigned(2449, 12), 31 => to_unsigned(1514, 12), 32 => to_unsigned(136, 12), 33 => to_unsigned(2581, 12), 34 => to_unsigned(740, 12), 35 => to_unsigned(1293, 12), 36 => to_unsigned(4080, 12), 37 => to_unsigned(1639, 12), 38 => to_unsigned(3811, 12), 39 => to_unsigned(2128, 12), 40 => to_unsigned(2597, 12), 41 => to_unsigned(3768, 12), 42 => to_unsigned(1485, 12), 43 => to_unsigned(2209, 12), 44 => to_unsigned(1867, 12), 45 => to_unsigned(1856, 12), 46 => to_unsigned(910, 12), 47 => to_unsigned(3115, 12), 48 => to_unsigned(920, 12), 49 => to_unsigned(1115, 12), 50 => to_unsigned(1812, 12), 51 => to_unsigned(3870, 12), 52 => to_unsigned(782, 12), 53 => to_unsigned(684, 12), 54 => to_unsigned(2142, 12), 55 => to_unsigned(4095, 12), 56 => to_unsigned(144, 12), 57 => to_unsigned(639, 12), 58 => to_unsigned(1662, 12), 59 => to_unsigned(2432, 12), 60 => to_unsigned(1659, 12), 61 => to_unsigned(3827, 12), 62 => to_unsigned(688, 12), 63 => to_unsigned(2475, 12), 64 => to_unsigned(3967, 12), 65 => to_unsigned(2180, 12), 66 => to_unsigned(2244, 12), 67 => to_unsigned(658, 12), 68 => to_unsigned(1571, 12), 69 => to_unsigned(2962, 12), 70 => to_unsigned(3457, 12), 71 => to_unsigned(1979, 12), 72 => to_unsigned(2337, 12), 73 => to_unsigned(1452, 12), 74 => to_unsigned(852, 12), 75 => to_unsigned(2011, 12), 76 => to_unsigned(1780, 12), 77 => to_unsigned(169, 12), 78 => to_unsigned(1867, 12), 79 => to_unsigned(416, 12), 80 => to_unsigned(2855, 12), 81 => to_unsigned(2055, 12), 82 => to_unsigned(2803, 12), 83 => to_unsigned(1077, 12), 84 => to_unsigned(1833, 12), 85 => to_unsigned(281, 12), 86 => to_unsigned(2238, 12), 87 => to_unsigned(981, 12), 88 => to_unsigned(822, 12), 89 => to_unsigned(297, 12), 90 => to_unsigned(2336, 12), 91 => to_unsigned(878, 12), 92 => to_unsigned(521, 12), 93 => to_unsigned(639, 12), 94 => to_unsigned(1261, 12), 95 => to_unsigned(3497, 12), 96 => to_unsigned(4074, 12), 97 => to_unsigned(1607, 12), 98 => to_unsigned(1337, 12), 99 => to_unsigned(305, 12), 100 => to_unsigned(108, 12), 101 => to_unsigned(1743, 12), 102 => to_unsigned(800, 12), 103 => to_unsigned(1847, 12), 104 => to_unsigned(2136, 12), 105 => to_unsigned(3854, 12), 106 => to_unsigned(2004, 12), 107 => to_unsigned(2840, 12), 108 => to_unsigned(598, 12), 109 => to_unsigned(2786, 12), 110 => to_unsigned(2614, 12), 111 => to_unsigned(607, 12), 112 => to_unsigned(1794, 12), 113 => to_unsigned(2546, 12), 114 => to_unsigned(1586, 12), 115 => to_unsigned(1592, 12), 116 => to_unsigned(1675, 12), 117 => to_unsigned(2611, 12), 118 => to_unsigned(663, 12), 119 => to_unsigned(2859, 12), 120 => to_unsigned(1851, 12), 121 => to_unsigned(1208, 12), 122 => to_unsigned(387, 12), 123 => to_unsigned(967, 12), 124 => to_unsigned(521, 12), 125 => to_unsigned(2186, 12), 126 => to_unsigned(4062, 12), 127 => to_unsigned(3329, 12), 128 => to_unsigned(1428, 12), 129 => to_unsigned(1234, 12), 130 => to_unsigned(638, 12), 131 => to_unsigned(1325, 12), 132 => to_unsigned(293, 12), 133 => to_unsigned(23, 12), 134 => to_unsigned(3518, 12), 135 => to_unsigned(248, 12), 136 => to_unsigned(940, 12), 137 => to_unsigned(3688, 12), 138 => to_unsigned(441, 12), 139 => to_unsigned(2394, 12), 140 => to_unsigned(1580, 12), 141 => to_unsigned(381, 12), 142 => to_unsigned(3909, 12), 143 => to_unsigned(2477, 12), 144 => to_unsigned(2708, 12), 145 => to_unsigned(3121, 12), 146 => to_unsigned(2374, 12), 147 => to_unsigned(3379, 12), 148 => to_unsigned(1221, 12), 149 => to_unsigned(2189, 12), 150 => to_unsigned(3459, 12), 151 => to_unsigned(2144, 12), 152 => to_unsigned(2101, 12), 153 => to_unsigned(284, 12), 154 => to_unsigned(817, 12), 155 => to_unsigned(511, 12), 156 => to_unsigned(2200, 12), 157 => to_unsigned(1847, 12), 158 => to_unsigned(1468, 12), 159 => to_unsigned(2366, 12), 160 => to_unsigned(315, 12), 161 => to_unsigned(2605, 12), 162 => to_unsigned(3867, 12), 163 => to_unsigned(3557, 12), 164 => to_unsigned(1850, 12), 165 => to_unsigned(1666, 12), 166 => to_unsigned(557, 12), 167 => to_unsigned(3297, 12), 168 => to_unsigned(3433, 12), 169 => to_unsigned(2940, 12), 170 => to_unsigned(531, 12), 171 => to_unsigned(4048, 12), 172 => to_unsigned(3789, 12), 173 => to_unsigned(4048, 12), 174 => to_unsigned(3105, 12), 175 => to_unsigned(3127, 12), 176 => to_unsigned(2611, 12), 177 => to_unsigned(2349, 12), 178 => to_unsigned(1654, 12), 179 => to_unsigned(2807, 12), 180 => to_unsigned(3206, 12), 181 => to_unsigned(2908, 12), 182 => to_unsigned(2624, 12), 183 => to_unsigned(1950, 12), 184 => to_unsigned(2741, 12), 185 => to_unsigned(3757, 12), 186 => to_unsigned(1259, 12), 187 => to_unsigned(2248, 12), 188 => to_unsigned(3780, 12), 189 => to_unsigned(634, 12), 190 => to_unsigned(201, 12), 191 => to_unsigned(1939, 12), 192 => to_unsigned(3271, 12), 193 => to_unsigned(3621, 12), 194 => to_unsigned(1749, 12), 195 => to_unsigned(1333, 12), 196 => to_unsigned(999, 12), 197 => to_unsigned(1426, 12), 198 => to_unsigned(2083, 12), 199 => to_unsigned(858, 12), 200 => to_unsigned(2217, 12), 201 => to_unsigned(2112, 12), 202 => to_unsigned(1666, 12), 203 => to_unsigned(2911, 12), 204 => to_unsigned(2916, 12), 205 => to_unsigned(3233, 12), 206 => to_unsigned(3526, 12), 207 => to_unsigned(2409, 12), 208 => to_unsigned(589, 12), 209 => to_unsigned(3745, 12), 210 => to_unsigned(2367, 12), 211 => to_unsigned(2328, 12), 212 => to_unsigned(3814, 12), 213 => to_unsigned(2274, 12), 214 => to_unsigned(1236, 12), 215 => to_unsigned(3216, 12), 216 => to_unsigned(398, 12), 217 => to_unsigned(3982, 12), 218 => to_unsigned(1748, 12), 219 => to_unsigned(524, 12), 220 => to_unsigned(1684, 12), 221 => to_unsigned(272, 12), 222 => to_unsigned(500, 12), 223 => to_unsigned(2157, 12), 224 => to_unsigned(348, 12), 225 => to_unsigned(766, 12), 226 => to_unsigned(398, 12), 227 => to_unsigned(1701, 12), 228 => to_unsigned(3989, 12), 229 => to_unsigned(3849, 12), 230 => to_unsigned(3132, 12), 231 => to_unsigned(3180, 12), 232 => to_unsigned(484, 12), 233 => to_unsigned(3094, 12), 234 => to_unsigned(2774, 12), 235 => to_unsigned(3206, 12), 236 => to_unsigned(2543, 12), 237 => to_unsigned(1881, 12), 238 => to_unsigned(2630, 12), 239 => to_unsigned(3216, 12), 240 => to_unsigned(969, 12), 241 => to_unsigned(2360, 12), 242 => to_unsigned(3701, 12), 243 => to_unsigned(1636, 12), 244 => to_unsigned(1605, 12), 245 => to_unsigned(2340, 12), 246 => to_unsigned(1569, 12), 247 => to_unsigned(4079, 12), 248 => to_unsigned(1045, 12), 249 => to_unsigned(495, 12), 250 => to_unsigned(2874, 12), 251 => to_unsigned(253, 12), 252 => to_unsigned(1498, 12), 253 => to_unsigned(1594, 12), 254 => to_unsigned(3907, 12), 255 => to_unsigned(2249, 12), 256 => to_unsigned(831, 12), 257 => to_unsigned(3784, 12), 258 => to_unsigned(1348, 12), 259 => to_unsigned(3205, 12), 260 => to_unsigned(3919, 12), 261 => to_unsigned(1447, 12), 262 => to_unsigned(2691, 12), 263 => to_unsigned(2348, 12), 264 => to_unsigned(1680, 12), 265 => to_unsigned(2035, 12), 266 => to_unsigned(123, 12), 267 => to_unsigned(2722, 12), 268 => to_unsigned(1567, 12), 269 => to_unsigned(1270, 12), 270 => to_unsigned(1353, 12), 271 => to_unsigned(2479, 12), 272 => to_unsigned(2468, 12), 273 => to_unsigned(3486, 12), 274 => to_unsigned(1673, 12), 275 => to_unsigned(1446, 12), 276 => to_unsigned(3744, 12), 277 => to_unsigned(514, 12), 278 => to_unsigned(953, 12), 279 => to_unsigned(3595, 12), 280 => to_unsigned(3822, 12), 281 => to_unsigned(822, 12), 282 => to_unsigned(2291, 12), 283 => to_unsigned(344, 12), 284 => to_unsigned(3288, 12), 285 => to_unsigned(1979, 12), 286 => to_unsigned(183, 12), 287 => to_unsigned(2985, 12), 288 => to_unsigned(2801, 12), 289 => to_unsigned(3739, 12), 290 => to_unsigned(1101, 12), 291 => to_unsigned(2219, 12), 292 => to_unsigned(3455, 12), 293 => to_unsigned(107, 12), 294 => to_unsigned(3247, 12), 295 => to_unsigned(3524, 12), 296 => to_unsigned(274, 12), 297 => to_unsigned(3525, 12), 298 => to_unsigned(2310, 12), 299 => to_unsigned(3148, 12), 300 => to_unsigned(3428, 12), 301 => to_unsigned(2091, 12), 302 => to_unsigned(714, 12), 303 => to_unsigned(3631, 12), 304 => to_unsigned(1771, 12), 305 => to_unsigned(3067, 12), 306 => to_unsigned(4024, 12), 307 => to_unsigned(2274, 12), 308 => to_unsigned(1313, 12), 309 => to_unsigned(3283, 12), 310 => to_unsigned(1426, 12), 311 => to_unsigned(141, 12), 312 => to_unsigned(488, 12), 313 => to_unsigned(3125, 12), 314 => to_unsigned(401, 12), 315 => to_unsigned(2494, 12), 316 => to_unsigned(181, 12), 317 => to_unsigned(4089, 12), 318 => to_unsigned(1510, 12), 319 => to_unsigned(129, 12), 320 => to_unsigned(3274, 12), 321 => to_unsigned(3723, 12), 322 => to_unsigned(2935, 12), 323 => to_unsigned(784, 12), 324 => to_unsigned(2735, 12), 325 => to_unsigned(1813, 12), 326 => to_unsigned(403, 12), 327 => to_unsigned(1854, 12), 328 => to_unsigned(1631, 12), 329 => to_unsigned(818, 12), 330 => to_unsigned(1898, 12), 331 => to_unsigned(1609, 12), 332 => to_unsigned(1701, 12), 333 => to_unsigned(429, 12), 334 => to_unsigned(854, 12), 335 => to_unsigned(1875, 12), 336 => to_unsigned(2688, 12), 337 => to_unsigned(2310, 12), 338 => to_unsigned(3330, 12), 339 => to_unsigned(3699, 12), 340 => to_unsigned(3498, 12), 341 => to_unsigned(3191, 12), 342 => to_unsigned(2096, 12), 343 => to_unsigned(1345, 12), 344 => to_unsigned(3913, 12), 345 => to_unsigned(2225, 12), 346 => to_unsigned(1623, 12), 347 => to_unsigned(2647, 12), 348 => to_unsigned(3173, 12), 349 => to_unsigned(2587, 12), 350 => to_unsigned(1116, 12), 351 => to_unsigned(2238, 12), 352 => to_unsigned(2299, 12), 353 => to_unsigned(3429, 12), 354 => to_unsigned(4005, 12), 355 => to_unsigned(4071, 12), 356 => to_unsigned(2857, 12), 357 => to_unsigned(2799, 12), 358 => to_unsigned(706, 12), 359 => to_unsigned(1879, 12), 360 => to_unsigned(947, 12), 361 => to_unsigned(2018, 12), 362 => to_unsigned(576, 12), 363 => to_unsigned(2916, 12), 364 => to_unsigned(1987, 12), 365 => to_unsigned(2028, 12), 366 => to_unsigned(2240, 12), 367 => to_unsigned(3063, 12), 368 => to_unsigned(2585, 12), 369 => to_unsigned(1051, 12), 370 => to_unsigned(3172, 12), 371 => to_unsigned(1200, 12), 372 => to_unsigned(321, 12), 373 => to_unsigned(760, 12), 374 => to_unsigned(1543, 12), 375 => to_unsigned(2913, 12), 376 => to_unsigned(2716, 12), 377 => to_unsigned(3748, 12), 378 => to_unsigned(3821, 12), 379 => to_unsigned(1446, 12), 380 => to_unsigned(2664, 12), 381 => to_unsigned(573, 12), 382 => to_unsigned(2085, 12), 383 => to_unsigned(2147, 12), 384 => to_unsigned(465, 12), 385 => to_unsigned(3259, 12), 386 => to_unsigned(90, 12), 387 => to_unsigned(3637, 12), 388 => to_unsigned(2610, 12), 389 => to_unsigned(2367, 12), 390 => to_unsigned(4095, 12), 391 => to_unsigned(2317, 12), 392 => to_unsigned(542, 12), 393 => to_unsigned(83, 12), 394 => to_unsigned(3348, 12), 395 => to_unsigned(1326, 12), 396 => to_unsigned(1036, 12), 397 => to_unsigned(1969, 12), 398 => to_unsigned(1324, 12), 399 => to_unsigned(1641, 12), 400 => to_unsigned(509, 12), 401 => to_unsigned(1011, 12), 402 => to_unsigned(2236, 12), 403 => to_unsigned(1994, 12), 404 => to_unsigned(3885, 12), 405 => to_unsigned(1270, 12), 406 => to_unsigned(2349, 12), 407 => to_unsigned(532, 12), 408 => to_unsigned(2366, 12), 409 => to_unsigned(603, 12), 410 => to_unsigned(1431, 12), 411 => to_unsigned(1186, 12), 412 => to_unsigned(1186, 12), 413 => to_unsigned(977, 12), 414 => to_unsigned(1598, 12), 415 => to_unsigned(486, 12), 416 => to_unsigned(348, 12), 417 => to_unsigned(64, 12), 418 => to_unsigned(3516, 12), 419 => to_unsigned(826, 12), 420 => to_unsigned(3065, 12), 421 => to_unsigned(3308, 12), 422 => to_unsigned(2483, 12), 423 => to_unsigned(423, 12), 424 => to_unsigned(2895, 12), 425 => to_unsigned(3427, 12), 426 => to_unsigned(1291, 12), 427 => to_unsigned(1558, 12), 428 => to_unsigned(444, 12), 429 => to_unsigned(1336, 12), 430 => to_unsigned(1293, 12), 431 => to_unsigned(3326, 12), 432 => to_unsigned(1404, 12), 433 => to_unsigned(1065, 12), 434 => to_unsigned(1509, 12), 435 => to_unsigned(2295, 12), 436 => to_unsigned(392, 12), 437 => to_unsigned(1985, 12), 438 => to_unsigned(3303, 12), 439 => to_unsigned(1510, 12), 440 => to_unsigned(2585, 12), 441 => to_unsigned(928, 12), 442 => to_unsigned(2577, 12), 443 => to_unsigned(2773, 12), 444 => to_unsigned(364, 12), 445 => to_unsigned(2754, 12), 446 => to_unsigned(12, 12), 447 => to_unsigned(484, 12), 448 => to_unsigned(3852, 12), 449 => to_unsigned(3072, 12), 450 => to_unsigned(3267, 12), 451 => to_unsigned(1124, 12), 452 => to_unsigned(3006, 12), 453 => to_unsigned(3189, 12), 454 => to_unsigned(506, 12), 455 => to_unsigned(1785, 12), 456 => to_unsigned(193, 12), 457 => to_unsigned(4008, 12), 458 => to_unsigned(1351, 12), 459 => to_unsigned(3016, 12), 460 => to_unsigned(3036, 12), 461 => to_unsigned(3364, 12), 462 => to_unsigned(1023, 12), 463 => to_unsigned(1505, 12), 464 => to_unsigned(3717, 12), 465 => to_unsigned(1629, 12), 466 => to_unsigned(4038, 12), 467 => to_unsigned(1693, 12), 468 => to_unsigned(3029, 12), 469 => to_unsigned(637, 12), 470 => to_unsigned(2536, 12), 471 => to_unsigned(142, 12), 472 => to_unsigned(182, 12), 473 => to_unsigned(34, 12), 474 => to_unsigned(4012, 12), 475 => to_unsigned(2735, 12), 476 => to_unsigned(1696, 12), 477 => to_unsigned(2779, 12), 478 => to_unsigned(140, 12), 479 => to_unsigned(2271, 12), 480 => to_unsigned(575, 12), 481 => to_unsigned(3535, 12), 482 => to_unsigned(1099, 12), 483 => to_unsigned(1531, 12), 484 => to_unsigned(3308, 12), 485 => to_unsigned(2225, 12), 486 => to_unsigned(369, 12), 487 => to_unsigned(1440, 12), 488 => to_unsigned(1857, 12), 489 => to_unsigned(1358, 12), 490 => to_unsigned(3881, 12), 491 => to_unsigned(2529, 12), 492 => to_unsigned(219, 12), 493 => to_unsigned(2875, 12), 494 => to_unsigned(597, 12), 495 => to_unsigned(2299, 12), 496 => to_unsigned(353, 12), 497 => to_unsigned(3306, 12), 498 => to_unsigned(4010, 12), 499 => to_unsigned(4069, 12), 500 => to_unsigned(3585, 12), 501 => to_unsigned(19, 12), 502 => to_unsigned(3467, 12), 503 => to_unsigned(1668, 12), 504 => to_unsigned(777, 12), 505 => to_unsigned(795, 12), 506 => to_unsigned(2895, 12), 507 => to_unsigned(705, 12), 508 => to_unsigned(2915, 12), 509 => to_unsigned(2048, 12), 510 => to_unsigned(3408, 12), 511 => to_unsigned(1608, 12), 512 => to_unsigned(3345, 12), 513 => to_unsigned(742, 12), 514 => to_unsigned(1748, 12), 515 => to_unsigned(1787, 12), 516 => to_unsigned(50, 12), 517 => to_unsigned(3328, 12), 518 => to_unsigned(279, 12), 519 => to_unsigned(2605, 12), 520 => to_unsigned(337, 12), 521 => to_unsigned(625, 12), 522 => to_unsigned(1224, 12), 523 => to_unsigned(3081, 12), 524 => to_unsigned(1371, 12), 525 => to_unsigned(2889, 12), 526 => to_unsigned(1394, 12), 527 => to_unsigned(178, 12), 528 => to_unsigned(4006, 12), 529 => to_unsigned(3359, 12), 530 => to_unsigned(2439, 12), 531 => to_unsigned(1021, 12), 532 => to_unsigned(3530, 12), 533 => to_unsigned(3309, 12), 534 => to_unsigned(198, 12), 535 => to_unsigned(2175, 12), 536 => to_unsigned(1222, 12), 537 => to_unsigned(2939, 12), 538 => to_unsigned(1637, 12), 539 => to_unsigned(4030, 12), 540 => to_unsigned(2611, 12), 541 => to_unsigned(2514, 12), 542 => to_unsigned(2475, 12), 543 => to_unsigned(4013, 12), 544 => to_unsigned(3889, 12), 545 => to_unsigned(1375, 12), 546 => to_unsigned(3033, 12), 547 => to_unsigned(2608, 12), 548 => to_unsigned(1509, 12), 549 => to_unsigned(3790, 12), 550 => to_unsigned(805, 12), 551 => to_unsigned(2480, 12), 552 => to_unsigned(1240, 12), 553 => to_unsigned(3523, 12), 554 => to_unsigned(2942, 12), 555 => to_unsigned(490, 12), 556 => to_unsigned(1579, 12), 557 => to_unsigned(1722, 12), 558 => to_unsigned(1566, 12), 559 => to_unsigned(3528, 12), 560 => to_unsigned(3664, 12), 561 => to_unsigned(2709, 12), 562 => to_unsigned(3718, 12), 563 => to_unsigned(1277, 12), 564 => to_unsigned(1604, 12), 565 => to_unsigned(1694, 12), 566 => to_unsigned(3580, 12), 567 => to_unsigned(2391, 12), 568 => to_unsigned(369, 12), 569 => to_unsigned(1718, 12), 570 => to_unsigned(377, 12), 571 => to_unsigned(1724, 12), 572 => to_unsigned(1217, 12), 573 => to_unsigned(2418, 12), 574 => to_unsigned(1832, 12), 575 => to_unsigned(2439, 12), 576 => to_unsigned(329, 12), 577 => to_unsigned(3966, 12), 578 => to_unsigned(2855, 12), 579 => to_unsigned(1010, 12), 580 => to_unsigned(2285, 12), 581 => to_unsigned(1928, 12), 582 => to_unsigned(3356, 12), 583 => to_unsigned(1552, 12), 584 => to_unsigned(1556, 12), 585 => to_unsigned(2308, 12), 586 => to_unsigned(1443, 12), 587 => to_unsigned(827, 12), 588 => to_unsigned(3578, 12), 589 => to_unsigned(3560, 12), 590 => to_unsigned(233, 12), 591 => to_unsigned(463, 12), 592 => to_unsigned(622, 12), 593 => to_unsigned(2403, 12), 594 => to_unsigned(1953, 12), 595 => to_unsigned(1356, 12), 596 => to_unsigned(3278, 12), 597 => to_unsigned(3250, 12), 598 => to_unsigned(3938, 12), 599 => to_unsigned(3779, 12), 600 => to_unsigned(2437, 12), 601 => to_unsigned(927, 12), 602 => to_unsigned(4055, 12), 603 => to_unsigned(50, 12), 604 => to_unsigned(4072, 12), 605 => to_unsigned(2124, 12), 606 => to_unsigned(2752, 12), 607 => to_unsigned(2074, 12), 608 => to_unsigned(3159, 12), 609 => to_unsigned(1038, 12), 610 => to_unsigned(2841, 12), 611 => to_unsigned(3663, 12), 612 => to_unsigned(584, 12), 613 => to_unsigned(667, 12), 614 => to_unsigned(2211, 12), 615 => to_unsigned(2941, 12), 616 => to_unsigned(279, 12), 617 => to_unsigned(2763, 12), 618 => to_unsigned(2155, 12), 619 => to_unsigned(901, 12), 620 => to_unsigned(2818, 12), 621 => to_unsigned(1204, 12), 622 => to_unsigned(3345, 12), 623 => to_unsigned(1252, 12), 624 => to_unsigned(1191, 12), 625 => to_unsigned(3015, 12), 626 => to_unsigned(2145, 12), 627 => to_unsigned(2719, 12), 628 => to_unsigned(1564, 12), 629 => to_unsigned(907, 12), 630 => to_unsigned(1659, 12), 631 => to_unsigned(3959, 12), 632 => to_unsigned(2236, 12), 633 => to_unsigned(3819, 12), 634 => to_unsigned(884, 12), 635 => to_unsigned(3901, 12), 636 => to_unsigned(2332, 12), 637 => to_unsigned(2715, 12), 638 => to_unsigned(2135, 12), 639 => to_unsigned(2016, 12), 640 => to_unsigned(2543, 12), 641 => to_unsigned(3284, 12), 642 => to_unsigned(2494, 12), 643 => to_unsigned(3580, 12), 644 => to_unsigned(611, 12), 645 => to_unsigned(1274, 12), 646 => to_unsigned(2784, 12), 647 => to_unsigned(380, 12), 648 => to_unsigned(3331, 12), 649 => to_unsigned(716, 12), 650 => to_unsigned(3191, 12), 651 => to_unsigned(3233, 12), 652 => to_unsigned(486, 12), 653 => to_unsigned(2023, 12), 654 => to_unsigned(2363, 12), 655 => to_unsigned(2110, 12), 656 => to_unsigned(540, 12), 657 => to_unsigned(115, 12), 658 => to_unsigned(849, 12), 659 => to_unsigned(1753, 12), 660 => to_unsigned(2234, 12), 661 => to_unsigned(2586, 12), 662 => to_unsigned(3547, 12), 663 => to_unsigned(1090, 12), 664 => to_unsigned(3386, 12), 665 => to_unsigned(892, 12), 666 => to_unsigned(3731, 12), 667 => to_unsigned(3424, 12), 668 => to_unsigned(729, 12), 669 => to_unsigned(3035, 12), 670 => to_unsigned(2572, 12), 671 => to_unsigned(3567, 12), 672 => to_unsigned(3965, 12), 673 => to_unsigned(1963, 12), 674 => to_unsigned(1348, 12), 675 => to_unsigned(1029, 12), 676 => to_unsigned(566, 12), 677 => to_unsigned(1586, 12), 678 => to_unsigned(1428, 12), 679 => to_unsigned(1853, 12), 680 => to_unsigned(1691, 12), 681 => to_unsigned(3459, 12), 682 => to_unsigned(2240, 12), 683 => to_unsigned(98, 12), 684 => to_unsigned(1838, 12), 685 => to_unsigned(2417, 12), 686 => to_unsigned(1481, 12), 687 => to_unsigned(4030, 12), 688 => to_unsigned(1827, 12), 689 => to_unsigned(677, 12), 690 => to_unsigned(2049, 12), 691 => to_unsigned(3501, 12), 692 => to_unsigned(1889, 12), 693 => to_unsigned(2522, 12), 694 => to_unsigned(4044, 12), 695 => to_unsigned(2584, 12), 696 => to_unsigned(1175, 12), 697 => to_unsigned(2913, 12), 698 => to_unsigned(926, 12), 699 => to_unsigned(2184, 12), 700 => to_unsigned(3772, 12), 701 => to_unsigned(3559, 12), 702 => to_unsigned(159, 12), 703 => to_unsigned(2500, 12), 704 => to_unsigned(3883, 12), 705 => to_unsigned(3022, 12), 706 => to_unsigned(4027, 12), 707 => to_unsigned(3979, 12), 708 => to_unsigned(733, 12), 709 => to_unsigned(1565, 12), 710 => to_unsigned(1937, 12), 711 => to_unsigned(3177, 12), 712 => to_unsigned(452, 12), 713 => to_unsigned(3586, 12), 714 => to_unsigned(2444, 12), 715 => to_unsigned(646, 12), 716 => to_unsigned(2957, 12), 717 => to_unsigned(371, 12), 718 => to_unsigned(3502, 12), 719 => to_unsigned(1998, 12), 720 => to_unsigned(263, 12), 721 => to_unsigned(493, 12), 722 => to_unsigned(1587, 12), 723 => to_unsigned(598, 12), 724 => to_unsigned(1128, 12), 725 => to_unsigned(1131, 12), 726 => to_unsigned(3846, 12), 727 => to_unsigned(3654, 12), 728 => to_unsigned(2114, 12), 729 => to_unsigned(2743, 12), 730 => to_unsigned(1808, 12), 731 => to_unsigned(2968, 12), 732 => to_unsigned(3842, 12), 733 => to_unsigned(1559, 12), 734 => to_unsigned(1631, 12), 735 => to_unsigned(4010, 12), 736 => to_unsigned(1418, 12), 737 => to_unsigned(245, 12), 738 => to_unsigned(1797, 12), 739 => to_unsigned(1118, 12), 740 => to_unsigned(3081, 12), 741 => to_unsigned(767, 12), 742 => to_unsigned(818, 12), 743 => to_unsigned(1142, 12), 744 => to_unsigned(1261, 12), 745 => to_unsigned(2890, 12), 746 => to_unsigned(940, 12), 747 => to_unsigned(2992, 12), 748 => to_unsigned(4058, 12), 749 => to_unsigned(2753, 12), 750 => to_unsigned(1276, 12), 751 => to_unsigned(3490, 12), 752 => to_unsigned(3964, 12), 753 => to_unsigned(2984, 12), 754 => to_unsigned(3266, 12), 755 => to_unsigned(3379, 12), 756 => to_unsigned(1728, 12), 757 => to_unsigned(4051, 12), 758 => to_unsigned(1451, 12), 759 => to_unsigned(3176, 12), 760 => to_unsigned(3841, 12), 761 => to_unsigned(2030, 12), 762 => to_unsigned(3145, 12), 763 => to_unsigned(659, 12), 764 => to_unsigned(2156, 12), 765 => to_unsigned(3270, 12), 766 => to_unsigned(884, 12), 767 => to_unsigned(3786, 12), 768 => to_unsigned(481, 12), 769 => to_unsigned(2646, 12), 770 => to_unsigned(3744, 12), 771 => to_unsigned(1356, 12), 772 => to_unsigned(3970, 12), 773 => to_unsigned(1607, 12), 774 => to_unsigned(1351, 12), 775 => to_unsigned(1352, 12), 776 => to_unsigned(1011, 12), 777 => to_unsigned(2819, 12), 778 => to_unsigned(3761, 12), 779 => to_unsigned(512, 12), 780 => to_unsigned(850, 12), 781 => to_unsigned(2256, 12), 782 => to_unsigned(1810, 12), 783 => to_unsigned(2304, 12), 784 => to_unsigned(3355, 12), 785 => to_unsigned(2260, 12), 786 => to_unsigned(2042, 12), 787 => to_unsigned(1994, 12), 788 => to_unsigned(1901, 12), 789 => to_unsigned(52, 12), 790 => to_unsigned(1987, 12), 791 => to_unsigned(1509, 12), 792 => to_unsigned(531, 12), 793 => to_unsigned(2387, 12), 794 => to_unsigned(338, 12), 795 => to_unsigned(2544, 12), 796 => to_unsigned(837, 12), 797 => to_unsigned(2546, 12), 798 => to_unsigned(3714, 12), 799 => to_unsigned(2581, 12), 800 => to_unsigned(103, 12), 801 => to_unsigned(802, 12), 802 => to_unsigned(810, 12), 803 => to_unsigned(3609, 12), 804 => to_unsigned(3938, 12), 805 => to_unsigned(2267, 12), 806 => to_unsigned(1512, 12), 807 => to_unsigned(3326, 12), 808 => to_unsigned(3647, 12), 809 => to_unsigned(2598, 12), 810 => to_unsigned(2713, 12), 811 => to_unsigned(2923, 12), 812 => to_unsigned(205, 12), 813 => to_unsigned(2350, 12), 814 => to_unsigned(1119, 12), 815 => to_unsigned(3633, 12), 816 => to_unsigned(843, 12), 817 => to_unsigned(3827, 12), 818 => to_unsigned(2381, 12), 819 => to_unsigned(1342, 12), 820 => to_unsigned(551, 12), 821 => to_unsigned(3714, 12), 822 => to_unsigned(2691, 12), 823 => to_unsigned(1052, 12), 824 => to_unsigned(1497, 12), 825 => to_unsigned(774, 12), 826 => to_unsigned(2501, 12), 827 => to_unsigned(3341, 12), 828 => to_unsigned(562, 12), 829 => to_unsigned(864, 12), 830 => to_unsigned(1587, 12), 831 => to_unsigned(1451, 12), 832 => to_unsigned(2773, 12), 833 => to_unsigned(1874, 12), 834 => to_unsigned(3164, 12), 835 => to_unsigned(2089, 12), 836 => to_unsigned(2454, 12), 837 => to_unsigned(3963, 12), 838 => to_unsigned(205, 12), 839 => to_unsigned(2092, 12), 840 => to_unsigned(549, 12), 841 => to_unsigned(534, 12), 842 => to_unsigned(2624, 12), 843 => to_unsigned(1570, 12), 844 => to_unsigned(2629, 12), 845 => to_unsigned(1535, 12), 846 => to_unsigned(1128, 12), 847 => to_unsigned(495, 12), 848 => to_unsigned(3100, 12), 849 => to_unsigned(3603, 12), 850 => to_unsigned(661, 12), 851 => to_unsigned(2672, 12), 852 => to_unsigned(811, 12), 853 => to_unsigned(3589, 12), 854 => to_unsigned(958, 12), 855 => to_unsigned(1040, 12), 856 => to_unsigned(2843, 12), 857 => to_unsigned(808, 12), 858 => to_unsigned(3027, 12), 859 => to_unsigned(1498, 12), 860 => to_unsigned(203, 12), 861 => to_unsigned(2840, 12), 862 => to_unsigned(1197, 12), 863 => to_unsigned(383, 12), 864 => to_unsigned(3948, 12), 865 => to_unsigned(3246, 12), 866 => to_unsigned(2095, 12), 867 => to_unsigned(1775, 12), 868 => to_unsigned(633, 12), 869 => to_unsigned(3700, 12), 870 => to_unsigned(1894, 12), 871 => to_unsigned(2313, 12), 872 => to_unsigned(3435, 12), 873 => to_unsigned(2661, 12), 874 => to_unsigned(80, 12), 875 => to_unsigned(776, 12), 876 => to_unsigned(1432, 12), 877 => to_unsigned(1640, 12), 878 => to_unsigned(250, 12), 879 => to_unsigned(1083, 12), 880 => to_unsigned(3457, 12), 881 => to_unsigned(1740, 12), 882 => to_unsigned(3225, 12), 883 => to_unsigned(2371, 12), 884 => to_unsigned(3613, 12), 885 => to_unsigned(3758, 12), 886 => to_unsigned(2252, 12), 887 => to_unsigned(3785, 12), 888 => to_unsigned(2355, 12), 889 => to_unsigned(2514, 12), 890 => to_unsigned(3995, 12), 891 => to_unsigned(1841, 12), 892 => to_unsigned(569, 12), 893 => to_unsigned(4024, 12), 894 => to_unsigned(2776, 12), 895 => to_unsigned(3677, 12), 896 => to_unsigned(3382, 12), 897 => to_unsigned(2357, 12), 898 => to_unsigned(399, 12), 899 => to_unsigned(3678, 12), 900 => to_unsigned(2782, 12), 901 => to_unsigned(2578, 12), 902 => to_unsigned(1460, 12), 903 => to_unsigned(3789, 12), 904 => to_unsigned(3691, 12), 905 => to_unsigned(1038, 12), 906 => to_unsigned(1160, 12), 907 => to_unsigned(1490, 12), 908 => to_unsigned(1540, 12), 909 => to_unsigned(1357, 12), 910 => to_unsigned(502, 12), 911 => to_unsigned(2778, 12), 912 => to_unsigned(569, 12), 913 => to_unsigned(1118, 12), 914 => to_unsigned(3984, 12), 915 => to_unsigned(1806, 12), 916 => to_unsigned(1401, 12), 917 => to_unsigned(938, 12), 918 => to_unsigned(3297, 12), 919 => to_unsigned(424, 12), 920 => to_unsigned(3350, 12), 921 => to_unsigned(97, 12), 922 => to_unsigned(2362, 12), 923 => to_unsigned(3838, 12), 924 => to_unsigned(1133, 12), 925 => to_unsigned(1831, 12), 926 => to_unsigned(3100, 12), 927 => to_unsigned(3935, 12), 928 => to_unsigned(3821, 12), 929 => to_unsigned(53, 12), 930 => to_unsigned(2556, 12), 931 => to_unsigned(3465, 12), 932 => to_unsigned(1891, 12), 933 => to_unsigned(3556, 12), 934 => to_unsigned(2230, 12), 935 => to_unsigned(3904, 12), 936 => to_unsigned(169, 12), 937 => to_unsigned(2968, 12), 938 => to_unsigned(3683, 12), 939 => to_unsigned(2856, 12), 940 => to_unsigned(1286, 12), 941 => to_unsigned(1681, 12), 942 => to_unsigned(225, 12), 943 => to_unsigned(3948, 12), 944 => to_unsigned(2424, 12), 945 => to_unsigned(1085, 12), 946 => to_unsigned(3531, 12), 947 => to_unsigned(1595, 12), 948 => to_unsigned(2279, 12), 949 => to_unsigned(1592, 12), 950 => to_unsigned(3780, 12), 951 => to_unsigned(2873, 12), 952 => to_unsigned(117, 12), 953 => to_unsigned(1397, 12), 954 => to_unsigned(2217, 12), 955 => to_unsigned(3548, 12), 956 => to_unsigned(3897, 12), 957 => to_unsigned(864, 12), 958 => to_unsigned(3857, 12), 959 => to_unsigned(9, 12), 960 => to_unsigned(3633, 12), 961 => to_unsigned(2460, 12), 962 => to_unsigned(2984, 12), 963 => to_unsigned(3795, 12), 964 => to_unsigned(1645, 12), 965 => to_unsigned(329, 12), 966 => to_unsigned(651, 12), 967 => to_unsigned(282, 12), 968 => to_unsigned(2540, 12), 969 => to_unsigned(150, 12), 970 => to_unsigned(2031, 12), 971 => to_unsigned(1224, 12), 972 => to_unsigned(104, 12), 973 => to_unsigned(53, 12), 974 => to_unsigned(3778, 12), 975 => to_unsigned(2191, 12), 976 => to_unsigned(410, 12), 977 => to_unsigned(3246, 12), 978 => to_unsigned(1565, 12), 979 => to_unsigned(2955, 12), 980 => to_unsigned(3514, 12), 981 => to_unsigned(187, 12), 982 => to_unsigned(273, 12), 983 => to_unsigned(2801, 12), 984 => to_unsigned(1326, 12), 985 => to_unsigned(4064, 12), 986 => to_unsigned(1191, 12), 987 => to_unsigned(1212, 12), 988 => to_unsigned(135, 12), 989 => to_unsigned(709, 12), 990 => to_unsigned(1274, 12), 991 => to_unsigned(529, 12), 992 => to_unsigned(264, 12), 993 => to_unsigned(1438, 12), 994 => to_unsigned(4012, 12), 995 => to_unsigned(1264, 12), 996 => to_unsigned(893, 12), 997 => to_unsigned(3722, 12), 998 => to_unsigned(1378, 12), 999 => to_unsigned(2796, 12), 1000 => to_unsigned(1938, 12), 1001 => to_unsigned(3567, 12), 1002 => to_unsigned(2109, 12), 1003 => to_unsigned(3205, 12), 1004 => to_unsigned(29, 12), 1005 => to_unsigned(3639, 12), 1006 => to_unsigned(2689, 12), 1007 => to_unsigned(3175, 12), 1008 => to_unsigned(932, 12), 1009 => to_unsigned(1182, 12), 1010 => to_unsigned(2126, 12), 1011 => to_unsigned(2824, 12), 1012 => to_unsigned(3304, 12), 1013 => to_unsigned(3165, 12), 1014 => to_unsigned(1154, 12), 1015 => to_unsigned(1787, 12), 1016 => to_unsigned(3224, 12), 1017 => to_unsigned(3559, 12), 1018 => to_unsigned(298, 12), 1019 => to_unsigned(1474, 12), 1020 => to_unsigned(1218, 12), 1021 => to_unsigned(727, 12), 1022 => to_unsigned(614, 12), 1023 => to_unsigned(3912, 12), 1024 => to_unsigned(124, 12), 1025 => to_unsigned(1634, 12), 1026 => to_unsigned(1353, 12), 1027 => to_unsigned(542, 12), 1028 => to_unsigned(514, 12), 1029 => to_unsigned(432, 12), 1030 => to_unsigned(2961, 12), 1031 => to_unsigned(1436, 12), 1032 => to_unsigned(403, 12), 1033 => to_unsigned(2545, 12), 1034 => to_unsigned(2573, 12), 1035 => to_unsigned(880, 12), 1036 => to_unsigned(1092, 12), 1037 => to_unsigned(172, 12), 1038 => to_unsigned(650, 12), 1039 => to_unsigned(3907, 12), 1040 => to_unsigned(4045, 12), 1041 => to_unsigned(712, 12), 1042 => to_unsigned(1033, 12), 1043 => to_unsigned(1269, 12), 1044 => to_unsigned(2186, 12), 1045 => to_unsigned(1986, 12), 1046 => to_unsigned(2423, 12), 1047 => to_unsigned(3762, 12), 1048 => to_unsigned(564, 12), 1049 => to_unsigned(966, 12), 1050 => to_unsigned(2996, 12), 1051 => to_unsigned(1701, 12), 1052 => to_unsigned(1600, 12), 1053 => to_unsigned(1561, 12), 1054 => to_unsigned(925, 12), 1055 => to_unsigned(648, 12), 1056 => to_unsigned(230, 12), 1057 => to_unsigned(774, 12), 1058 => to_unsigned(2382, 12), 1059 => to_unsigned(1786, 12), 1060 => to_unsigned(305, 12), 1061 => to_unsigned(717, 12), 1062 => to_unsigned(937, 12), 1063 => to_unsigned(994, 12), 1064 => to_unsigned(3280, 12), 1065 => to_unsigned(3054, 12), 1066 => to_unsigned(1373, 12), 1067 => to_unsigned(2241, 12), 1068 => to_unsigned(3128, 12), 1069 => to_unsigned(3846, 12), 1070 => to_unsigned(1650, 12), 1071 => to_unsigned(760, 12), 1072 => to_unsigned(1837, 12), 1073 => to_unsigned(679, 12), 1074 => to_unsigned(390, 12), 1075 => to_unsigned(3801, 12), 1076 => to_unsigned(716, 12), 1077 => to_unsigned(1468, 12), 1078 => to_unsigned(3709, 12), 1079 => to_unsigned(193, 12), 1080 => to_unsigned(3877, 12), 1081 => to_unsigned(2878, 12), 1082 => to_unsigned(1976, 12), 1083 => to_unsigned(2909, 12), 1084 => to_unsigned(474, 12), 1085 => to_unsigned(2235, 12), 1086 => to_unsigned(3166, 12), 1087 => to_unsigned(205, 12), 1088 => to_unsigned(2287, 12), 1089 => to_unsigned(527, 12), 1090 => to_unsigned(2610, 12), 1091 => to_unsigned(3901, 12), 1092 => to_unsigned(1176, 12), 1093 => to_unsigned(3360, 12), 1094 => to_unsigned(3964, 12), 1095 => to_unsigned(3757, 12), 1096 => to_unsigned(370, 12), 1097 => to_unsigned(2886, 12), 1098 => to_unsigned(3222, 12), 1099 => to_unsigned(2322, 12), 1100 => to_unsigned(494, 12), 1101 => to_unsigned(2384, 12), 1102 => to_unsigned(2875, 12), 1103 => to_unsigned(1340, 12), 1104 => to_unsigned(3512, 12), 1105 => to_unsigned(10, 12), 1106 => to_unsigned(1872, 12), 1107 => to_unsigned(1068, 12), 1108 => to_unsigned(2991, 12), 1109 => to_unsigned(2751, 12), 1110 => to_unsigned(2147, 12), 1111 => to_unsigned(890, 12), 1112 => to_unsigned(3286, 12), 1113 => to_unsigned(2889, 12), 1114 => to_unsigned(841, 12), 1115 => to_unsigned(3519, 12), 1116 => to_unsigned(3839, 12), 1117 => to_unsigned(1847, 12), 1118 => to_unsigned(2408, 12), 1119 => to_unsigned(2046, 12), 1120 => to_unsigned(3891, 12), 1121 => to_unsigned(2069, 12), 1122 => to_unsigned(889, 12), 1123 => to_unsigned(110, 12), 1124 => to_unsigned(3998, 12), 1125 => to_unsigned(1634, 12), 1126 => to_unsigned(728, 12), 1127 => to_unsigned(1477, 12), 1128 => to_unsigned(2598, 12), 1129 => to_unsigned(2269, 12), 1130 => to_unsigned(2347, 12), 1131 => to_unsigned(1886, 12), 1132 => to_unsigned(1353, 12), 1133 => to_unsigned(3015, 12), 1134 => to_unsigned(2187, 12), 1135 => to_unsigned(3098, 12), 1136 => to_unsigned(612, 12), 1137 => to_unsigned(3436, 12), 1138 => to_unsigned(2167, 12), 1139 => to_unsigned(2342, 12), 1140 => to_unsigned(758, 12), 1141 => to_unsigned(2896, 12), 1142 => to_unsigned(769, 12), 1143 => to_unsigned(1010, 12), 1144 => to_unsigned(1317, 12), 1145 => to_unsigned(579, 12), 1146 => to_unsigned(3121, 12), 1147 => to_unsigned(3690, 12), 1148 => to_unsigned(2391, 12), 1149 => to_unsigned(2979, 12), 1150 => to_unsigned(1845, 12), 1151 => to_unsigned(1641, 12), 1152 => to_unsigned(537, 12), 1153 => to_unsigned(1804, 12), 1154 => to_unsigned(3186, 12), 1155 => to_unsigned(2397, 12), 1156 => to_unsigned(1874, 12), 1157 => to_unsigned(3015, 12), 1158 => to_unsigned(3276, 12), 1159 => to_unsigned(2784, 12), 1160 => to_unsigned(2120, 12), 1161 => to_unsigned(3291, 12), 1162 => to_unsigned(688, 12), 1163 => to_unsigned(3578, 12), 1164 => to_unsigned(1565, 12), 1165 => to_unsigned(3600, 12), 1166 => to_unsigned(87, 12), 1167 => to_unsigned(2546, 12), 1168 => to_unsigned(1502, 12), 1169 => to_unsigned(2679, 12), 1170 => to_unsigned(1997, 12), 1171 => to_unsigned(49, 12), 1172 => to_unsigned(1736, 12), 1173 => to_unsigned(3941, 12), 1174 => to_unsigned(2320, 12), 1175 => to_unsigned(1394, 12), 1176 => to_unsigned(552, 12), 1177 => to_unsigned(4062, 12), 1178 => to_unsigned(1633, 12), 1179 => to_unsigned(419, 12), 1180 => to_unsigned(894, 12), 1181 => to_unsigned(1515, 12), 1182 => to_unsigned(3536, 12), 1183 => to_unsigned(2667, 12), 1184 => to_unsigned(43, 12), 1185 => to_unsigned(1115, 12), 1186 => to_unsigned(1698, 12), 1187 => to_unsigned(140, 12), 1188 => to_unsigned(3145, 12), 1189 => to_unsigned(1381, 12), 1190 => to_unsigned(1148, 12), 1191 => to_unsigned(2507, 12), 1192 => to_unsigned(2656, 12), 1193 => to_unsigned(1410, 12), 1194 => to_unsigned(2141, 12), 1195 => to_unsigned(1958, 12), 1196 => to_unsigned(3324, 12), 1197 => to_unsigned(3482, 12), 1198 => to_unsigned(2128, 12), 1199 => to_unsigned(1479, 12), 1200 => to_unsigned(489, 12), 1201 => to_unsigned(3674, 12), 1202 => to_unsigned(2633, 12), 1203 => to_unsigned(3659, 12), 1204 => to_unsigned(963, 12), 1205 => to_unsigned(2631, 12), 1206 => to_unsigned(117, 12), 1207 => to_unsigned(3107, 12), 1208 => to_unsigned(1403, 12), 1209 => to_unsigned(1409, 12), 1210 => to_unsigned(1839, 12), 1211 => to_unsigned(2268, 12), 1212 => to_unsigned(3867, 12), 1213 => to_unsigned(2643, 12), 1214 => to_unsigned(1972, 12), 1215 => to_unsigned(3060, 12), 1216 => to_unsigned(1435, 12), 1217 => to_unsigned(758, 12), 1218 => to_unsigned(520, 12), 1219 => to_unsigned(684, 12), 1220 => to_unsigned(1805, 12), 1221 => to_unsigned(3970, 12), 1222 => to_unsigned(1337, 12), 1223 => to_unsigned(3643, 12), 1224 => to_unsigned(3893, 12), 1225 => to_unsigned(1758, 12), 1226 => to_unsigned(2603, 12), 1227 => to_unsigned(3738, 12), 1228 => to_unsigned(1528, 12), 1229 => to_unsigned(773, 12), 1230 => to_unsigned(3943, 12), 1231 => to_unsigned(3056, 12), 1232 => to_unsigned(2460, 12), 1233 => to_unsigned(281, 12), 1234 => to_unsigned(1619, 12), 1235 => to_unsigned(451, 12), 1236 => to_unsigned(994, 12), 1237 => to_unsigned(229, 12), 1238 => to_unsigned(2579, 12), 1239 => to_unsigned(3277, 12), 1240 => to_unsigned(1714, 12), 1241 => to_unsigned(3518, 12), 1242 => to_unsigned(621, 12), 1243 => to_unsigned(3476, 12), 1244 => to_unsigned(733, 12), 1245 => to_unsigned(3413, 12), 1246 => to_unsigned(1120, 12), 1247 => to_unsigned(3058, 12), 1248 => to_unsigned(896, 12), 1249 => to_unsigned(1219, 12), 1250 => to_unsigned(409, 12), 1251 => to_unsigned(507, 12), 1252 => to_unsigned(376, 12), 1253 => to_unsigned(703, 12), 1254 => to_unsigned(2640, 12), 1255 => to_unsigned(1891, 12), 1256 => to_unsigned(1329, 12), 1257 => to_unsigned(579, 12), 1258 => to_unsigned(1731, 12), 1259 => to_unsigned(1736, 12), 1260 => to_unsigned(2421, 12), 1261 => to_unsigned(1696, 12), 1262 => to_unsigned(3690, 12), 1263 => to_unsigned(3448, 12), 1264 => to_unsigned(1999, 12), 1265 => to_unsigned(4049, 12), 1266 => to_unsigned(2007, 12), 1267 => to_unsigned(2915, 12), 1268 => to_unsigned(184, 12), 1269 => to_unsigned(1849, 12), 1270 => to_unsigned(3217, 12), 1271 => to_unsigned(3355, 12), 1272 => to_unsigned(3903, 12), 1273 => to_unsigned(2108, 12), 1274 => to_unsigned(2426, 12), 1275 => to_unsigned(2324, 12), 1276 => to_unsigned(1596, 12), 1277 => to_unsigned(1946, 12), 1278 => to_unsigned(2869, 12), 1279 => to_unsigned(1038, 12), 1280 => to_unsigned(2462, 12), 1281 => to_unsigned(945, 12), 1282 => to_unsigned(3307, 12), 1283 => to_unsigned(3222, 12), 1284 => to_unsigned(3073, 12), 1285 => to_unsigned(953, 12), 1286 => to_unsigned(1053, 12), 1287 => to_unsigned(1965, 12), 1288 => to_unsigned(118, 12), 1289 => to_unsigned(3995, 12), 1290 => to_unsigned(485, 12), 1291 => to_unsigned(2952, 12), 1292 => to_unsigned(157, 12), 1293 => to_unsigned(419, 12), 1294 => to_unsigned(1917, 12), 1295 => to_unsigned(3498, 12), 1296 => to_unsigned(2010, 12), 1297 => to_unsigned(2090, 12), 1298 => to_unsigned(3113, 12), 1299 => to_unsigned(592, 12), 1300 => to_unsigned(343, 12), 1301 => to_unsigned(911, 12), 1302 => to_unsigned(1849, 12), 1303 => to_unsigned(3151, 12), 1304 => to_unsigned(1959, 12), 1305 => to_unsigned(1940, 12), 1306 => to_unsigned(3947, 12), 1307 => to_unsigned(2415, 12), 1308 => to_unsigned(2473, 12), 1309 => to_unsigned(2476, 12), 1310 => to_unsigned(3146, 12), 1311 => to_unsigned(886, 12), 1312 => to_unsigned(331, 12), 1313 => to_unsigned(2684, 12), 1314 => to_unsigned(2539, 12), 1315 => to_unsigned(2702, 12), 1316 => to_unsigned(217, 12), 1317 => to_unsigned(971, 12), 1318 => to_unsigned(1101, 12), 1319 => to_unsigned(4025, 12), 1320 => to_unsigned(691, 12), 1321 => to_unsigned(3588, 12), 1322 => to_unsigned(1634, 12), 1323 => to_unsigned(831, 12), 1324 => to_unsigned(322, 12), 1325 => to_unsigned(3605, 12), 1326 => to_unsigned(3372, 12), 1327 => to_unsigned(3124, 12), 1328 => to_unsigned(1134, 12), 1329 => to_unsigned(2898, 12), 1330 => to_unsigned(3315, 12), 1331 => to_unsigned(2971, 12), 1332 => to_unsigned(521, 12), 1333 => to_unsigned(1329, 12), 1334 => to_unsigned(3029, 12), 1335 => to_unsigned(4092, 12), 1336 => to_unsigned(2745, 12), 1337 => to_unsigned(863, 12), 1338 => to_unsigned(3091, 12), 1339 => to_unsigned(1629, 12), 1340 => to_unsigned(1469, 12), 1341 => to_unsigned(3449, 12), 1342 => to_unsigned(2261, 12), 1343 => to_unsigned(3927, 12), 1344 => to_unsigned(166, 12), 1345 => to_unsigned(2002, 12), 1346 => to_unsigned(141, 12), 1347 => to_unsigned(1736, 12), 1348 => to_unsigned(706, 12), 1349 => to_unsigned(3104, 12), 1350 => to_unsigned(3972, 12), 1351 => to_unsigned(2565, 12), 1352 => to_unsigned(3367, 12), 1353 => to_unsigned(2858, 12), 1354 => to_unsigned(1871, 12), 1355 => to_unsigned(50, 12), 1356 => to_unsigned(623, 12), 1357 => to_unsigned(354, 12), 1358 => to_unsigned(3658, 12), 1359 => to_unsigned(3178, 12), 1360 => to_unsigned(3202, 12), 1361 => to_unsigned(3184, 12), 1362 => to_unsigned(3225, 12), 1363 => to_unsigned(2466, 12), 1364 => to_unsigned(3650, 12), 1365 => to_unsigned(139, 12), 1366 => to_unsigned(675, 12), 1367 => to_unsigned(2795, 12), 1368 => to_unsigned(3648, 12), 1369 => to_unsigned(1211, 12), 1370 => to_unsigned(488, 12), 1371 => to_unsigned(3943, 12), 1372 => to_unsigned(3888, 12), 1373 => to_unsigned(2116, 12), 1374 => to_unsigned(673, 12), 1375 => to_unsigned(3145, 12), 1376 => to_unsigned(1542, 12), 1377 => to_unsigned(2297, 12), 1378 => to_unsigned(922, 12), 1379 => to_unsigned(2179, 12), 1380 => to_unsigned(767, 12), 1381 => to_unsigned(1186, 12), 1382 => to_unsigned(2892, 12), 1383 => to_unsigned(3232, 12), 1384 => to_unsigned(1955, 12), 1385 => to_unsigned(3619, 12), 1386 => to_unsigned(1277, 12), 1387 => to_unsigned(536, 12), 1388 => to_unsigned(1459, 12), 1389 => to_unsigned(121, 12), 1390 => to_unsigned(3986, 12), 1391 => to_unsigned(3171, 12), 1392 => to_unsigned(1449, 12), 1393 => to_unsigned(3687, 12), 1394 => to_unsigned(2214, 12), 1395 => to_unsigned(3735, 12), 1396 => to_unsigned(1372, 12), 1397 => to_unsigned(1720, 12), 1398 => to_unsigned(4091, 12), 1399 => to_unsigned(2042, 12), 1400 => to_unsigned(266, 12), 1401 => to_unsigned(2214, 12), 1402 => to_unsigned(2804, 12), 1403 => to_unsigned(3398, 12), 1404 => to_unsigned(1653, 12), 1405 => to_unsigned(49, 12), 1406 => to_unsigned(835, 12), 1407 => to_unsigned(1368, 12), 1408 => to_unsigned(2827, 12), 1409 => to_unsigned(2844, 12), 1410 => to_unsigned(3252, 12), 1411 => to_unsigned(349, 12), 1412 => to_unsigned(3166, 12), 1413 => to_unsigned(2493, 12), 1414 => to_unsigned(3852, 12), 1415 => to_unsigned(307, 12), 1416 => to_unsigned(2110, 12), 1417 => to_unsigned(919, 12), 1418 => to_unsigned(2342, 12), 1419 => to_unsigned(1533, 12), 1420 => to_unsigned(2847, 12), 1421 => to_unsigned(769, 12), 1422 => to_unsigned(2536, 12), 1423 => to_unsigned(2552, 12), 1424 => to_unsigned(2363, 12), 1425 => to_unsigned(3516, 12), 1426 => to_unsigned(2423, 12), 1427 => to_unsigned(693, 12), 1428 => to_unsigned(2163, 12), 1429 => to_unsigned(1117, 12), 1430 => to_unsigned(4016, 12), 1431 => to_unsigned(679, 12), 1432 => to_unsigned(362, 12), 1433 => to_unsigned(377, 12), 1434 => to_unsigned(3811, 12), 1435 => to_unsigned(1513, 12), 1436 => to_unsigned(805, 12), 1437 => to_unsigned(2141, 12), 1438 => to_unsigned(3097, 12), 1439 => to_unsigned(4005, 12), 1440 => to_unsigned(1141, 12), 1441 => to_unsigned(3502, 12), 1442 => to_unsigned(1332, 12), 1443 => to_unsigned(1884, 12), 1444 => to_unsigned(3674, 12), 1445 => to_unsigned(1955, 12), 1446 => to_unsigned(1318, 12), 1447 => to_unsigned(2163, 12), 1448 => to_unsigned(256, 12), 1449 => to_unsigned(1946, 12), 1450 => to_unsigned(1390, 12), 1451 => to_unsigned(623, 12), 1452 => to_unsigned(3182, 12), 1453 => to_unsigned(2485, 12), 1454 => to_unsigned(3396, 12), 1455 => to_unsigned(3775, 12), 1456 => to_unsigned(1822, 12), 1457 => to_unsigned(3980, 12), 1458 => to_unsigned(202, 12), 1459 => to_unsigned(832, 12), 1460 => to_unsigned(2494, 12), 1461 => to_unsigned(1965, 12), 1462 => to_unsigned(2323, 12), 1463 => to_unsigned(433, 12), 1464 => to_unsigned(1976, 12), 1465 => to_unsigned(3712, 12), 1466 => to_unsigned(703, 12), 1467 => to_unsigned(373, 12), 1468 => to_unsigned(480, 12), 1469 => to_unsigned(1427, 12), 1470 => to_unsigned(806, 12), 1471 => to_unsigned(1333, 12), 1472 => to_unsigned(615, 12), 1473 => to_unsigned(1943, 12), 1474 => to_unsigned(3502, 12), 1475 => to_unsigned(2682, 12), 1476 => to_unsigned(3920, 12), 1477 => to_unsigned(756, 12), 1478 => to_unsigned(3826, 12), 1479 => to_unsigned(112, 12), 1480 => to_unsigned(2650, 12), 1481 => to_unsigned(1469, 12), 1482 => to_unsigned(72, 12), 1483 => to_unsigned(924, 12), 1484 => to_unsigned(3606, 12), 1485 => to_unsigned(4007, 12), 1486 => to_unsigned(226, 12), 1487 => to_unsigned(310, 12), 1488 => to_unsigned(1359, 12), 1489 => to_unsigned(1095, 12), 1490 => to_unsigned(1601, 12), 1491 => to_unsigned(3868, 12), 1492 => to_unsigned(1850, 12), 1493 => to_unsigned(322, 12), 1494 => to_unsigned(2440, 12), 1495 => to_unsigned(3961, 12), 1496 => to_unsigned(303, 12), 1497 => to_unsigned(2715, 12), 1498 => to_unsigned(1427, 12), 1499 => to_unsigned(228, 12), 1500 => to_unsigned(1490, 12), 1501 => to_unsigned(1958, 12), 1502 => to_unsigned(3491, 12), 1503 => to_unsigned(3567, 12), 1504 => to_unsigned(2544, 12), 1505 => to_unsigned(938, 12), 1506 => to_unsigned(3320, 12), 1507 => to_unsigned(3199, 12), 1508 => to_unsigned(2055, 12), 1509 => to_unsigned(4086, 12), 1510 => to_unsigned(3696, 12), 1511 => to_unsigned(621, 12), 1512 => to_unsigned(880, 12), 1513 => to_unsigned(1764, 12), 1514 => to_unsigned(1846, 12), 1515 => to_unsigned(1789, 12), 1516 => to_unsigned(3167, 12), 1517 => to_unsigned(2564, 12), 1518 => to_unsigned(2501, 12), 1519 => to_unsigned(3463, 12), 1520 => to_unsigned(279, 12), 1521 => to_unsigned(948, 12), 1522 => to_unsigned(220, 12), 1523 => to_unsigned(313, 12), 1524 => to_unsigned(3650, 12), 1525 => to_unsigned(3844, 12), 1526 => to_unsigned(3396, 12), 1527 => to_unsigned(1498, 12), 1528 => to_unsigned(3597, 12), 1529 => to_unsigned(1562, 12), 1530 => to_unsigned(3308, 12), 1531 => to_unsigned(2689, 12), 1532 => to_unsigned(1558, 12), 1533 => to_unsigned(1078, 12), 1534 => to_unsigned(762, 12), 1535 => to_unsigned(2094, 12), 1536 => to_unsigned(2632, 12), 1537 => to_unsigned(2053, 12), 1538 => to_unsigned(2244, 12), 1539 => to_unsigned(3837, 12), 1540 => to_unsigned(2700, 12), 1541 => to_unsigned(402, 12), 1542 => to_unsigned(3566, 12), 1543 => to_unsigned(2785, 12), 1544 => to_unsigned(2178, 12), 1545 => to_unsigned(1373, 12), 1546 => to_unsigned(1471, 12), 1547 => to_unsigned(1327, 12), 1548 => to_unsigned(3417, 12), 1549 => to_unsigned(3746, 12), 1550 => to_unsigned(2490, 12), 1551 => to_unsigned(1173, 12), 1552 => to_unsigned(2940, 12), 1553 => to_unsigned(4040, 12), 1554 => to_unsigned(3601, 12), 1555 => to_unsigned(922, 12), 1556 => to_unsigned(760, 12), 1557 => to_unsigned(2276, 12), 1558 => to_unsigned(107, 12), 1559 => to_unsigned(157, 12), 1560 => to_unsigned(2428, 12), 1561 => to_unsigned(2507, 12), 1562 => to_unsigned(224, 12), 1563 => to_unsigned(2135, 12), 1564 => to_unsigned(1107, 12), 1565 => to_unsigned(768, 12), 1566 => to_unsigned(1813, 12), 1567 => to_unsigned(668, 12), 1568 => to_unsigned(289, 12), 1569 => to_unsigned(1206, 12), 1570 => to_unsigned(1003, 12), 1571 => to_unsigned(2813, 12), 1572 => to_unsigned(3218, 12), 1573 => to_unsigned(256, 12), 1574 => to_unsigned(2086, 12), 1575 => to_unsigned(2898, 12), 1576 => to_unsigned(1970, 12), 1577 => to_unsigned(986, 12), 1578 => to_unsigned(1869, 12), 1579 => to_unsigned(2739, 12), 1580 => to_unsigned(2755, 12), 1581 => to_unsigned(3841, 12), 1582 => to_unsigned(167, 12), 1583 => to_unsigned(3991, 12), 1584 => to_unsigned(3244, 12), 1585 => to_unsigned(415, 12), 1586 => to_unsigned(1031, 12), 1587 => to_unsigned(158, 12), 1588 => to_unsigned(1398, 12), 1589 => to_unsigned(540, 12), 1590 => to_unsigned(182, 12), 1591 => to_unsigned(3376, 12), 1592 => to_unsigned(1800, 12), 1593 => to_unsigned(218, 12), 1594 => to_unsigned(133, 12), 1595 => to_unsigned(3845, 12), 1596 => to_unsigned(3317, 12), 1597 => to_unsigned(1059, 12), 1598 => to_unsigned(1434, 12), 1599 => to_unsigned(3187, 12), 1600 => to_unsigned(2100, 12), 1601 => to_unsigned(869, 12), 1602 => to_unsigned(2128, 12), 1603 => to_unsigned(441, 12), 1604 => to_unsigned(1909, 12), 1605 => to_unsigned(995, 12), 1606 => to_unsigned(744, 12), 1607 => to_unsigned(2572, 12), 1608 => to_unsigned(924, 12), 1609 => to_unsigned(2821, 12), 1610 => to_unsigned(2818, 12), 1611 => to_unsigned(50, 12), 1612 => to_unsigned(1876, 12), 1613 => to_unsigned(2232, 12), 1614 => to_unsigned(3326, 12), 1615 => to_unsigned(2830, 12), 1616 => to_unsigned(1105, 12), 1617 => to_unsigned(90, 12), 1618 => to_unsigned(3700, 12), 1619 => to_unsigned(2308, 12), 1620 => to_unsigned(174, 12), 1621 => to_unsigned(520, 12), 1622 => to_unsigned(3272, 12), 1623 => to_unsigned(531, 12), 1624 => to_unsigned(15, 12), 1625 => to_unsigned(1171, 12), 1626 => to_unsigned(3442, 12), 1627 => to_unsigned(1654, 12), 1628 => to_unsigned(530, 12), 1629 => to_unsigned(1881, 12), 1630 => to_unsigned(485, 12), 1631 => to_unsigned(1486, 12), 1632 => to_unsigned(2712, 12), 1633 => to_unsigned(446, 12), 1634 => to_unsigned(1276, 12), 1635 => to_unsigned(453, 12), 1636 => to_unsigned(1586, 12), 1637 => to_unsigned(2057, 12), 1638 => to_unsigned(1051, 12), 1639 => to_unsigned(2138, 12), 1640 => to_unsigned(3791, 12), 1641 => to_unsigned(3875, 12), 1642 => to_unsigned(717, 12), 1643 => to_unsigned(3850, 12), 1644 => to_unsigned(3595, 12), 1645 => to_unsigned(99, 12), 1646 => to_unsigned(1038, 12), 1647 => to_unsigned(242, 12), 1648 => to_unsigned(1472, 12), 1649 => to_unsigned(1481, 12), 1650 => to_unsigned(3506, 12), 1651 => to_unsigned(1983, 12), 1652 => to_unsigned(3437, 12), 1653 => to_unsigned(577, 12), 1654 => to_unsigned(2244, 12), 1655 => to_unsigned(4057, 12), 1656 => to_unsigned(3739, 12), 1657 => to_unsigned(3381, 12), 1658 => to_unsigned(2357, 12), 1659 => to_unsigned(4092, 12), 1660 => to_unsigned(100, 12), 1661 => to_unsigned(3283, 12), 1662 => to_unsigned(2829, 12), 1663 => to_unsigned(1496, 12), 1664 => to_unsigned(1009, 12), 1665 => to_unsigned(175, 12), 1666 => to_unsigned(1684, 12), 1667 => to_unsigned(384, 12), 1668 => to_unsigned(1888, 12), 1669 => to_unsigned(3112, 12), 1670 => to_unsigned(3550, 12), 1671 => to_unsigned(2914, 12), 1672 => to_unsigned(1189, 12), 1673 => to_unsigned(3812, 12), 1674 => to_unsigned(3561, 12), 1675 => to_unsigned(2158, 12), 1676 => to_unsigned(548, 12), 1677 => to_unsigned(482, 12), 1678 => to_unsigned(3216, 12), 1679 => to_unsigned(612, 12), 1680 => to_unsigned(3383, 12), 1681 => to_unsigned(1925, 12), 1682 => to_unsigned(1369, 12), 1683 => to_unsigned(3576, 12), 1684 => to_unsigned(625, 12), 1685 => to_unsigned(1793, 12), 1686 => to_unsigned(2047, 12), 1687 => to_unsigned(3862, 12), 1688 => to_unsigned(3927, 12), 1689 => to_unsigned(1228, 12), 1690 => to_unsigned(3912, 12), 1691 => to_unsigned(1337, 12), 1692 => to_unsigned(2468, 12), 1693 => to_unsigned(2518, 12), 1694 => to_unsigned(3562, 12), 1695 => to_unsigned(433, 12), 1696 => to_unsigned(1180, 12), 1697 => to_unsigned(390, 12), 1698 => to_unsigned(142, 12), 1699 => to_unsigned(2607, 12), 1700 => to_unsigned(2547, 12), 1701 => to_unsigned(2268, 12), 1702 => to_unsigned(1141, 12), 1703 => to_unsigned(2061, 12), 1704 => to_unsigned(1506, 12), 1705 => to_unsigned(3391, 12), 1706 => to_unsigned(501, 12), 1707 => to_unsigned(3398, 12), 1708 => to_unsigned(3550, 12), 1709 => to_unsigned(1802, 12), 1710 => to_unsigned(3712, 12), 1711 => to_unsigned(2872, 12), 1712 => to_unsigned(3719, 12), 1713 => to_unsigned(770, 12), 1714 => to_unsigned(1306, 12), 1715 => to_unsigned(592, 12), 1716 => to_unsigned(869, 12), 1717 => to_unsigned(3266, 12), 1718 => to_unsigned(2989, 12), 1719 => to_unsigned(1119, 12), 1720 => to_unsigned(1396, 12), 1721 => to_unsigned(1155, 12), 1722 => to_unsigned(2789, 12), 1723 => to_unsigned(2497, 12), 1724 => to_unsigned(879, 12), 1725 => to_unsigned(37, 12), 1726 => to_unsigned(2170, 12), 1727 => to_unsigned(1549, 12), 1728 => to_unsigned(3772, 12), 1729 => to_unsigned(447, 12), 1730 => to_unsigned(2245, 12), 1731 => to_unsigned(3346, 12), 1732 => to_unsigned(3887, 12), 1733 => to_unsigned(2593, 12), 1734 => to_unsigned(1239, 12), 1735 => to_unsigned(2548, 12), 1736 => to_unsigned(4002, 12), 1737 => to_unsigned(3562, 12), 1738 => to_unsigned(65, 12), 1739 => to_unsigned(1394, 12), 1740 => to_unsigned(3119, 12), 1741 => to_unsigned(2398, 12), 1742 => to_unsigned(2196, 12), 1743 => to_unsigned(3224, 12), 1744 => to_unsigned(2575, 12), 1745 => to_unsigned(1472, 12), 1746 => to_unsigned(403, 12), 1747 => to_unsigned(3716, 12), 1748 => to_unsigned(1800, 12), 1749 => to_unsigned(3330, 12), 1750 => to_unsigned(2715, 12), 1751 => to_unsigned(3201, 12), 1752 => to_unsigned(60, 12), 1753 => to_unsigned(1407, 12), 1754 => to_unsigned(2339, 12), 1755 => to_unsigned(3228, 12), 1756 => to_unsigned(3052, 12), 1757 => to_unsigned(2087, 12), 1758 => to_unsigned(784, 12), 1759 => to_unsigned(2599, 12), 1760 => to_unsigned(1141, 12), 1761 => to_unsigned(2986, 12), 1762 => to_unsigned(1329, 12), 1763 => to_unsigned(1797, 12), 1764 => to_unsigned(2113, 12), 1765 => to_unsigned(4074, 12), 1766 => to_unsigned(1629, 12), 1767 => to_unsigned(2639, 12), 1768 => to_unsigned(3570, 12), 1769 => to_unsigned(349, 12), 1770 => to_unsigned(2266, 12), 1771 => to_unsigned(354, 12), 1772 => to_unsigned(3572, 12), 1773 => to_unsigned(2802, 12), 1774 => to_unsigned(2773, 12), 1775 => to_unsigned(1108, 12), 1776 => to_unsigned(3639, 12), 1777 => to_unsigned(346, 12), 1778 => to_unsigned(357, 12), 1779 => to_unsigned(2712, 12), 1780 => to_unsigned(1053, 12), 1781 => to_unsigned(305, 12), 1782 => to_unsigned(1212, 12), 1783 => to_unsigned(948, 12), 1784 => to_unsigned(2654, 12), 1785 => to_unsigned(2815, 12), 1786 => to_unsigned(3280, 12), 1787 => to_unsigned(3276, 12), 1788 => to_unsigned(3691, 12), 1789 => to_unsigned(2635, 12), 1790 => to_unsigned(2194, 12), 1791 => to_unsigned(830, 12), 1792 => to_unsigned(486, 12), 1793 => to_unsigned(2786, 12), 1794 => to_unsigned(2707, 12), 1795 => to_unsigned(1609, 12), 1796 => to_unsigned(2592, 12), 1797 => to_unsigned(2060, 12), 1798 => to_unsigned(3627, 12), 1799 => to_unsigned(2066, 12), 1800 => to_unsigned(323, 12), 1801 => to_unsigned(3947, 12), 1802 => to_unsigned(1198, 12), 1803 => to_unsigned(2676, 12), 1804 => to_unsigned(1540, 12), 1805 => to_unsigned(779, 12), 1806 => to_unsigned(1668, 12), 1807 => to_unsigned(2711, 12), 1808 => to_unsigned(2745, 12), 1809 => to_unsigned(3289, 12), 1810 => to_unsigned(1581, 12), 1811 => to_unsigned(1050, 12), 1812 => to_unsigned(2497, 12), 1813 => to_unsigned(3462, 12), 1814 => to_unsigned(2773, 12), 1815 => to_unsigned(1748, 12), 1816 => to_unsigned(990, 12), 1817 => to_unsigned(2531, 12), 1818 => to_unsigned(1374, 12), 1819 => to_unsigned(3592, 12), 1820 => to_unsigned(2872, 12), 1821 => to_unsigned(2315, 12), 1822 => to_unsigned(189, 12), 1823 => to_unsigned(3492, 12), 1824 => to_unsigned(2674, 12), 1825 => to_unsigned(1726, 12), 1826 => to_unsigned(2178, 12), 1827 => to_unsigned(1643, 12), 1828 => to_unsigned(719, 12), 1829 => to_unsigned(1774, 12), 1830 => to_unsigned(3401, 12), 1831 => to_unsigned(3656, 12), 1832 => to_unsigned(963, 12), 1833 => to_unsigned(3924, 12), 1834 => to_unsigned(665, 12), 1835 => to_unsigned(1077, 12), 1836 => to_unsigned(1408, 12), 1837 => to_unsigned(329, 12), 1838 => to_unsigned(2610, 12), 1839 => to_unsigned(1668, 12), 1840 => to_unsigned(70, 12), 1841 => to_unsigned(1610, 12), 1842 => to_unsigned(650, 12), 1843 => to_unsigned(800, 12), 1844 => to_unsigned(114, 12), 1845 => to_unsigned(3495, 12), 1846 => to_unsigned(2430, 12), 1847 => to_unsigned(2307, 12), 1848 => to_unsigned(2005, 12), 1849 => to_unsigned(3708, 12), 1850 => to_unsigned(1235, 12), 1851 => to_unsigned(1677, 12), 1852 => to_unsigned(3861, 12), 1853 => to_unsigned(2676, 12), 1854 => to_unsigned(2824, 12), 1855 => to_unsigned(252, 12), 1856 => to_unsigned(1994, 12), 1857 => to_unsigned(1338, 12), 1858 => to_unsigned(1322, 12), 1859 => to_unsigned(2589, 12), 1860 => to_unsigned(605, 12), 1861 => to_unsigned(231, 12), 1862 => to_unsigned(2562, 12), 1863 => to_unsigned(2560, 12), 1864 => to_unsigned(652, 12), 1865 => to_unsigned(2746, 12), 1866 => to_unsigned(524, 12), 1867 => to_unsigned(1994, 12), 1868 => to_unsigned(2576, 12), 1869 => to_unsigned(742, 12), 1870 => to_unsigned(1881, 12), 1871 => to_unsigned(1947, 12), 1872 => to_unsigned(733, 12), 1873 => to_unsigned(1345, 12), 1874 => to_unsigned(496, 12), 1875 => to_unsigned(1029, 12), 1876 => to_unsigned(604, 12), 1877 => to_unsigned(2578, 12), 1878 => to_unsigned(348, 12), 1879 => to_unsigned(3522, 12), 1880 => to_unsigned(141, 12), 1881 => to_unsigned(1746, 12), 1882 => to_unsigned(707, 12), 1883 => to_unsigned(716, 12), 1884 => to_unsigned(1557, 12), 1885 => to_unsigned(1161, 12), 1886 => to_unsigned(2525, 12), 1887 => to_unsigned(1148, 12), 1888 => to_unsigned(3799, 12), 1889 => to_unsigned(3873, 12), 1890 => to_unsigned(3400, 12), 1891 => to_unsigned(1031, 12), 1892 => to_unsigned(1373, 12), 1893 => to_unsigned(137, 12), 1894 => to_unsigned(3315, 12), 1895 => to_unsigned(2736, 12), 1896 => to_unsigned(243, 12), 1897 => to_unsigned(2463, 12), 1898 => to_unsigned(1819, 12), 1899 => to_unsigned(1785, 12), 1900 => to_unsigned(3950, 12), 1901 => to_unsigned(3108, 12), 1902 => to_unsigned(1854, 12), 1903 => to_unsigned(3761, 12), 1904 => to_unsigned(3915, 12), 1905 => to_unsigned(1902, 12), 1906 => to_unsigned(3782, 12), 1907 => to_unsigned(2973, 12), 1908 => to_unsigned(637, 12), 1909 => to_unsigned(3337, 12), 1910 => to_unsigned(14, 12), 1911 => to_unsigned(1972, 12), 1912 => to_unsigned(2142, 12), 1913 => to_unsigned(1654, 12), 1914 => to_unsigned(3771, 12), 1915 => to_unsigned(1881, 12), 1916 => to_unsigned(4, 12), 1917 => to_unsigned(3134, 12), 1918 => to_unsigned(1049, 12), 1919 => to_unsigned(2110, 12), 1920 => to_unsigned(2257, 12), 1921 => to_unsigned(1811, 12), 1922 => to_unsigned(1647, 12), 1923 => to_unsigned(2091, 12), 1924 => to_unsigned(4077, 12), 1925 => to_unsigned(3600, 12), 1926 => to_unsigned(2528, 12), 1927 => to_unsigned(254, 12), 1928 => to_unsigned(3735, 12), 1929 => to_unsigned(929, 12), 1930 => to_unsigned(616, 12), 1931 => to_unsigned(3223, 12), 1932 => to_unsigned(2175, 12), 1933 => to_unsigned(2706, 12), 1934 => to_unsigned(189, 12), 1935 => to_unsigned(109, 12), 1936 => to_unsigned(2157, 12), 1937 => to_unsigned(2785, 12), 1938 => to_unsigned(2724, 12), 1939 => to_unsigned(4049, 12), 1940 => to_unsigned(132, 12), 1941 => to_unsigned(3225, 12), 1942 => to_unsigned(3412, 12), 1943 => to_unsigned(1464, 12), 1944 => to_unsigned(1510, 12), 1945 => to_unsigned(359, 12), 1946 => to_unsigned(2046, 12), 1947 => to_unsigned(968, 12), 1948 => to_unsigned(4094, 12), 1949 => to_unsigned(419, 12), 1950 => to_unsigned(3725, 12), 1951 => to_unsigned(3701, 12), 1952 => to_unsigned(1446, 12), 1953 => to_unsigned(1815, 12), 1954 => to_unsigned(3354, 12), 1955 => to_unsigned(2504, 12), 1956 => to_unsigned(467, 12), 1957 => to_unsigned(480, 12), 1958 => to_unsigned(757, 12), 1959 => to_unsigned(3844, 12), 1960 => to_unsigned(3617, 12), 1961 => to_unsigned(1495, 12), 1962 => to_unsigned(1457, 12), 1963 => to_unsigned(4007, 12), 1964 => to_unsigned(3796, 12), 1965 => to_unsigned(1424, 12), 1966 => to_unsigned(2024, 12), 1967 => to_unsigned(2719, 12), 1968 => to_unsigned(2553, 12), 1969 => to_unsigned(1847, 12), 1970 => to_unsigned(15, 12), 1971 => to_unsigned(227, 12), 1972 => to_unsigned(1401, 12), 1973 => to_unsigned(900, 12), 1974 => to_unsigned(3726, 12), 1975 => to_unsigned(68, 12), 1976 => to_unsigned(3891, 12), 1977 => to_unsigned(672, 12), 1978 => to_unsigned(387, 12), 1979 => to_unsigned(935, 12), 1980 => to_unsigned(1205, 12), 1981 => to_unsigned(2503, 12), 1982 => to_unsigned(2614, 12), 1983 => to_unsigned(920, 12), 1984 => to_unsigned(827, 12), 1985 => to_unsigned(1018, 12), 1986 => to_unsigned(3890, 12), 1987 => to_unsigned(4065, 12), 1988 => to_unsigned(2729, 12), 1989 => to_unsigned(587, 12), 1990 => to_unsigned(3026, 12), 1991 => to_unsigned(710, 12), 1992 => to_unsigned(2052, 12), 1993 => to_unsigned(1085, 12), 1994 => to_unsigned(343, 12), 1995 => to_unsigned(215, 12), 1996 => to_unsigned(1180, 12), 1997 => to_unsigned(3590, 12), 1998 => to_unsigned(3730, 12), 1999 => to_unsigned(2498, 12), 2000 => to_unsigned(822, 12), 2001 => to_unsigned(2050, 12), 2002 => to_unsigned(868, 12), 2003 => to_unsigned(1139, 12), 2004 => to_unsigned(3497, 12), 2005 => to_unsigned(2812, 12), 2006 => to_unsigned(100, 12), 2007 => to_unsigned(1119, 12), 2008 => to_unsigned(1472, 12), 2009 => to_unsigned(3453, 12), 2010 => to_unsigned(732, 12), 2011 => to_unsigned(42, 12), 2012 => to_unsigned(265, 12), 2013 => to_unsigned(3885, 12), 2014 => to_unsigned(3667, 12), 2015 => to_unsigned(431, 12), 2016 => to_unsigned(649, 12), 2017 => to_unsigned(3310, 12), 2018 => to_unsigned(15, 12), 2019 => to_unsigned(3197, 12), 2020 => to_unsigned(615, 12), 2021 => to_unsigned(3900, 12), 2022 => to_unsigned(2440, 12), 2023 => to_unsigned(3193, 12), 2024 => to_unsigned(2789, 12), 2025 => to_unsigned(3005, 12), 2026 => to_unsigned(3815, 12), 2027 => to_unsigned(2148, 12), 2028 => to_unsigned(3332, 12), 2029 => to_unsigned(3852, 12), 2030 => to_unsigned(3120, 12), 2031 => to_unsigned(1566, 12), 2032 => to_unsigned(758, 12), 2033 => to_unsigned(3518, 12), 2034 => to_unsigned(300, 12), 2035 => to_unsigned(833, 12), 2036 => to_unsigned(2760, 12), 2037 => to_unsigned(3569, 12), 2038 => to_unsigned(1979, 12), 2039 => to_unsigned(3178, 12), 2040 => to_unsigned(3931, 12), 2041 => to_unsigned(2554, 12), 2042 => to_unsigned(3995, 12), 2043 => to_unsigned(1568, 12), 2044 => to_unsigned(4055, 12), 2045 => to_unsigned(3634, 12), 2046 => to_unsigned(3944, 12), 2047 => to_unsigned(3813, 12)),
            7 => (0 => to_unsigned(143, 12), 1 => to_unsigned(1166, 12), 2 => to_unsigned(82, 12), 3 => to_unsigned(4049, 12), 4 => to_unsigned(2528, 12), 5 => to_unsigned(3747, 12), 6 => to_unsigned(3629, 12), 7 => to_unsigned(3358, 12), 8 => to_unsigned(3453, 12), 9 => to_unsigned(985, 12), 10 => to_unsigned(11, 12), 11 => to_unsigned(1607, 12), 12 => to_unsigned(2881, 12), 13 => to_unsigned(3301, 12), 14 => to_unsigned(466, 12), 15 => to_unsigned(562, 12), 16 => to_unsigned(3504, 12), 17 => to_unsigned(1636, 12), 18 => to_unsigned(2982, 12), 19 => to_unsigned(731, 12), 20 => to_unsigned(1531, 12), 21 => to_unsigned(2208, 12), 22 => to_unsigned(3227, 12), 23 => to_unsigned(1051, 12), 24 => to_unsigned(3302, 12), 25 => to_unsigned(2926, 12), 26 => to_unsigned(1658, 12), 27 => to_unsigned(979, 12), 28 => to_unsigned(1668, 12), 29 => to_unsigned(1263, 12), 30 => to_unsigned(440, 12), 31 => to_unsigned(2860, 12), 32 => to_unsigned(3944, 12), 33 => to_unsigned(2124, 12), 34 => to_unsigned(3623, 12), 35 => to_unsigned(3054, 12), 36 => to_unsigned(3688, 12), 37 => to_unsigned(1251, 12), 38 => to_unsigned(3843, 12), 39 => to_unsigned(1028, 12), 40 => to_unsigned(3820, 12), 41 => to_unsigned(3111, 12), 42 => to_unsigned(1581, 12), 43 => to_unsigned(3887, 12), 44 => to_unsigned(3062, 12), 45 => to_unsigned(3571, 12), 46 => to_unsigned(2714, 12), 47 => to_unsigned(1219, 12), 48 => to_unsigned(3607, 12), 49 => to_unsigned(892, 12), 50 => to_unsigned(4067, 12), 51 => to_unsigned(2003, 12), 52 => to_unsigned(1054, 12), 53 => to_unsigned(1725, 12), 54 => to_unsigned(1135, 12), 55 => to_unsigned(2694, 12), 56 => to_unsigned(3565, 12), 57 => to_unsigned(1195, 12), 58 => to_unsigned(1760, 12), 59 => to_unsigned(1759, 12), 60 => to_unsigned(2880, 12), 61 => to_unsigned(1341, 12), 62 => to_unsigned(305, 12), 63 => to_unsigned(1916, 12), 64 => to_unsigned(3813, 12), 65 => to_unsigned(433, 12), 66 => to_unsigned(3255, 12), 67 => to_unsigned(2309, 12), 68 => to_unsigned(3386, 12), 69 => to_unsigned(906, 12), 70 => to_unsigned(1297, 12), 71 => to_unsigned(1273, 12), 72 => to_unsigned(3257, 12), 73 => to_unsigned(1146, 12), 74 => to_unsigned(1897, 12), 75 => to_unsigned(3522, 12), 76 => to_unsigned(3904, 12), 77 => to_unsigned(514, 12), 78 => to_unsigned(152, 12), 79 => to_unsigned(3052, 12), 80 => to_unsigned(3928, 12), 81 => to_unsigned(2537, 12), 82 => to_unsigned(311, 12), 83 => to_unsigned(1706, 12), 84 => to_unsigned(1976, 12), 85 => to_unsigned(2551, 12), 86 => to_unsigned(1242, 12), 87 => to_unsigned(755, 12), 88 => to_unsigned(2784, 12), 89 => to_unsigned(1902, 12), 90 => to_unsigned(953, 12), 91 => to_unsigned(1466, 12), 92 => to_unsigned(1688, 12), 93 => to_unsigned(3921, 12), 94 => to_unsigned(1454, 12), 95 => to_unsigned(2037, 12), 96 => to_unsigned(530, 12), 97 => to_unsigned(2191, 12), 98 => to_unsigned(1347, 12), 99 => to_unsigned(2757, 12), 100 => to_unsigned(1482, 12), 101 => to_unsigned(3939, 12), 102 => to_unsigned(2273, 12), 103 => to_unsigned(1666, 12), 104 => to_unsigned(881, 12), 105 => to_unsigned(3232, 12), 106 => to_unsigned(473, 12), 107 => to_unsigned(3317, 12), 108 => to_unsigned(536, 12), 109 => to_unsigned(1924, 12), 110 => to_unsigned(1541, 12), 111 => to_unsigned(1793, 12), 112 => to_unsigned(733, 12), 113 => to_unsigned(1018, 12), 114 => to_unsigned(2011, 12), 115 => to_unsigned(3253, 12), 116 => to_unsigned(2313, 12), 117 => to_unsigned(2785, 12), 118 => to_unsigned(4048, 12), 119 => to_unsigned(1938, 12), 120 => to_unsigned(2263, 12), 121 => to_unsigned(3711, 12), 122 => to_unsigned(1041, 12), 123 => to_unsigned(2256, 12), 124 => to_unsigned(1914, 12), 125 => to_unsigned(1637, 12), 126 => to_unsigned(3630, 12), 127 => to_unsigned(64, 12), 128 => to_unsigned(3469, 12), 129 => to_unsigned(3610, 12), 130 => to_unsigned(1339, 12), 131 => to_unsigned(2613, 12), 132 => to_unsigned(970, 12), 133 => to_unsigned(1578, 12), 134 => to_unsigned(3933, 12), 135 => to_unsigned(1305, 12), 136 => to_unsigned(1089, 12), 137 => to_unsigned(167, 12), 138 => to_unsigned(3323, 12), 139 => to_unsigned(2246, 12), 140 => to_unsigned(3229, 12), 141 => to_unsigned(3759, 12), 142 => to_unsigned(2459, 12), 143 => to_unsigned(2789, 12), 144 => to_unsigned(2880, 12), 145 => to_unsigned(1433, 12), 146 => to_unsigned(2908, 12), 147 => to_unsigned(1367, 12), 148 => to_unsigned(1154, 12), 149 => to_unsigned(1922, 12), 150 => to_unsigned(975, 12), 151 => to_unsigned(2331, 12), 152 => to_unsigned(2374, 12), 153 => to_unsigned(3809, 12), 154 => to_unsigned(3145, 12), 155 => to_unsigned(2217, 12), 156 => to_unsigned(192, 12), 157 => to_unsigned(3419, 12), 158 => to_unsigned(1013, 12), 159 => to_unsigned(3741, 12), 160 => to_unsigned(77, 12), 161 => to_unsigned(4085, 12), 162 => to_unsigned(3281, 12), 163 => to_unsigned(922, 12), 164 => to_unsigned(1600, 12), 165 => to_unsigned(1154, 12), 166 => to_unsigned(3052, 12), 167 => to_unsigned(1436, 12), 168 => to_unsigned(3958, 12), 169 => to_unsigned(1344, 12), 170 => to_unsigned(1671, 12), 171 => to_unsigned(1492, 12), 172 => to_unsigned(2944, 12), 173 => to_unsigned(1045, 12), 174 => to_unsigned(4076, 12), 175 => to_unsigned(162, 12), 176 => to_unsigned(573, 12), 177 => to_unsigned(3324, 12), 178 => to_unsigned(670, 12), 179 => to_unsigned(1754, 12), 180 => to_unsigned(3219, 12), 181 => to_unsigned(821, 12), 182 => to_unsigned(1957, 12), 183 => to_unsigned(3880, 12), 184 => to_unsigned(1011, 12), 185 => to_unsigned(849, 12), 186 => to_unsigned(2284, 12), 187 => to_unsigned(1988, 12), 188 => to_unsigned(3856, 12), 189 => to_unsigned(2194, 12), 190 => to_unsigned(1464, 12), 191 => to_unsigned(654, 12), 192 => to_unsigned(3027, 12), 193 => to_unsigned(1914, 12), 194 => to_unsigned(367, 12), 195 => to_unsigned(2807, 12), 196 => to_unsigned(3917, 12), 197 => to_unsigned(520, 12), 198 => to_unsigned(2215, 12), 199 => to_unsigned(3694, 12), 200 => to_unsigned(1264, 12), 201 => to_unsigned(3210, 12), 202 => to_unsigned(3237, 12), 203 => to_unsigned(2647, 12), 204 => to_unsigned(983, 12), 205 => to_unsigned(1518, 12), 206 => to_unsigned(3257, 12), 207 => to_unsigned(2237, 12), 208 => to_unsigned(2555, 12), 209 => to_unsigned(2223, 12), 210 => to_unsigned(1407, 12), 211 => to_unsigned(65, 12), 212 => to_unsigned(3670, 12), 213 => to_unsigned(2780, 12), 214 => to_unsigned(2653, 12), 215 => to_unsigned(521, 12), 216 => to_unsigned(336, 12), 217 => to_unsigned(2958, 12), 218 => to_unsigned(475, 12), 219 => to_unsigned(2300, 12), 220 => to_unsigned(767, 12), 221 => to_unsigned(1207, 12), 222 => to_unsigned(2622, 12), 223 => to_unsigned(1740, 12), 224 => to_unsigned(706, 12), 225 => to_unsigned(976, 12), 226 => to_unsigned(1001, 12), 227 => to_unsigned(2472, 12), 228 => to_unsigned(3879, 12), 229 => to_unsigned(3713, 12), 230 => to_unsigned(2351, 12), 231 => to_unsigned(1769, 12), 232 => to_unsigned(2906, 12), 233 => to_unsigned(4011, 12), 234 => to_unsigned(1195, 12), 235 => to_unsigned(3096, 12), 236 => to_unsigned(925, 12), 237 => to_unsigned(2193, 12), 238 => to_unsigned(1663, 12), 239 => to_unsigned(1708, 12), 240 => to_unsigned(484, 12), 241 => to_unsigned(1255, 12), 242 => to_unsigned(3762, 12), 243 => to_unsigned(2853, 12), 244 => to_unsigned(1491, 12), 245 => to_unsigned(3003, 12), 246 => to_unsigned(2025, 12), 247 => to_unsigned(2486, 12), 248 => to_unsigned(2169, 12), 249 => to_unsigned(3517, 12), 250 => to_unsigned(1934, 12), 251 => to_unsigned(1062, 12), 252 => to_unsigned(2874, 12), 253 => to_unsigned(1645, 12), 254 => to_unsigned(1417, 12), 255 => to_unsigned(1496, 12), 256 => to_unsigned(1547, 12), 257 => to_unsigned(272, 12), 258 => to_unsigned(751, 12), 259 => to_unsigned(3669, 12), 260 => to_unsigned(1150, 12), 261 => to_unsigned(2987, 12), 262 => to_unsigned(1805, 12), 263 => to_unsigned(1430, 12), 264 => to_unsigned(2037, 12), 265 => to_unsigned(536, 12), 266 => to_unsigned(907, 12), 267 => to_unsigned(339, 12), 268 => to_unsigned(1373, 12), 269 => to_unsigned(2223, 12), 270 => to_unsigned(3676, 12), 271 => to_unsigned(2428, 12), 272 => to_unsigned(344, 12), 273 => to_unsigned(1588, 12), 274 => to_unsigned(182, 12), 275 => to_unsigned(98, 12), 276 => to_unsigned(74, 12), 277 => to_unsigned(2462, 12), 278 => to_unsigned(3051, 12), 279 => to_unsigned(753, 12), 280 => to_unsigned(1458, 12), 281 => to_unsigned(323, 12), 282 => to_unsigned(2217, 12), 283 => to_unsigned(2291, 12), 284 => to_unsigned(3401, 12), 285 => to_unsigned(306, 12), 286 => to_unsigned(1894, 12), 287 => to_unsigned(3575, 12), 288 => to_unsigned(2614, 12), 289 => to_unsigned(2651, 12), 290 => to_unsigned(2942, 12), 291 => to_unsigned(3076, 12), 292 => to_unsigned(129, 12), 293 => to_unsigned(3038, 12), 294 => to_unsigned(3836, 12), 295 => to_unsigned(1137, 12), 296 => to_unsigned(3931, 12), 297 => to_unsigned(3863, 12), 298 => to_unsigned(729, 12), 299 => to_unsigned(3730, 12), 300 => to_unsigned(922, 12), 301 => to_unsigned(340, 12), 302 => to_unsigned(1349, 12), 303 => to_unsigned(4024, 12), 304 => to_unsigned(2316, 12), 305 => to_unsigned(3308, 12), 306 => to_unsigned(3087, 12), 307 => to_unsigned(3854, 12), 308 => to_unsigned(2462, 12), 309 => to_unsigned(1992, 12), 310 => to_unsigned(2355, 12), 311 => to_unsigned(737, 12), 312 => to_unsigned(1434, 12), 313 => to_unsigned(2158, 12), 314 => to_unsigned(3276, 12), 315 => to_unsigned(3443, 12), 316 => to_unsigned(2607, 12), 317 => to_unsigned(2114, 12), 318 => to_unsigned(1136, 12), 319 => to_unsigned(3987, 12), 320 => to_unsigned(132, 12), 321 => to_unsigned(1723, 12), 322 => to_unsigned(654, 12), 323 => to_unsigned(1722, 12), 324 => to_unsigned(1315, 12), 325 => to_unsigned(263, 12), 326 => to_unsigned(3469, 12), 327 => to_unsigned(1472, 12), 328 => to_unsigned(3367, 12), 329 => to_unsigned(1927, 12), 330 => to_unsigned(1273, 12), 331 => to_unsigned(1507, 12), 332 => to_unsigned(2367, 12), 333 => to_unsigned(1410, 12), 334 => to_unsigned(3815, 12), 335 => to_unsigned(138, 12), 336 => to_unsigned(1878, 12), 337 => to_unsigned(1949, 12), 338 => to_unsigned(1454, 12), 339 => to_unsigned(136, 12), 340 => to_unsigned(3747, 12), 341 => to_unsigned(824, 12), 342 => to_unsigned(640, 12), 343 => to_unsigned(95, 12), 344 => to_unsigned(3270, 12), 345 => to_unsigned(2917, 12), 346 => to_unsigned(16, 12), 347 => to_unsigned(3785, 12), 348 => to_unsigned(3263, 12), 349 => to_unsigned(862, 12), 350 => to_unsigned(21, 12), 351 => to_unsigned(2494, 12), 352 => to_unsigned(3420, 12), 353 => to_unsigned(3105, 12), 354 => to_unsigned(4093, 12), 355 => to_unsigned(3335, 12), 356 => to_unsigned(398, 12), 357 => to_unsigned(3056, 12), 358 => to_unsigned(1718, 12), 359 => to_unsigned(3215, 12), 360 => to_unsigned(3482, 12), 361 => to_unsigned(523, 12), 362 => to_unsigned(3790, 12), 363 => to_unsigned(1577, 12), 364 => to_unsigned(312, 12), 365 => to_unsigned(3792, 12), 366 => to_unsigned(2026, 12), 367 => to_unsigned(3352, 12), 368 => to_unsigned(2434, 12), 369 => to_unsigned(4031, 12), 370 => to_unsigned(3935, 12), 371 => to_unsigned(4082, 12), 372 => to_unsigned(3908, 12), 373 => to_unsigned(43, 12), 374 => to_unsigned(3187, 12), 375 => to_unsigned(649, 12), 376 => to_unsigned(3929, 12), 377 => to_unsigned(1211, 12), 378 => to_unsigned(2337, 12), 379 => to_unsigned(3355, 12), 380 => to_unsigned(3850, 12), 381 => to_unsigned(370, 12), 382 => to_unsigned(1511, 12), 383 => to_unsigned(222, 12), 384 => to_unsigned(1006, 12), 385 => to_unsigned(829, 12), 386 => to_unsigned(2202, 12), 387 => to_unsigned(800, 12), 388 => to_unsigned(2129, 12), 389 => to_unsigned(3741, 12), 390 => to_unsigned(2796, 12), 391 => to_unsigned(3549, 12), 392 => to_unsigned(440, 12), 393 => to_unsigned(1318, 12), 394 => to_unsigned(3304, 12), 395 => to_unsigned(901, 12), 396 => to_unsigned(289, 12), 397 => to_unsigned(288, 12), 398 => to_unsigned(1738, 12), 399 => to_unsigned(114, 12), 400 => to_unsigned(3497, 12), 401 => to_unsigned(1662, 12), 402 => to_unsigned(3626, 12), 403 => to_unsigned(3707, 12), 404 => to_unsigned(2738, 12), 405 => to_unsigned(1526, 12), 406 => to_unsigned(3662, 12), 407 => to_unsigned(2331, 12), 408 => to_unsigned(2352, 12), 409 => to_unsigned(779, 12), 410 => to_unsigned(2611, 12), 411 => to_unsigned(1479, 12), 412 => to_unsigned(1036, 12), 413 => to_unsigned(3168, 12), 414 => to_unsigned(566, 12), 415 => to_unsigned(2231, 12), 416 => to_unsigned(11, 12), 417 => to_unsigned(443, 12), 418 => to_unsigned(2138, 12), 419 => to_unsigned(883, 12), 420 => to_unsigned(2053, 12), 421 => to_unsigned(4093, 12), 422 => to_unsigned(170, 12), 423 => to_unsigned(1527, 12), 424 => to_unsigned(1839, 12), 425 => to_unsigned(2312, 12), 426 => to_unsigned(533, 12), 427 => to_unsigned(2758, 12), 428 => to_unsigned(2776, 12), 429 => to_unsigned(2792, 12), 430 => to_unsigned(1253, 12), 431 => to_unsigned(3613, 12), 432 => to_unsigned(781, 12), 433 => to_unsigned(547, 12), 434 => to_unsigned(3077, 12), 435 => to_unsigned(1012, 12), 436 => to_unsigned(2165, 12), 437 => to_unsigned(3277, 12), 438 => to_unsigned(3749, 12), 439 => to_unsigned(3614, 12), 440 => to_unsigned(2656, 12), 441 => to_unsigned(1474, 12), 442 => to_unsigned(2100, 12), 443 => to_unsigned(77, 12), 444 => to_unsigned(118, 12), 445 => to_unsigned(3003, 12), 446 => to_unsigned(381, 12), 447 => to_unsigned(4062, 12), 448 => to_unsigned(1920, 12), 449 => to_unsigned(1673, 12), 450 => to_unsigned(1426, 12), 451 => to_unsigned(3503, 12), 452 => to_unsigned(1424, 12), 453 => to_unsigned(2091, 12), 454 => to_unsigned(1577, 12), 455 => to_unsigned(1231, 12), 456 => to_unsigned(3605, 12), 457 => to_unsigned(2069, 12), 458 => to_unsigned(1270, 12), 459 => to_unsigned(2667, 12), 460 => to_unsigned(3739, 12), 461 => to_unsigned(3006, 12), 462 => to_unsigned(2542, 12), 463 => to_unsigned(3225, 12), 464 => to_unsigned(1796, 12), 465 => to_unsigned(1752, 12), 466 => to_unsigned(3720, 12), 467 => to_unsigned(2357, 12), 468 => to_unsigned(215, 12), 469 => to_unsigned(2395, 12), 470 => to_unsigned(3944, 12), 471 => to_unsigned(3173, 12), 472 => to_unsigned(156, 12), 473 => to_unsigned(3562, 12), 474 => to_unsigned(2927, 12), 475 => to_unsigned(1822, 12), 476 => to_unsigned(737, 12), 477 => to_unsigned(973, 12), 478 => to_unsigned(307, 12), 479 => to_unsigned(1256, 12), 480 => to_unsigned(2006, 12), 481 => to_unsigned(1489, 12), 482 => to_unsigned(2986, 12), 483 => to_unsigned(1603, 12), 484 => to_unsigned(1575, 12), 485 => to_unsigned(3796, 12), 486 => to_unsigned(1794, 12), 487 => to_unsigned(799, 12), 488 => to_unsigned(3791, 12), 489 => to_unsigned(2558, 12), 490 => to_unsigned(777, 12), 491 => to_unsigned(1362, 12), 492 => to_unsigned(1508, 12), 493 => to_unsigned(599, 12), 494 => to_unsigned(337, 12), 495 => to_unsigned(2131, 12), 496 => to_unsigned(2627, 12), 497 => to_unsigned(3045, 12), 498 => to_unsigned(1417, 12), 499 => to_unsigned(1219, 12), 500 => to_unsigned(3574, 12), 501 => to_unsigned(2502, 12), 502 => to_unsigned(3152, 12), 503 => to_unsigned(1384, 12), 504 => to_unsigned(3307, 12), 505 => to_unsigned(3031, 12), 506 => to_unsigned(4062, 12), 507 => to_unsigned(3172, 12), 508 => to_unsigned(2522, 12), 509 => to_unsigned(1049, 12), 510 => to_unsigned(739, 12), 511 => to_unsigned(44, 12), 512 => to_unsigned(1249, 12), 513 => to_unsigned(560, 12), 514 => to_unsigned(4064, 12), 515 => to_unsigned(3140, 12), 516 => to_unsigned(1377, 12), 517 => to_unsigned(3086, 12), 518 => to_unsigned(216, 12), 519 => to_unsigned(1009, 12), 520 => to_unsigned(135, 12), 521 => to_unsigned(45, 12), 522 => to_unsigned(242, 12), 523 => to_unsigned(740, 12), 524 => to_unsigned(3841, 12), 525 => to_unsigned(2659, 12), 526 => to_unsigned(80, 12), 527 => to_unsigned(3042, 12), 528 => to_unsigned(2416, 12), 529 => to_unsigned(3960, 12), 530 => to_unsigned(262, 12), 531 => to_unsigned(968, 12), 532 => to_unsigned(3181, 12), 533 => to_unsigned(502, 12), 534 => to_unsigned(1694, 12), 535 => to_unsigned(2185, 12), 536 => to_unsigned(265, 12), 537 => to_unsigned(1261, 12), 538 => to_unsigned(3470, 12), 539 => to_unsigned(240, 12), 540 => to_unsigned(3142, 12), 541 => to_unsigned(1034, 12), 542 => to_unsigned(3979, 12), 543 => to_unsigned(3766, 12), 544 => to_unsigned(1890, 12), 545 => to_unsigned(1772, 12), 546 => to_unsigned(3525, 12), 547 => to_unsigned(879, 12), 548 => to_unsigned(1432, 12), 549 => to_unsigned(470, 12), 550 => to_unsigned(1306, 12), 551 => to_unsigned(114, 12), 552 => to_unsigned(3520, 12), 553 => to_unsigned(2234, 12), 554 => to_unsigned(2339, 12), 555 => to_unsigned(3691, 12), 556 => to_unsigned(3842, 12), 557 => to_unsigned(2099, 12), 558 => to_unsigned(1089, 12), 559 => to_unsigned(2874, 12), 560 => to_unsigned(135, 12), 561 => to_unsigned(338, 12), 562 => to_unsigned(3820, 12), 563 => to_unsigned(613, 12), 564 => to_unsigned(3440, 12), 565 => to_unsigned(3088, 12), 566 => to_unsigned(1752, 12), 567 => to_unsigned(1077, 12), 568 => to_unsigned(2260, 12), 569 => to_unsigned(3812, 12), 570 => to_unsigned(3713, 12), 571 => to_unsigned(687, 12), 572 => to_unsigned(522, 12), 573 => to_unsigned(517, 12), 574 => to_unsigned(2397, 12), 575 => to_unsigned(3214, 12), 576 => to_unsigned(3217, 12), 577 => to_unsigned(3166, 12), 578 => to_unsigned(3087, 12), 579 => to_unsigned(766, 12), 580 => to_unsigned(2478, 12), 581 => to_unsigned(175, 12), 582 => to_unsigned(3731, 12), 583 => to_unsigned(767, 12), 584 => to_unsigned(3637, 12), 585 => to_unsigned(2998, 12), 586 => to_unsigned(4008, 12), 587 => to_unsigned(381, 12), 588 => to_unsigned(430, 12), 589 => to_unsigned(2712, 12), 590 => to_unsigned(49, 12), 591 => to_unsigned(464, 12), 592 => to_unsigned(2584, 12), 593 => to_unsigned(1740, 12), 594 => to_unsigned(993, 12), 595 => to_unsigned(243, 12), 596 => to_unsigned(1468, 12), 597 => to_unsigned(1021, 12), 598 => to_unsigned(3524, 12), 599 => to_unsigned(2196, 12), 600 => to_unsigned(3381, 12), 601 => to_unsigned(1621, 12), 602 => to_unsigned(3513, 12), 603 => to_unsigned(69, 12), 604 => to_unsigned(4007, 12), 605 => to_unsigned(1887, 12), 606 => to_unsigned(128, 12), 607 => to_unsigned(652, 12), 608 => to_unsigned(3173, 12), 609 => to_unsigned(982, 12), 610 => to_unsigned(3246, 12), 611 => to_unsigned(985, 12), 612 => to_unsigned(3159, 12), 613 => to_unsigned(748, 12), 614 => to_unsigned(2775, 12), 615 => to_unsigned(732, 12), 616 => to_unsigned(1511, 12), 617 => to_unsigned(28, 12), 618 => to_unsigned(4007, 12), 619 => to_unsigned(1416, 12), 620 => to_unsigned(1381, 12), 621 => to_unsigned(740, 12), 622 => to_unsigned(785, 12), 623 => to_unsigned(207, 12), 624 => to_unsigned(1461, 12), 625 => to_unsigned(1364, 12), 626 => to_unsigned(1345, 12), 627 => to_unsigned(1268, 12), 628 => to_unsigned(3087, 12), 629 => to_unsigned(3314, 12), 630 => to_unsigned(3685, 12), 631 => to_unsigned(2364, 12), 632 => to_unsigned(1658, 12), 633 => to_unsigned(1800, 12), 634 => to_unsigned(3772, 12), 635 => to_unsigned(1601, 12), 636 => to_unsigned(1206, 12), 637 => to_unsigned(3536, 12), 638 => to_unsigned(3279, 12), 639 => to_unsigned(1449, 12), 640 => to_unsigned(641, 12), 641 => to_unsigned(2280, 12), 642 => to_unsigned(639, 12), 643 => to_unsigned(3007, 12), 644 => to_unsigned(2686, 12), 645 => to_unsigned(142, 12), 646 => to_unsigned(2324, 12), 647 => to_unsigned(1795, 12), 648 => to_unsigned(156, 12), 649 => to_unsigned(3424, 12), 650 => to_unsigned(2744, 12), 651 => to_unsigned(3935, 12), 652 => to_unsigned(161, 12), 653 => to_unsigned(1438, 12), 654 => to_unsigned(347, 12), 655 => to_unsigned(1047, 12), 656 => to_unsigned(2609, 12), 657 => to_unsigned(701, 12), 658 => to_unsigned(2302, 12), 659 => to_unsigned(3525, 12), 660 => to_unsigned(2923, 12), 661 => to_unsigned(3189, 12), 662 => to_unsigned(671, 12), 663 => to_unsigned(1027, 12), 664 => to_unsigned(38, 12), 665 => to_unsigned(3895, 12), 666 => to_unsigned(1138, 12), 667 => to_unsigned(3686, 12), 668 => to_unsigned(1073, 12), 669 => to_unsigned(2126, 12), 670 => to_unsigned(1282, 12), 671 => to_unsigned(2147, 12), 672 => to_unsigned(1261, 12), 673 => to_unsigned(2007, 12), 674 => to_unsigned(12, 12), 675 => to_unsigned(841, 12), 676 => to_unsigned(1334, 12), 677 => to_unsigned(607, 12), 678 => to_unsigned(1750, 12), 679 => to_unsigned(512, 12), 680 => to_unsigned(2849, 12), 681 => to_unsigned(1379, 12), 682 => to_unsigned(2018, 12), 683 => to_unsigned(35, 12), 684 => to_unsigned(4032, 12), 685 => to_unsigned(2220, 12), 686 => to_unsigned(2397, 12), 687 => to_unsigned(3116, 12), 688 => to_unsigned(638, 12), 689 => to_unsigned(3856, 12), 690 => to_unsigned(2498, 12), 691 => to_unsigned(2435, 12), 692 => to_unsigned(1953, 12), 693 => to_unsigned(47, 12), 694 => to_unsigned(1045, 12), 695 => to_unsigned(1506, 12), 696 => to_unsigned(157, 12), 697 => to_unsigned(1275, 12), 698 => to_unsigned(3257, 12), 699 => to_unsigned(3953, 12), 700 => to_unsigned(686, 12), 701 => to_unsigned(2512, 12), 702 => to_unsigned(769, 12), 703 => to_unsigned(2077, 12), 704 => to_unsigned(795, 12), 705 => to_unsigned(3218, 12), 706 => to_unsigned(1575, 12), 707 => to_unsigned(2294, 12), 708 => to_unsigned(3244, 12), 709 => to_unsigned(1876, 12), 710 => to_unsigned(2826, 12), 711 => to_unsigned(2368, 12), 712 => to_unsigned(2490, 12), 713 => to_unsigned(417, 12), 714 => to_unsigned(3884, 12), 715 => to_unsigned(589, 12), 716 => to_unsigned(3731, 12), 717 => to_unsigned(2684, 12), 718 => to_unsigned(1614, 12), 719 => to_unsigned(3502, 12), 720 => to_unsigned(849, 12), 721 => to_unsigned(981, 12), 722 => to_unsigned(3661, 12), 723 => to_unsigned(924, 12), 724 => to_unsigned(3342, 12), 725 => to_unsigned(3010, 12), 726 => to_unsigned(1651, 12), 727 => to_unsigned(1583, 12), 728 => to_unsigned(1822, 12), 729 => to_unsigned(946, 12), 730 => to_unsigned(1854, 12), 731 => to_unsigned(247, 12), 732 => to_unsigned(1407, 12), 733 => to_unsigned(3105, 12), 734 => to_unsigned(714, 12), 735 => to_unsigned(3199, 12), 736 => to_unsigned(762, 12), 737 => to_unsigned(616, 12), 738 => to_unsigned(229, 12), 739 => to_unsigned(1241, 12), 740 => to_unsigned(3119, 12), 741 => to_unsigned(1644, 12), 742 => to_unsigned(2027, 12), 743 => to_unsigned(937, 12), 744 => to_unsigned(631, 12), 745 => to_unsigned(2593, 12), 746 => to_unsigned(3584, 12), 747 => to_unsigned(3333, 12), 748 => to_unsigned(618, 12), 749 => to_unsigned(1598, 12), 750 => to_unsigned(3243, 12), 751 => to_unsigned(794, 12), 752 => to_unsigned(3903, 12), 753 => to_unsigned(553, 12), 754 => to_unsigned(2843, 12), 755 => to_unsigned(526, 12), 756 => to_unsigned(1519, 12), 757 => to_unsigned(1648, 12), 758 => to_unsigned(258, 12), 759 => to_unsigned(1043, 12), 760 => to_unsigned(1164, 12), 761 => to_unsigned(880, 12), 762 => to_unsigned(287, 12), 763 => to_unsigned(1713, 12), 764 => to_unsigned(550, 12), 765 => to_unsigned(478, 12), 766 => to_unsigned(1590, 12), 767 => to_unsigned(1771, 12), 768 => to_unsigned(2817, 12), 769 => to_unsigned(634, 12), 770 => to_unsigned(801, 12), 771 => to_unsigned(3647, 12), 772 => to_unsigned(3559, 12), 773 => to_unsigned(2481, 12), 774 => to_unsigned(3920, 12), 775 => to_unsigned(4090, 12), 776 => to_unsigned(3884, 12), 777 => to_unsigned(2162, 12), 778 => to_unsigned(2060, 12), 779 => to_unsigned(3227, 12), 780 => to_unsigned(3158, 12), 781 => to_unsigned(1134, 12), 782 => to_unsigned(3822, 12), 783 => to_unsigned(716, 12), 784 => to_unsigned(1637, 12), 785 => to_unsigned(2163, 12), 786 => to_unsigned(1165, 12), 787 => to_unsigned(2678, 12), 788 => to_unsigned(839, 12), 789 => to_unsigned(931, 12), 790 => to_unsigned(2796, 12), 791 => to_unsigned(3006, 12), 792 => to_unsigned(1085, 12), 793 => to_unsigned(2262, 12), 794 => to_unsigned(235, 12), 795 => to_unsigned(468, 12), 796 => to_unsigned(1824, 12), 797 => to_unsigned(2877, 12), 798 => to_unsigned(1022, 12), 799 => to_unsigned(1267, 12), 800 => to_unsigned(3762, 12), 801 => to_unsigned(415, 12), 802 => to_unsigned(181, 12), 803 => to_unsigned(1362, 12), 804 => to_unsigned(2279, 12), 805 => to_unsigned(1467, 12), 806 => to_unsigned(563, 12), 807 => to_unsigned(906, 12), 808 => to_unsigned(4042, 12), 809 => to_unsigned(1254, 12), 810 => to_unsigned(92, 12), 811 => to_unsigned(2362, 12), 812 => to_unsigned(4001, 12), 813 => to_unsigned(3679, 12), 814 => to_unsigned(3644, 12), 815 => to_unsigned(2332, 12), 816 => to_unsigned(2640, 12), 817 => to_unsigned(2409, 12), 818 => to_unsigned(3836, 12), 819 => to_unsigned(2673, 12), 820 => to_unsigned(3345, 12), 821 => to_unsigned(1360, 12), 822 => to_unsigned(2266, 12), 823 => to_unsigned(1869, 12), 824 => to_unsigned(1987, 12), 825 => to_unsigned(1478, 12), 826 => to_unsigned(145, 12), 827 => to_unsigned(2312, 12), 828 => to_unsigned(1756, 12), 829 => to_unsigned(2519, 12), 830 => to_unsigned(551, 12), 831 => to_unsigned(3354, 12), 832 => to_unsigned(2139, 12), 833 => to_unsigned(1186, 12), 834 => to_unsigned(287, 12), 835 => to_unsigned(2238, 12), 836 => to_unsigned(1374, 12), 837 => to_unsigned(2473, 12), 838 => to_unsigned(223, 12), 839 => to_unsigned(2390, 12), 840 => to_unsigned(1725, 12), 841 => to_unsigned(3083, 12), 842 => to_unsigned(356, 12), 843 => to_unsigned(1107, 12), 844 => to_unsigned(999, 12), 845 => to_unsigned(563, 12), 846 => to_unsigned(2846, 12), 847 => to_unsigned(23, 12), 848 => to_unsigned(1667, 12), 849 => to_unsigned(59, 12), 850 => to_unsigned(1535, 12), 851 => to_unsigned(1363, 12), 852 => to_unsigned(885, 12), 853 => to_unsigned(609, 12), 854 => to_unsigned(827, 12), 855 => to_unsigned(2053, 12), 856 => to_unsigned(171, 12), 857 => to_unsigned(26, 12), 858 => to_unsigned(2035, 12), 859 => to_unsigned(1394, 12), 860 => to_unsigned(3117, 12), 861 => to_unsigned(2709, 12), 862 => to_unsigned(186, 12), 863 => to_unsigned(1263, 12), 864 => to_unsigned(2625, 12), 865 => to_unsigned(1987, 12), 866 => to_unsigned(2603, 12), 867 => to_unsigned(4049, 12), 868 => to_unsigned(2509, 12), 869 => to_unsigned(432, 12), 870 => to_unsigned(1506, 12), 871 => to_unsigned(3398, 12), 872 => to_unsigned(4048, 12), 873 => to_unsigned(2638, 12), 874 => to_unsigned(2092, 12), 875 => to_unsigned(3900, 12), 876 => to_unsigned(479, 12), 877 => to_unsigned(3109, 12), 878 => to_unsigned(601, 12), 879 => to_unsigned(734, 12), 880 => to_unsigned(3297, 12), 881 => to_unsigned(2366, 12), 882 => to_unsigned(658, 12), 883 => to_unsigned(2624, 12), 884 => to_unsigned(939, 12), 885 => to_unsigned(3158, 12), 886 => to_unsigned(3699, 12), 887 => to_unsigned(3559, 12), 888 => to_unsigned(4004, 12), 889 => to_unsigned(3394, 12), 890 => to_unsigned(1489, 12), 891 => to_unsigned(3506, 12), 892 => to_unsigned(2763, 12), 893 => to_unsigned(3329, 12), 894 => to_unsigned(3722, 12), 895 => to_unsigned(328, 12), 896 => to_unsigned(175, 12), 897 => to_unsigned(481, 12), 898 => to_unsigned(51, 12), 899 => to_unsigned(2339, 12), 900 => to_unsigned(865, 12), 901 => to_unsigned(2509, 12), 902 => to_unsigned(71, 12), 903 => to_unsigned(1266, 12), 904 => to_unsigned(2474, 12), 905 => to_unsigned(1582, 12), 906 => to_unsigned(1643, 12), 907 => to_unsigned(2668, 12), 908 => to_unsigned(1695, 12), 909 => to_unsigned(2474, 12), 910 => to_unsigned(2174, 12), 911 => to_unsigned(2616, 12), 912 => to_unsigned(468, 12), 913 => to_unsigned(3033, 12), 914 => to_unsigned(3188, 12), 915 => to_unsigned(1760, 12), 916 => to_unsigned(1024, 12), 917 => to_unsigned(637, 12), 918 => to_unsigned(1217, 12), 919 => to_unsigned(430, 12), 920 => to_unsigned(892, 12), 921 => to_unsigned(2499, 12), 922 => to_unsigned(578, 12), 923 => to_unsigned(3275, 12), 924 => to_unsigned(942, 12), 925 => to_unsigned(1784, 12), 926 => to_unsigned(3684, 12), 927 => to_unsigned(1369, 12), 928 => to_unsigned(3608, 12), 929 => to_unsigned(2366, 12), 930 => to_unsigned(3910, 12), 931 => to_unsigned(746, 12), 932 => to_unsigned(885, 12), 933 => to_unsigned(3326, 12), 934 => to_unsigned(1715, 12), 935 => to_unsigned(1252, 12), 936 => to_unsigned(1784, 12), 937 => to_unsigned(1373, 12), 938 => to_unsigned(3542, 12), 939 => to_unsigned(3438, 12), 940 => to_unsigned(4006, 12), 941 => to_unsigned(2404, 12), 942 => to_unsigned(1421, 12), 943 => to_unsigned(2600, 12), 944 => to_unsigned(3675, 12), 945 => to_unsigned(237, 12), 946 => to_unsigned(2603, 12), 947 => to_unsigned(529, 12), 948 => to_unsigned(310, 12), 949 => to_unsigned(237, 12), 950 => to_unsigned(712, 12), 951 => to_unsigned(2703, 12), 952 => to_unsigned(1864, 12), 953 => to_unsigned(3650, 12), 954 => to_unsigned(3224, 12), 955 => to_unsigned(1998, 12), 956 => to_unsigned(975, 12), 957 => to_unsigned(810, 12), 958 => to_unsigned(3443, 12), 959 => to_unsigned(3278, 12), 960 => to_unsigned(11, 12), 961 => to_unsigned(3632, 12), 962 => to_unsigned(3704, 12), 963 => to_unsigned(3518, 12), 964 => to_unsigned(238, 12), 965 => to_unsigned(2474, 12), 966 => to_unsigned(2141, 12), 967 => to_unsigned(2651, 12), 968 => to_unsigned(3036, 12), 969 => to_unsigned(3801, 12), 970 => to_unsigned(2285, 12), 971 => to_unsigned(1540, 12), 972 => to_unsigned(3881, 12), 973 => to_unsigned(3920, 12), 974 => to_unsigned(3376, 12), 975 => to_unsigned(2165, 12), 976 => to_unsigned(3402, 12), 977 => to_unsigned(2428, 12), 978 => to_unsigned(76, 12), 979 => to_unsigned(2278, 12), 980 => to_unsigned(3315, 12), 981 => to_unsigned(332, 12), 982 => to_unsigned(3640, 12), 983 => to_unsigned(392, 12), 984 => to_unsigned(3416, 12), 985 => to_unsigned(951, 12), 986 => to_unsigned(442, 12), 987 => to_unsigned(1629, 12), 988 => to_unsigned(2667, 12), 989 => to_unsigned(2538, 12), 990 => to_unsigned(3628, 12), 991 => to_unsigned(1908, 12), 992 => to_unsigned(614, 12), 993 => to_unsigned(3644, 12), 994 => to_unsigned(702, 12), 995 => to_unsigned(1842, 12), 996 => to_unsigned(2902, 12), 997 => to_unsigned(348, 12), 998 => to_unsigned(3675, 12), 999 => to_unsigned(819, 12), 1000 => to_unsigned(3664, 12), 1001 => to_unsigned(2817, 12), 1002 => to_unsigned(1304, 12), 1003 => to_unsigned(2101, 12), 1004 => to_unsigned(2021, 12), 1005 => to_unsigned(536, 12), 1006 => to_unsigned(963, 12), 1007 => to_unsigned(2103, 12), 1008 => to_unsigned(3942, 12), 1009 => to_unsigned(2987, 12), 1010 => to_unsigned(991, 12), 1011 => to_unsigned(2207, 12), 1012 => to_unsigned(2214, 12), 1013 => to_unsigned(850, 12), 1014 => to_unsigned(2509, 12), 1015 => to_unsigned(2398, 12), 1016 => to_unsigned(2756, 12), 1017 => to_unsigned(777, 12), 1018 => to_unsigned(2141, 12), 1019 => to_unsigned(2842, 12), 1020 => to_unsigned(3058, 12), 1021 => to_unsigned(3555, 12), 1022 => to_unsigned(3363, 12), 1023 => to_unsigned(671, 12), 1024 => to_unsigned(3788, 12), 1025 => to_unsigned(1297, 12), 1026 => to_unsigned(3016, 12), 1027 => to_unsigned(2780, 12), 1028 => to_unsigned(3599, 12), 1029 => to_unsigned(1884, 12), 1030 => to_unsigned(3112, 12), 1031 => to_unsigned(893, 12), 1032 => to_unsigned(180, 12), 1033 => to_unsigned(4095, 12), 1034 => to_unsigned(994, 12), 1035 => to_unsigned(447, 12), 1036 => to_unsigned(1684, 12), 1037 => to_unsigned(210, 12), 1038 => to_unsigned(1967, 12), 1039 => to_unsigned(1152, 12), 1040 => to_unsigned(2159, 12), 1041 => to_unsigned(4051, 12), 1042 => to_unsigned(1164, 12), 1043 => to_unsigned(917, 12), 1044 => to_unsigned(2069, 12), 1045 => to_unsigned(1586, 12), 1046 => to_unsigned(3898, 12), 1047 => to_unsigned(2375, 12), 1048 => to_unsigned(890, 12), 1049 => to_unsigned(370, 12), 1050 => to_unsigned(1686, 12), 1051 => to_unsigned(2569, 12), 1052 => to_unsigned(192, 12), 1053 => to_unsigned(1745, 12), 1054 => to_unsigned(2437, 12), 1055 => to_unsigned(588, 12), 1056 => to_unsigned(3376, 12), 1057 => to_unsigned(1281, 12), 1058 => to_unsigned(701, 12), 1059 => to_unsigned(903, 12), 1060 => to_unsigned(2019, 12), 1061 => to_unsigned(1116, 12), 1062 => to_unsigned(2873, 12), 1063 => to_unsigned(2896, 12), 1064 => to_unsigned(157, 12), 1065 => to_unsigned(2658, 12), 1066 => to_unsigned(193, 12), 1067 => to_unsigned(3876, 12), 1068 => to_unsigned(1296, 12), 1069 => to_unsigned(1964, 12), 1070 => to_unsigned(220, 12), 1071 => to_unsigned(2946, 12), 1072 => to_unsigned(1152, 12), 1073 => to_unsigned(2195, 12), 1074 => to_unsigned(746, 12), 1075 => to_unsigned(1303, 12), 1076 => to_unsigned(3689, 12), 1077 => to_unsigned(3218, 12), 1078 => to_unsigned(388, 12), 1079 => to_unsigned(771, 12), 1080 => to_unsigned(900, 12), 1081 => to_unsigned(2157, 12), 1082 => to_unsigned(2301, 12), 1083 => to_unsigned(1370, 12), 1084 => to_unsigned(2279, 12), 1085 => to_unsigned(2383, 12), 1086 => to_unsigned(3974, 12), 1087 => to_unsigned(3828, 12), 1088 => to_unsigned(3199, 12), 1089 => to_unsigned(1626, 12), 1090 => to_unsigned(2561, 12), 1091 => to_unsigned(1780, 12), 1092 => to_unsigned(4028, 12), 1093 => to_unsigned(70, 12), 1094 => to_unsigned(800, 12), 1095 => to_unsigned(173, 12), 1096 => to_unsigned(2645, 12), 1097 => to_unsigned(2757, 12), 1098 => to_unsigned(2061, 12), 1099 => to_unsigned(999, 12), 1100 => to_unsigned(3198, 12), 1101 => to_unsigned(3226, 12), 1102 => to_unsigned(2074, 12), 1103 => to_unsigned(2838, 12), 1104 => to_unsigned(2637, 12), 1105 => to_unsigned(3124, 12), 1106 => to_unsigned(3432, 12), 1107 => to_unsigned(1908, 12), 1108 => to_unsigned(1814, 12), 1109 => to_unsigned(1680, 12), 1110 => to_unsigned(24, 12), 1111 => to_unsigned(3820, 12), 1112 => to_unsigned(2572, 12), 1113 => to_unsigned(77, 12), 1114 => to_unsigned(1963, 12), 1115 => to_unsigned(868, 12), 1116 => to_unsigned(2264, 12), 1117 => to_unsigned(1191, 12), 1118 => to_unsigned(1021, 12), 1119 => to_unsigned(1572, 12), 1120 => to_unsigned(2426, 12), 1121 => to_unsigned(3946, 12), 1122 => to_unsigned(2285, 12), 1123 => to_unsigned(2629, 12), 1124 => to_unsigned(2244, 12), 1125 => to_unsigned(2408, 12), 1126 => to_unsigned(2679, 12), 1127 => to_unsigned(2322, 12), 1128 => to_unsigned(1571, 12), 1129 => to_unsigned(1, 12), 1130 => to_unsigned(2298, 12), 1131 => to_unsigned(674, 12), 1132 => to_unsigned(708, 12), 1133 => to_unsigned(1260, 12), 1134 => to_unsigned(2264, 12), 1135 => to_unsigned(3651, 12), 1136 => to_unsigned(51, 12), 1137 => to_unsigned(3824, 12), 1138 => to_unsigned(729, 12), 1139 => to_unsigned(764, 12), 1140 => to_unsigned(1515, 12), 1141 => to_unsigned(2761, 12), 1142 => to_unsigned(3605, 12), 1143 => to_unsigned(3319, 12), 1144 => to_unsigned(3473, 12), 1145 => to_unsigned(1551, 12), 1146 => to_unsigned(2847, 12), 1147 => to_unsigned(495, 12), 1148 => to_unsigned(790, 12), 1149 => to_unsigned(3221, 12), 1150 => to_unsigned(576, 12), 1151 => to_unsigned(2925, 12), 1152 => to_unsigned(3817, 12), 1153 => to_unsigned(3071, 12), 1154 => to_unsigned(88, 12), 1155 => to_unsigned(1171, 12), 1156 => to_unsigned(1763, 12), 1157 => to_unsigned(2916, 12), 1158 => to_unsigned(385, 12), 1159 => to_unsigned(3630, 12), 1160 => to_unsigned(1846, 12), 1161 => to_unsigned(2171, 12), 1162 => to_unsigned(3371, 12), 1163 => to_unsigned(925, 12), 1164 => to_unsigned(3769, 12), 1165 => to_unsigned(2326, 12), 1166 => to_unsigned(3484, 12), 1167 => to_unsigned(596, 12), 1168 => to_unsigned(3411, 12), 1169 => to_unsigned(1329, 12), 1170 => to_unsigned(1586, 12), 1171 => to_unsigned(1033, 12), 1172 => to_unsigned(3043, 12), 1173 => to_unsigned(3874, 12), 1174 => to_unsigned(82, 12), 1175 => to_unsigned(105, 12), 1176 => to_unsigned(4004, 12), 1177 => to_unsigned(1780, 12), 1178 => to_unsigned(2729, 12), 1179 => to_unsigned(1099, 12), 1180 => to_unsigned(949, 12), 1181 => to_unsigned(2647, 12), 1182 => to_unsigned(1999, 12), 1183 => to_unsigned(462, 12), 1184 => to_unsigned(1167, 12), 1185 => to_unsigned(1265, 12), 1186 => to_unsigned(2902, 12), 1187 => to_unsigned(2565, 12), 1188 => to_unsigned(1959, 12), 1189 => to_unsigned(1825, 12), 1190 => to_unsigned(677, 12), 1191 => to_unsigned(1945, 12), 1192 => to_unsigned(3914, 12), 1193 => to_unsigned(3798, 12), 1194 => to_unsigned(1180, 12), 1195 => to_unsigned(2586, 12), 1196 => to_unsigned(1556, 12), 1197 => to_unsigned(869, 12), 1198 => to_unsigned(2951, 12), 1199 => to_unsigned(251, 12), 1200 => to_unsigned(374, 12), 1201 => to_unsigned(1760, 12), 1202 => to_unsigned(386, 12), 1203 => to_unsigned(501, 12), 1204 => to_unsigned(557, 12), 1205 => to_unsigned(3181, 12), 1206 => to_unsigned(3662, 12), 1207 => to_unsigned(3464, 12), 1208 => to_unsigned(2857, 12), 1209 => to_unsigned(1934, 12), 1210 => to_unsigned(3204, 12), 1211 => to_unsigned(1186, 12), 1212 => to_unsigned(3271, 12), 1213 => to_unsigned(3217, 12), 1214 => to_unsigned(2182, 12), 1215 => to_unsigned(1146, 12), 1216 => to_unsigned(1172, 12), 1217 => to_unsigned(2759, 12), 1218 => to_unsigned(1296, 12), 1219 => to_unsigned(3069, 12), 1220 => to_unsigned(1364, 12), 1221 => to_unsigned(2378, 12), 1222 => to_unsigned(1821, 12), 1223 => to_unsigned(2266, 12), 1224 => to_unsigned(1497, 12), 1225 => to_unsigned(1577, 12), 1226 => to_unsigned(4060, 12), 1227 => to_unsigned(1357, 12), 1228 => to_unsigned(4052, 12), 1229 => to_unsigned(2905, 12), 1230 => to_unsigned(534, 12), 1231 => to_unsigned(3856, 12), 1232 => to_unsigned(2809, 12), 1233 => to_unsigned(3845, 12), 1234 => to_unsigned(482, 12), 1235 => to_unsigned(3693, 12), 1236 => to_unsigned(1629, 12), 1237 => to_unsigned(2586, 12), 1238 => to_unsigned(2034, 12), 1239 => to_unsigned(36, 12), 1240 => to_unsigned(1637, 12), 1241 => to_unsigned(2983, 12), 1242 => to_unsigned(1036, 12), 1243 => to_unsigned(550, 12), 1244 => to_unsigned(2915, 12), 1245 => to_unsigned(2500, 12), 1246 => to_unsigned(2479, 12), 1247 => to_unsigned(2398, 12), 1248 => to_unsigned(3187, 12), 1249 => to_unsigned(3475, 12), 1250 => to_unsigned(823, 12), 1251 => to_unsigned(2254, 12), 1252 => to_unsigned(502, 12), 1253 => to_unsigned(325, 12), 1254 => to_unsigned(251, 12), 1255 => to_unsigned(2898, 12), 1256 => to_unsigned(3262, 12), 1257 => to_unsigned(1677, 12), 1258 => to_unsigned(3258, 12), 1259 => to_unsigned(3102, 12), 1260 => to_unsigned(3810, 12), 1261 => to_unsigned(1937, 12), 1262 => to_unsigned(636, 12), 1263 => to_unsigned(237, 12), 1264 => to_unsigned(2168, 12), 1265 => to_unsigned(3997, 12), 1266 => to_unsigned(1864, 12), 1267 => to_unsigned(929, 12), 1268 => to_unsigned(2110, 12), 1269 => to_unsigned(576, 12), 1270 => to_unsigned(2370, 12), 1271 => to_unsigned(1445, 12), 1272 => to_unsigned(3299, 12), 1273 => to_unsigned(2502, 12), 1274 => to_unsigned(1780, 12), 1275 => to_unsigned(2272, 12), 1276 => to_unsigned(2948, 12), 1277 => to_unsigned(2930, 12), 1278 => to_unsigned(3210, 12), 1279 => to_unsigned(1200, 12), 1280 => to_unsigned(3396, 12), 1281 => to_unsigned(3603, 12), 1282 => to_unsigned(2533, 12), 1283 => to_unsigned(3295, 12), 1284 => to_unsigned(881, 12), 1285 => to_unsigned(3031, 12), 1286 => to_unsigned(3059, 12), 1287 => to_unsigned(2486, 12), 1288 => to_unsigned(1867, 12), 1289 => to_unsigned(2097, 12), 1290 => to_unsigned(1474, 12), 1291 => to_unsigned(332, 12), 1292 => to_unsigned(3096, 12), 1293 => to_unsigned(3649, 12), 1294 => to_unsigned(1478, 12), 1295 => to_unsigned(1677, 12), 1296 => to_unsigned(481, 12), 1297 => to_unsigned(3773, 12), 1298 => to_unsigned(1574, 12), 1299 => to_unsigned(383, 12), 1300 => to_unsigned(1734, 12), 1301 => to_unsigned(2023, 12), 1302 => to_unsigned(105, 12), 1303 => to_unsigned(2161, 12), 1304 => to_unsigned(247, 12), 1305 => to_unsigned(998, 12), 1306 => to_unsigned(3502, 12), 1307 => to_unsigned(3067, 12), 1308 => to_unsigned(3713, 12), 1309 => to_unsigned(3048, 12), 1310 => to_unsigned(3303, 12), 1311 => to_unsigned(2628, 12), 1312 => to_unsigned(2137, 12), 1313 => to_unsigned(2398, 12), 1314 => to_unsigned(32, 12), 1315 => to_unsigned(441, 12), 1316 => to_unsigned(2049, 12), 1317 => to_unsigned(2802, 12), 1318 => to_unsigned(475, 12), 1319 => to_unsigned(2364, 12), 1320 => to_unsigned(3101, 12), 1321 => to_unsigned(3997, 12), 1322 => to_unsigned(1806, 12), 1323 => to_unsigned(3296, 12), 1324 => to_unsigned(1725, 12), 1325 => to_unsigned(1161, 12), 1326 => to_unsigned(1886, 12), 1327 => to_unsigned(2889, 12), 1328 => to_unsigned(1690, 12), 1329 => to_unsigned(1136, 12), 1330 => to_unsigned(1485, 12), 1331 => to_unsigned(2565, 12), 1332 => to_unsigned(3664, 12), 1333 => to_unsigned(395, 12), 1334 => to_unsigned(778, 12), 1335 => to_unsigned(1946, 12), 1336 => to_unsigned(1413, 12), 1337 => to_unsigned(1600, 12), 1338 => to_unsigned(2577, 12), 1339 => to_unsigned(3044, 12), 1340 => to_unsigned(2357, 12), 1341 => to_unsigned(675, 12), 1342 => to_unsigned(1505, 12), 1343 => to_unsigned(842, 12), 1344 => to_unsigned(2168, 12), 1345 => to_unsigned(2560, 12), 1346 => to_unsigned(2904, 12), 1347 => to_unsigned(1486, 12), 1348 => to_unsigned(1845, 12), 1349 => to_unsigned(3187, 12), 1350 => to_unsigned(2470, 12), 1351 => to_unsigned(3110, 12), 1352 => to_unsigned(1280, 12), 1353 => to_unsigned(3141, 12), 1354 => to_unsigned(502, 12), 1355 => to_unsigned(531, 12), 1356 => to_unsigned(1713, 12), 1357 => to_unsigned(1669, 12), 1358 => to_unsigned(1718, 12), 1359 => to_unsigned(458, 12), 1360 => to_unsigned(2455, 12), 1361 => to_unsigned(866, 12), 1362 => to_unsigned(1593, 12), 1363 => to_unsigned(3849, 12), 1364 => to_unsigned(3569, 12), 1365 => to_unsigned(367, 12), 1366 => to_unsigned(1623, 12), 1367 => to_unsigned(2192, 12), 1368 => to_unsigned(3809, 12), 1369 => to_unsigned(3732, 12), 1370 => to_unsigned(3767, 12), 1371 => to_unsigned(3178, 12), 1372 => to_unsigned(206, 12), 1373 => to_unsigned(3517, 12), 1374 => to_unsigned(3875, 12), 1375 => to_unsigned(2527, 12), 1376 => to_unsigned(1610, 12), 1377 => to_unsigned(4019, 12), 1378 => to_unsigned(2645, 12), 1379 => to_unsigned(2101, 12), 1380 => to_unsigned(4016, 12), 1381 => to_unsigned(2321, 12), 1382 => to_unsigned(1165, 12), 1383 => to_unsigned(2744, 12), 1384 => to_unsigned(4049, 12), 1385 => to_unsigned(2498, 12), 1386 => to_unsigned(3051, 12), 1387 => to_unsigned(1692, 12), 1388 => to_unsigned(1615, 12), 1389 => to_unsigned(1370, 12), 1390 => to_unsigned(516, 12), 1391 => to_unsigned(3157, 12), 1392 => to_unsigned(3465, 12), 1393 => to_unsigned(493, 12), 1394 => to_unsigned(4069, 12), 1395 => to_unsigned(1270, 12), 1396 => to_unsigned(2666, 12), 1397 => to_unsigned(56, 12), 1398 => to_unsigned(2505, 12), 1399 => to_unsigned(813, 12), 1400 => to_unsigned(1265, 12), 1401 => to_unsigned(1267, 12), 1402 => to_unsigned(3348, 12), 1403 => to_unsigned(3121, 12), 1404 => to_unsigned(1673, 12), 1405 => to_unsigned(167, 12), 1406 => to_unsigned(485, 12), 1407 => to_unsigned(2475, 12), 1408 => to_unsigned(2651, 12), 1409 => to_unsigned(2951, 12), 1410 => to_unsigned(2138, 12), 1411 => to_unsigned(2253, 12), 1412 => to_unsigned(2009, 12), 1413 => to_unsigned(94, 12), 1414 => to_unsigned(2540, 12), 1415 => to_unsigned(2117, 12), 1416 => to_unsigned(2335, 12), 1417 => to_unsigned(1906, 12), 1418 => to_unsigned(630, 12), 1419 => to_unsigned(3290, 12), 1420 => to_unsigned(3893, 12), 1421 => to_unsigned(3024, 12), 1422 => to_unsigned(3020, 12), 1423 => to_unsigned(121, 12), 1424 => to_unsigned(2586, 12), 1425 => to_unsigned(442, 12), 1426 => to_unsigned(972, 12), 1427 => to_unsigned(792, 12), 1428 => to_unsigned(524, 12), 1429 => to_unsigned(3361, 12), 1430 => to_unsigned(917, 12), 1431 => to_unsigned(1199, 12), 1432 => to_unsigned(3060, 12), 1433 => to_unsigned(3453, 12), 1434 => to_unsigned(2085, 12), 1435 => to_unsigned(3169, 12), 1436 => to_unsigned(3979, 12), 1437 => to_unsigned(2941, 12), 1438 => to_unsigned(683, 12), 1439 => to_unsigned(2091, 12), 1440 => to_unsigned(3838, 12), 1441 => to_unsigned(1372, 12), 1442 => to_unsigned(3908, 12), 1443 => to_unsigned(42, 12), 1444 => to_unsigned(3656, 12), 1445 => to_unsigned(3269, 12), 1446 => to_unsigned(272, 12), 1447 => to_unsigned(971, 12), 1448 => to_unsigned(493, 12), 1449 => to_unsigned(916, 12), 1450 => to_unsigned(248, 12), 1451 => to_unsigned(2001, 12), 1452 => to_unsigned(1323, 12), 1453 => to_unsigned(2, 12), 1454 => to_unsigned(392, 12), 1455 => to_unsigned(2741, 12), 1456 => to_unsigned(2275, 12), 1457 => to_unsigned(3254, 12), 1458 => to_unsigned(1285, 12), 1459 => to_unsigned(823, 12), 1460 => to_unsigned(1732, 12), 1461 => to_unsigned(2691, 12), 1462 => to_unsigned(3652, 12), 1463 => to_unsigned(425, 12), 1464 => to_unsigned(1146, 12), 1465 => to_unsigned(2418, 12), 1466 => to_unsigned(3856, 12), 1467 => to_unsigned(2034, 12), 1468 => to_unsigned(1248, 12), 1469 => to_unsigned(883, 12), 1470 => to_unsigned(2940, 12), 1471 => to_unsigned(1874, 12), 1472 => to_unsigned(1819, 12), 1473 => to_unsigned(3061, 12), 1474 => to_unsigned(742, 12), 1475 => to_unsigned(3898, 12), 1476 => to_unsigned(3477, 12), 1477 => to_unsigned(1449, 12), 1478 => to_unsigned(3388, 12), 1479 => to_unsigned(2859, 12), 1480 => to_unsigned(2576, 12), 1481 => to_unsigned(2947, 12), 1482 => to_unsigned(115, 12), 1483 => to_unsigned(1335, 12), 1484 => to_unsigned(2765, 12), 1485 => to_unsigned(949, 12), 1486 => to_unsigned(1284, 12), 1487 => to_unsigned(3949, 12), 1488 => to_unsigned(2136, 12), 1489 => to_unsigned(695, 12), 1490 => to_unsigned(983, 12), 1491 => to_unsigned(2454, 12), 1492 => to_unsigned(3949, 12), 1493 => to_unsigned(1462, 12), 1494 => to_unsigned(2226, 12), 1495 => to_unsigned(280, 12), 1496 => to_unsigned(2563, 12), 1497 => to_unsigned(2114, 12), 1498 => to_unsigned(32, 12), 1499 => to_unsigned(1875, 12), 1500 => to_unsigned(447, 12), 1501 => to_unsigned(343, 12), 1502 => to_unsigned(3220, 12), 1503 => to_unsigned(498, 12), 1504 => to_unsigned(3725, 12), 1505 => to_unsigned(676, 12), 1506 => to_unsigned(2259, 12), 1507 => to_unsigned(1556, 12), 1508 => to_unsigned(2745, 12), 1509 => to_unsigned(3362, 12), 1510 => to_unsigned(999, 12), 1511 => to_unsigned(3, 12), 1512 => to_unsigned(3799, 12), 1513 => to_unsigned(828, 12), 1514 => to_unsigned(3509, 12), 1515 => to_unsigned(2274, 12), 1516 => to_unsigned(2361, 12), 1517 => to_unsigned(2139, 12), 1518 => to_unsigned(3585, 12), 1519 => to_unsigned(937, 12), 1520 => to_unsigned(473, 12), 1521 => to_unsigned(1043, 12), 1522 => to_unsigned(3887, 12), 1523 => to_unsigned(3690, 12), 1524 => to_unsigned(4030, 12), 1525 => to_unsigned(720, 12), 1526 => to_unsigned(1323, 12), 1527 => to_unsigned(3385, 12), 1528 => to_unsigned(2315, 12), 1529 => to_unsigned(685, 12), 1530 => to_unsigned(1940, 12), 1531 => to_unsigned(1949, 12), 1532 => to_unsigned(2986, 12), 1533 => to_unsigned(3655, 12), 1534 => to_unsigned(2610, 12), 1535 => to_unsigned(2187, 12), 1536 => to_unsigned(1612, 12), 1537 => to_unsigned(763, 12), 1538 => to_unsigned(530, 12), 1539 => to_unsigned(3014, 12), 1540 => to_unsigned(2159, 12), 1541 => to_unsigned(72, 12), 1542 => to_unsigned(4044, 12), 1543 => to_unsigned(3090, 12), 1544 => to_unsigned(3603, 12), 1545 => to_unsigned(576, 12), 1546 => to_unsigned(4084, 12), 1547 => to_unsigned(1930, 12), 1548 => to_unsigned(3430, 12), 1549 => to_unsigned(219, 12), 1550 => to_unsigned(348, 12), 1551 => to_unsigned(2319, 12), 1552 => to_unsigned(3432, 12), 1553 => to_unsigned(2979, 12), 1554 => to_unsigned(980, 12), 1555 => to_unsigned(3052, 12), 1556 => to_unsigned(2707, 12), 1557 => to_unsigned(623, 12), 1558 => to_unsigned(1814, 12), 1559 => to_unsigned(1855, 12), 1560 => to_unsigned(3469, 12), 1561 => to_unsigned(2429, 12), 1562 => to_unsigned(2188, 12), 1563 => to_unsigned(1475, 12), 1564 => to_unsigned(1025, 12), 1565 => to_unsigned(3543, 12), 1566 => to_unsigned(3012, 12), 1567 => to_unsigned(3968, 12), 1568 => to_unsigned(1609, 12), 1569 => to_unsigned(2773, 12), 1570 => to_unsigned(1426, 12), 1571 => to_unsigned(1052, 12), 1572 => to_unsigned(3484, 12), 1573 => to_unsigned(144, 12), 1574 => to_unsigned(601, 12), 1575 => to_unsigned(1158, 12), 1576 => to_unsigned(2731, 12), 1577 => to_unsigned(718, 12), 1578 => to_unsigned(932, 12), 1579 => to_unsigned(2764, 12), 1580 => to_unsigned(109, 12), 1581 => to_unsigned(3464, 12), 1582 => to_unsigned(2952, 12), 1583 => to_unsigned(3757, 12), 1584 => to_unsigned(50, 12), 1585 => to_unsigned(2092, 12), 1586 => to_unsigned(36, 12), 1587 => to_unsigned(1947, 12), 1588 => to_unsigned(2329, 12), 1589 => to_unsigned(3268, 12), 1590 => to_unsigned(3768, 12), 1591 => to_unsigned(3997, 12), 1592 => to_unsigned(286, 12), 1593 => to_unsigned(293, 12), 1594 => to_unsigned(101, 12), 1595 => to_unsigned(204, 12), 1596 => to_unsigned(2113, 12), 1597 => to_unsigned(2598, 12), 1598 => to_unsigned(398, 12), 1599 => to_unsigned(38, 12), 1600 => to_unsigned(3050, 12), 1601 => to_unsigned(3981, 12), 1602 => to_unsigned(677, 12), 1603 => to_unsigned(3805, 12), 1604 => to_unsigned(1246, 12), 1605 => to_unsigned(3367, 12), 1606 => to_unsigned(3579, 12), 1607 => to_unsigned(1035, 12), 1608 => to_unsigned(1279, 12), 1609 => to_unsigned(1057, 12), 1610 => to_unsigned(1979, 12), 1611 => to_unsigned(2421, 12), 1612 => to_unsigned(1852, 12), 1613 => to_unsigned(2223, 12), 1614 => to_unsigned(632, 12), 1615 => to_unsigned(1319, 12), 1616 => to_unsigned(2159, 12), 1617 => to_unsigned(1519, 12), 1618 => to_unsigned(489, 12), 1619 => to_unsigned(23, 12), 1620 => to_unsigned(1024, 12), 1621 => to_unsigned(1392, 12), 1622 => to_unsigned(117, 12), 1623 => to_unsigned(3194, 12), 1624 => to_unsigned(1014, 12), 1625 => to_unsigned(3842, 12), 1626 => to_unsigned(1067, 12), 1627 => to_unsigned(2383, 12), 1628 => to_unsigned(3846, 12), 1629 => to_unsigned(2249, 12), 1630 => to_unsigned(1917, 12), 1631 => to_unsigned(2572, 12), 1632 => to_unsigned(3639, 12), 1633 => to_unsigned(4015, 12), 1634 => to_unsigned(1762, 12), 1635 => to_unsigned(835, 12), 1636 => to_unsigned(3017, 12), 1637 => to_unsigned(282, 12), 1638 => to_unsigned(2479, 12), 1639 => to_unsigned(1521, 12), 1640 => to_unsigned(1367, 12), 1641 => to_unsigned(3949, 12), 1642 => to_unsigned(4030, 12), 1643 => to_unsigned(2832, 12), 1644 => to_unsigned(1676, 12), 1645 => to_unsigned(1100, 12), 1646 => to_unsigned(3384, 12), 1647 => to_unsigned(1758, 12), 1648 => to_unsigned(3628, 12), 1649 => to_unsigned(400, 12), 1650 => to_unsigned(3770, 12), 1651 => to_unsigned(2336, 12), 1652 => to_unsigned(1593, 12), 1653 => to_unsigned(3559, 12), 1654 => to_unsigned(3394, 12), 1655 => to_unsigned(2183, 12), 1656 => to_unsigned(2728, 12), 1657 => to_unsigned(2276, 12), 1658 => to_unsigned(440, 12), 1659 => to_unsigned(34, 12), 1660 => to_unsigned(2950, 12), 1661 => to_unsigned(882, 12), 1662 => to_unsigned(1526, 12), 1663 => to_unsigned(3789, 12), 1664 => to_unsigned(559, 12), 1665 => to_unsigned(2419, 12), 1666 => to_unsigned(3702, 12), 1667 => to_unsigned(486, 12), 1668 => to_unsigned(3768, 12), 1669 => to_unsigned(775, 12), 1670 => to_unsigned(3690, 12), 1671 => to_unsigned(174, 12), 1672 => to_unsigned(3507, 12), 1673 => to_unsigned(913, 12), 1674 => to_unsigned(1040, 12), 1675 => to_unsigned(4000, 12), 1676 => to_unsigned(2966, 12), 1677 => to_unsigned(1301, 12), 1678 => to_unsigned(4044, 12), 1679 => to_unsigned(429, 12), 1680 => to_unsigned(3602, 12), 1681 => to_unsigned(1680, 12), 1682 => to_unsigned(553, 12), 1683 => to_unsigned(2879, 12), 1684 => to_unsigned(2116, 12), 1685 => to_unsigned(1505, 12), 1686 => to_unsigned(2879, 12), 1687 => to_unsigned(3951, 12), 1688 => to_unsigned(166, 12), 1689 => to_unsigned(1259, 12), 1690 => to_unsigned(1766, 12), 1691 => to_unsigned(3082, 12), 1692 => to_unsigned(2439, 12), 1693 => to_unsigned(2646, 12), 1694 => to_unsigned(4038, 12), 1695 => to_unsigned(2846, 12), 1696 => to_unsigned(470, 12), 1697 => to_unsigned(3380, 12), 1698 => to_unsigned(690, 12), 1699 => to_unsigned(2370, 12), 1700 => to_unsigned(2060, 12), 1701 => to_unsigned(3357, 12), 1702 => to_unsigned(2619, 12), 1703 => to_unsigned(3682, 12), 1704 => to_unsigned(2323, 12), 1705 => to_unsigned(3352, 12), 1706 => to_unsigned(3789, 12), 1707 => to_unsigned(3645, 12), 1708 => to_unsigned(3801, 12), 1709 => to_unsigned(1876, 12), 1710 => to_unsigned(1396, 12), 1711 => to_unsigned(3831, 12), 1712 => to_unsigned(1300, 12), 1713 => to_unsigned(2620, 12), 1714 => to_unsigned(2616, 12), 1715 => to_unsigned(1449, 12), 1716 => to_unsigned(2977, 12), 1717 => to_unsigned(798, 12), 1718 => to_unsigned(2799, 12), 1719 => to_unsigned(1547, 12), 1720 => to_unsigned(3047, 12), 1721 => to_unsigned(2713, 12), 1722 => to_unsigned(2070, 12), 1723 => to_unsigned(2485, 12), 1724 => to_unsigned(4028, 12), 1725 => to_unsigned(335, 12), 1726 => to_unsigned(2233, 12), 1727 => to_unsigned(3712, 12), 1728 => to_unsigned(1221, 12), 1729 => to_unsigned(629, 12), 1730 => to_unsigned(1258, 12), 1731 => to_unsigned(3621, 12), 1732 => to_unsigned(3368, 12), 1733 => to_unsigned(2218, 12), 1734 => to_unsigned(3708, 12), 1735 => to_unsigned(2998, 12), 1736 => to_unsigned(770, 12), 1737 => to_unsigned(3752, 12), 1738 => to_unsigned(760, 12), 1739 => to_unsigned(708, 12), 1740 => to_unsigned(3198, 12), 1741 => to_unsigned(2105, 12), 1742 => to_unsigned(3113, 12), 1743 => to_unsigned(3787, 12), 1744 => to_unsigned(3569, 12), 1745 => to_unsigned(182, 12), 1746 => to_unsigned(3236, 12), 1747 => to_unsigned(2844, 12), 1748 => to_unsigned(948, 12), 1749 => to_unsigned(2401, 12), 1750 => to_unsigned(2569, 12), 1751 => to_unsigned(1151, 12), 1752 => to_unsigned(2819, 12), 1753 => to_unsigned(2654, 12), 1754 => to_unsigned(3019, 12), 1755 => to_unsigned(3933, 12), 1756 => to_unsigned(3622, 12), 1757 => to_unsigned(3695, 12), 1758 => to_unsigned(1808, 12), 1759 => to_unsigned(3694, 12), 1760 => to_unsigned(3344, 12), 1761 => to_unsigned(671, 12), 1762 => to_unsigned(2617, 12), 1763 => to_unsigned(2347, 12), 1764 => to_unsigned(1835, 12), 1765 => to_unsigned(2433, 12), 1766 => to_unsigned(1329, 12), 1767 => to_unsigned(3279, 12), 1768 => to_unsigned(3909, 12), 1769 => to_unsigned(2353, 12), 1770 => to_unsigned(1979, 12), 1771 => to_unsigned(517, 12), 1772 => to_unsigned(1026, 12), 1773 => to_unsigned(1504, 12), 1774 => to_unsigned(1026, 12), 1775 => to_unsigned(2833, 12), 1776 => to_unsigned(2758, 12), 1777 => to_unsigned(2719, 12), 1778 => to_unsigned(776, 12), 1779 => to_unsigned(3161, 12), 1780 => to_unsigned(887, 12), 1781 => to_unsigned(3162, 12), 1782 => to_unsigned(3494, 12), 1783 => to_unsigned(2305, 12), 1784 => to_unsigned(4028, 12), 1785 => to_unsigned(791, 12), 1786 => to_unsigned(3692, 12), 1787 => to_unsigned(783, 12), 1788 => to_unsigned(583, 12), 1789 => to_unsigned(3579, 12), 1790 => to_unsigned(2762, 12), 1791 => to_unsigned(2228, 12), 1792 => to_unsigned(443, 12), 1793 => to_unsigned(171, 12), 1794 => to_unsigned(2412, 12), 1795 => to_unsigned(1061, 12), 1796 => to_unsigned(2507, 12), 1797 => to_unsigned(1897, 12), 1798 => to_unsigned(2245, 12), 1799 => to_unsigned(378, 12), 1800 => to_unsigned(2224, 12), 1801 => to_unsigned(4063, 12), 1802 => to_unsigned(2848, 12), 1803 => to_unsigned(2897, 12), 1804 => to_unsigned(2148, 12), 1805 => to_unsigned(3531, 12), 1806 => to_unsigned(1369, 12), 1807 => to_unsigned(3191, 12), 1808 => to_unsigned(138, 12), 1809 => to_unsigned(819, 12), 1810 => to_unsigned(3408, 12), 1811 => to_unsigned(1102, 12), 1812 => to_unsigned(814, 12), 1813 => to_unsigned(2210, 12), 1814 => to_unsigned(3964, 12), 1815 => to_unsigned(1216, 12), 1816 => to_unsigned(360, 12), 1817 => to_unsigned(1422, 12), 1818 => to_unsigned(2588, 12), 1819 => to_unsigned(3166, 12), 1820 => to_unsigned(2332, 12), 1821 => to_unsigned(1649, 12), 1822 => to_unsigned(1599, 12), 1823 => to_unsigned(364, 12), 1824 => to_unsigned(585, 12), 1825 => to_unsigned(411, 12), 1826 => to_unsigned(3225, 12), 1827 => to_unsigned(3164, 12), 1828 => to_unsigned(2684, 12), 1829 => to_unsigned(2429, 12), 1830 => to_unsigned(4020, 12), 1831 => to_unsigned(885, 12), 1832 => to_unsigned(3294, 12), 1833 => to_unsigned(3406, 12), 1834 => to_unsigned(586, 12), 1835 => to_unsigned(3889, 12), 1836 => to_unsigned(1792, 12), 1837 => to_unsigned(555, 12), 1838 => to_unsigned(1559, 12), 1839 => to_unsigned(352, 12), 1840 => to_unsigned(2043, 12), 1841 => to_unsigned(2546, 12), 1842 => to_unsigned(355, 12), 1843 => to_unsigned(99, 12), 1844 => to_unsigned(1270, 12), 1845 => to_unsigned(1249, 12), 1846 => to_unsigned(1407, 12), 1847 => to_unsigned(342, 12), 1848 => to_unsigned(920, 12), 1849 => to_unsigned(3970, 12), 1850 => to_unsigned(693, 12), 1851 => to_unsigned(3927, 12), 1852 => to_unsigned(3597, 12), 1853 => to_unsigned(1852, 12), 1854 => to_unsigned(3587, 12), 1855 => to_unsigned(3751, 12), 1856 => to_unsigned(2951, 12), 1857 => to_unsigned(3630, 12), 1858 => to_unsigned(3685, 12), 1859 => to_unsigned(150, 12), 1860 => to_unsigned(2248, 12), 1861 => to_unsigned(2948, 12), 1862 => to_unsigned(546, 12), 1863 => to_unsigned(1727, 12), 1864 => to_unsigned(2439, 12), 1865 => to_unsigned(1715, 12), 1866 => to_unsigned(1302, 12), 1867 => to_unsigned(2993, 12), 1868 => to_unsigned(2595, 12), 1869 => to_unsigned(1220, 12), 1870 => to_unsigned(1348, 12), 1871 => to_unsigned(2841, 12), 1872 => to_unsigned(620, 12), 1873 => to_unsigned(481, 12), 1874 => to_unsigned(1525, 12), 1875 => to_unsigned(964, 12), 1876 => to_unsigned(1405, 12), 1877 => to_unsigned(3593, 12), 1878 => to_unsigned(1181, 12), 1879 => to_unsigned(868, 12), 1880 => to_unsigned(2979, 12), 1881 => to_unsigned(182, 12), 1882 => to_unsigned(1051, 12), 1883 => to_unsigned(2561, 12), 1884 => to_unsigned(406, 12), 1885 => to_unsigned(1736, 12), 1886 => to_unsigned(830, 12), 1887 => to_unsigned(488, 12), 1888 => to_unsigned(616, 12), 1889 => to_unsigned(3768, 12), 1890 => to_unsigned(338, 12), 1891 => to_unsigned(2671, 12), 1892 => to_unsigned(3105, 12), 1893 => to_unsigned(1041, 12), 1894 => to_unsigned(2806, 12), 1895 => to_unsigned(2805, 12), 1896 => to_unsigned(2025, 12), 1897 => to_unsigned(3366, 12), 1898 => to_unsigned(236, 12), 1899 => to_unsigned(316, 12), 1900 => to_unsigned(3060, 12), 1901 => to_unsigned(1205, 12), 1902 => to_unsigned(590, 12), 1903 => to_unsigned(3869, 12), 1904 => to_unsigned(319, 12), 1905 => to_unsigned(2813, 12), 1906 => to_unsigned(2040, 12), 1907 => to_unsigned(939, 12), 1908 => to_unsigned(3653, 12), 1909 => to_unsigned(2160, 12), 1910 => to_unsigned(2482, 12), 1911 => to_unsigned(2473, 12), 1912 => to_unsigned(2509, 12), 1913 => to_unsigned(428, 12), 1914 => to_unsigned(566, 12), 1915 => to_unsigned(1980, 12), 1916 => to_unsigned(2564, 12), 1917 => to_unsigned(3610, 12), 1918 => to_unsigned(2717, 12), 1919 => to_unsigned(3235, 12), 1920 => to_unsigned(858, 12), 1921 => to_unsigned(1993, 12), 1922 => to_unsigned(708, 12), 1923 => to_unsigned(1382, 12), 1924 => to_unsigned(3870, 12), 1925 => to_unsigned(3048, 12), 1926 => to_unsigned(1531, 12), 1927 => to_unsigned(3837, 12), 1928 => to_unsigned(2130, 12), 1929 => to_unsigned(1994, 12), 1930 => to_unsigned(597, 12), 1931 => to_unsigned(206, 12), 1932 => to_unsigned(4029, 12), 1933 => to_unsigned(3248, 12), 1934 => to_unsigned(444, 12), 1935 => to_unsigned(1550, 12), 1936 => to_unsigned(1380, 12), 1937 => to_unsigned(2313, 12), 1938 => to_unsigned(1243, 12), 1939 => to_unsigned(660, 12), 1940 => to_unsigned(1295, 12), 1941 => to_unsigned(3394, 12), 1942 => to_unsigned(2195, 12), 1943 => to_unsigned(790, 12), 1944 => to_unsigned(3190, 12), 1945 => to_unsigned(1408, 12), 1946 => to_unsigned(629, 12), 1947 => to_unsigned(3290, 12), 1948 => to_unsigned(1860, 12), 1949 => to_unsigned(1061, 12), 1950 => to_unsigned(1593, 12), 1951 => to_unsigned(2294, 12), 1952 => to_unsigned(1007, 12), 1953 => to_unsigned(2582, 12), 1954 => to_unsigned(1081, 12), 1955 => to_unsigned(2731, 12), 1956 => to_unsigned(3644, 12), 1957 => to_unsigned(547, 12), 1958 => to_unsigned(3532, 12), 1959 => to_unsigned(3283, 12), 1960 => to_unsigned(1657, 12), 1961 => to_unsigned(1623, 12), 1962 => to_unsigned(2075, 12), 1963 => to_unsigned(404, 12), 1964 => to_unsigned(2219, 12), 1965 => to_unsigned(3753, 12), 1966 => to_unsigned(1136, 12), 1967 => to_unsigned(895, 12), 1968 => to_unsigned(1597, 12), 1969 => to_unsigned(1974, 12), 1970 => to_unsigned(2358, 12), 1971 => to_unsigned(1659, 12), 1972 => to_unsigned(2324, 12), 1973 => to_unsigned(880, 12), 1974 => to_unsigned(1282, 12), 1975 => to_unsigned(2926, 12), 1976 => to_unsigned(249, 12), 1977 => to_unsigned(1303, 12), 1978 => to_unsigned(162, 12), 1979 => to_unsigned(442, 12), 1980 => to_unsigned(724, 12), 1981 => to_unsigned(512, 12), 1982 => to_unsigned(139, 12), 1983 => to_unsigned(3328, 12), 1984 => to_unsigned(2241, 12), 1985 => to_unsigned(2131, 12), 1986 => to_unsigned(1543, 12), 1987 => to_unsigned(2105, 12), 1988 => to_unsigned(1851, 12), 1989 => to_unsigned(2708, 12), 1990 => to_unsigned(2491, 12), 1991 => to_unsigned(2490, 12), 1992 => to_unsigned(1072, 12), 1993 => to_unsigned(1867, 12), 1994 => to_unsigned(1399, 12), 1995 => to_unsigned(200, 12), 1996 => to_unsigned(2928, 12), 1997 => to_unsigned(2852, 12), 1998 => to_unsigned(2361, 12), 1999 => to_unsigned(484, 12), 2000 => to_unsigned(928, 12), 2001 => to_unsigned(1707, 12), 2002 => to_unsigned(1609, 12), 2003 => to_unsigned(3893, 12), 2004 => to_unsigned(197, 12), 2005 => to_unsigned(277, 12), 2006 => to_unsigned(2950, 12), 2007 => to_unsigned(1174, 12), 2008 => to_unsigned(1933, 12), 2009 => to_unsigned(1901, 12), 2010 => to_unsigned(1476, 12), 2011 => to_unsigned(104, 12), 2012 => to_unsigned(3879, 12), 2013 => to_unsigned(1512, 12), 2014 => to_unsigned(940, 12), 2015 => to_unsigned(404, 12), 2016 => to_unsigned(987, 12), 2017 => to_unsigned(69, 12), 2018 => to_unsigned(4081, 12), 2019 => to_unsigned(1887, 12), 2020 => to_unsigned(3698, 12), 2021 => to_unsigned(838, 12), 2022 => to_unsigned(329, 12), 2023 => to_unsigned(2002, 12), 2024 => to_unsigned(3196, 12), 2025 => to_unsigned(2264, 12), 2026 => to_unsigned(1291, 12), 2027 => to_unsigned(1393, 12), 2028 => to_unsigned(3154, 12), 2029 => to_unsigned(2158, 12), 2030 => to_unsigned(3333, 12), 2031 => to_unsigned(1697, 12), 2032 => to_unsigned(1662, 12), 2033 => to_unsigned(3572, 12), 2034 => to_unsigned(3753, 12), 2035 => to_unsigned(4093, 12), 2036 => to_unsigned(2726, 12), 2037 => to_unsigned(2070, 12), 2038 => to_unsigned(3972, 12), 2039 => to_unsigned(1376, 12), 2040 => to_unsigned(874, 12), 2041 => to_unsigned(3365, 12), 2042 => to_unsigned(1620, 12), 2043 => to_unsigned(3069, 12), 2044 => to_unsigned(63, 12), 2045 => to_unsigned(774, 12), 2046 => to_unsigned(1392, 12), 2047 => to_unsigned(413, 12)),
            8 => (0 => to_unsigned(619, 12), 1 => to_unsigned(159, 12), 2 => to_unsigned(164, 12), 3 => to_unsigned(1083, 12), 4 => to_unsigned(2595, 12), 5 => to_unsigned(302, 12), 6 => to_unsigned(2613, 12), 7 => to_unsigned(3837, 12), 8 => to_unsigned(1152, 12), 9 => to_unsigned(3825, 12), 10 => to_unsigned(847, 12), 11 => to_unsigned(2169, 12), 12 => to_unsigned(2713, 12), 13 => to_unsigned(931, 12), 14 => to_unsigned(1387, 12), 15 => to_unsigned(2882, 12), 16 => to_unsigned(3908, 12), 17 => to_unsigned(1322, 12), 18 => to_unsigned(1045, 12), 19 => to_unsigned(3471, 12), 20 => to_unsigned(911, 12), 21 => to_unsigned(3850, 12), 22 => to_unsigned(2484, 12), 23 => to_unsigned(2993, 12), 24 => to_unsigned(3411, 12), 25 => to_unsigned(3654, 12), 26 => to_unsigned(155, 12), 27 => to_unsigned(1517, 12), 28 => to_unsigned(2899, 12), 29 => to_unsigned(3183, 12), 30 => to_unsigned(3633, 12), 31 => to_unsigned(93, 12), 32 => to_unsigned(2088, 12), 33 => to_unsigned(1304, 12), 34 => to_unsigned(2631, 12), 35 => to_unsigned(3238, 12), 36 => to_unsigned(2201, 12), 37 => to_unsigned(2284, 12), 38 => to_unsigned(2210, 12), 39 => to_unsigned(3463, 12), 40 => to_unsigned(786, 12), 41 => to_unsigned(3976, 12), 42 => to_unsigned(1961, 12), 43 => to_unsigned(1750, 12), 44 => to_unsigned(4030, 12), 45 => to_unsigned(2879, 12), 46 => to_unsigned(523, 12), 47 => to_unsigned(2283, 12), 48 => to_unsigned(339, 12), 49 => to_unsigned(3406, 12), 50 => to_unsigned(671, 12), 51 => to_unsigned(390, 12), 52 => to_unsigned(1064, 12), 53 => to_unsigned(2278, 12), 54 => to_unsigned(981, 12), 55 => to_unsigned(2425, 12), 56 => to_unsigned(4042, 12), 57 => to_unsigned(2281, 12), 58 => to_unsigned(3123, 12), 59 => to_unsigned(402, 12), 60 => to_unsigned(177, 12), 61 => to_unsigned(1851, 12), 62 => to_unsigned(1265, 12), 63 => to_unsigned(561, 12), 64 => to_unsigned(2516, 12), 65 => to_unsigned(511, 12), 66 => to_unsigned(108, 12), 67 => to_unsigned(1253, 12), 68 => to_unsigned(2230, 12), 69 => to_unsigned(905, 12), 70 => to_unsigned(1913, 12), 71 => to_unsigned(1963, 12), 72 => to_unsigned(3651, 12), 73 => to_unsigned(1465, 12), 74 => to_unsigned(3583, 12), 75 => to_unsigned(3000, 12), 76 => to_unsigned(643, 12), 77 => to_unsigned(2551, 12), 78 => to_unsigned(4034, 12), 79 => to_unsigned(2305, 12), 80 => to_unsigned(599, 12), 81 => to_unsigned(1596, 12), 82 => to_unsigned(1695, 12), 83 => to_unsigned(2546, 12), 84 => to_unsigned(2495, 12), 85 => to_unsigned(1591, 12), 86 => to_unsigned(1443, 12), 87 => to_unsigned(480, 12), 88 => to_unsigned(372, 12), 89 => to_unsigned(2987, 12), 90 => to_unsigned(2821, 12), 91 => to_unsigned(3238, 12), 92 => to_unsigned(1537, 12), 93 => to_unsigned(473, 12), 94 => to_unsigned(617, 12), 95 => to_unsigned(2531, 12), 96 => to_unsigned(3240, 12), 97 => to_unsigned(2849, 12), 98 => to_unsigned(2477, 12), 99 => to_unsigned(562, 12), 100 => to_unsigned(1743, 12), 101 => to_unsigned(17, 12), 102 => to_unsigned(2074, 12), 103 => to_unsigned(1867, 12), 104 => to_unsigned(2712, 12), 105 => to_unsigned(625, 12), 106 => to_unsigned(3188, 12), 107 => to_unsigned(3378, 12), 108 => to_unsigned(3900, 12), 109 => to_unsigned(2312, 12), 110 => to_unsigned(3505, 12), 111 => to_unsigned(156, 12), 112 => to_unsigned(301, 12), 113 => to_unsigned(3942, 12), 114 => to_unsigned(166, 12), 115 => to_unsigned(2320, 12), 116 => to_unsigned(2063, 12), 117 => to_unsigned(1515, 12), 118 => to_unsigned(3954, 12), 119 => to_unsigned(3883, 12), 120 => to_unsigned(3802, 12), 121 => to_unsigned(2085, 12), 122 => to_unsigned(3762, 12), 123 => to_unsigned(1541, 12), 124 => to_unsigned(643, 12), 125 => to_unsigned(1648, 12), 126 => to_unsigned(37, 12), 127 => to_unsigned(1751, 12), 128 => to_unsigned(766, 12), 129 => to_unsigned(3763, 12), 130 => to_unsigned(3711, 12), 131 => to_unsigned(2424, 12), 132 => to_unsigned(426, 12), 133 => to_unsigned(1800, 12), 134 => to_unsigned(873, 12), 135 => to_unsigned(3015, 12), 136 => to_unsigned(1723, 12), 137 => to_unsigned(3937, 12), 138 => to_unsigned(61, 12), 139 => to_unsigned(2681, 12), 140 => to_unsigned(1082, 12), 141 => to_unsigned(779, 12), 142 => to_unsigned(3184, 12), 143 => to_unsigned(2166, 12), 144 => to_unsigned(2613, 12), 145 => to_unsigned(3919, 12), 146 => to_unsigned(1946, 12), 147 => to_unsigned(3806, 12), 148 => to_unsigned(1693, 12), 149 => to_unsigned(210, 12), 150 => to_unsigned(2280, 12), 151 => to_unsigned(1129, 12), 152 => to_unsigned(2521, 12), 153 => to_unsigned(1056, 12), 154 => to_unsigned(2184, 12), 155 => to_unsigned(2272, 12), 156 => to_unsigned(1074, 12), 157 => to_unsigned(1789, 12), 158 => to_unsigned(460, 12), 159 => to_unsigned(896, 12), 160 => to_unsigned(2072, 12), 161 => to_unsigned(2303, 12), 162 => to_unsigned(1942, 12), 163 => to_unsigned(1501, 12), 164 => to_unsigned(1138, 12), 165 => to_unsigned(913, 12), 166 => to_unsigned(1468, 12), 167 => to_unsigned(3051, 12), 168 => to_unsigned(3384, 12), 169 => to_unsigned(1951, 12), 170 => to_unsigned(464, 12), 171 => to_unsigned(3543, 12), 172 => to_unsigned(2786, 12), 173 => to_unsigned(1241, 12), 174 => to_unsigned(2777, 12), 175 => to_unsigned(1864, 12), 176 => to_unsigned(1818, 12), 177 => to_unsigned(1095, 12), 178 => to_unsigned(2003, 12), 179 => to_unsigned(1636, 12), 180 => to_unsigned(3955, 12), 181 => to_unsigned(1915, 12), 182 => to_unsigned(3801, 12), 183 => to_unsigned(1315, 12), 184 => to_unsigned(1141, 12), 185 => to_unsigned(1997, 12), 186 => to_unsigned(530, 12), 187 => to_unsigned(1913, 12), 188 => to_unsigned(1370, 12), 189 => to_unsigned(2727, 12), 190 => to_unsigned(3315, 12), 191 => to_unsigned(1714, 12), 192 => to_unsigned(1997, 12), 193 => to_unsigned(2306, 12), 194 => to_unsigned(1747, 12), 195 => to_unsigned(3661, 12), 196 => to_unsigned(980, 12), 197 => to_unsigned(1196, 12), 198 => to_unsigned(681, 12), 199 => to_unsigned(47, 12), 200 => to_unsigned(196, 12), 201 => to_unsigned(3411, 12), 202 => to_unsigned(3257, 12), 203 => to_unsigned(554, 12), 204 => to_unsigned(2593, 12), 205 => to_unsigned(3691, 12), 206 => to_unsigned(1594, 12), 207 => to_unsigned(2577, 12), 208 => to_unsigned(2285, 12), 209 => to_unsigned(3687, 12), 210 => to_unsigned(193, 12), 211 => to_unsigned(1505, 12), 212 => to_unsigned(3396, 12), 213 => to_unsigned(2030, 12), 214 => to_unsigned(334, 12), 215 => to_unsigned(1603, 12), 216 => to_unsigned(3468, 12), 217 => to_unsigned(3007, 12), 218 => to_unsigned(3890, 12), 219 => to_unsigned(4040, 12), 220 => to_unsigned(1029, 12), 221 => to_unsigned(121, 12), 222 => to_unsigned(2527, 12), 223 => to_unsigned(2086, 12), 224 => to_unsigned(2196, 12), 225 => to_unsigned(507, 12), 226 => to_unsigned(1195, 12), 227 => to_unsigned(286, 12), 228 => to_unsigned(3827, 12), 229 => to_unsigned(3922, 12), 230 => to_unsigned(2801, 12), 231 => to_unsigned(3397, 12), 232 => to_unsigned(3577, 12), 233 => to_unsigned(478, 12), 234 => to_unsigned(527, 12), 235 => to_unsigned(1069, 12), 236 => to_unsigned(852, 12), 237 => to_unsigned(1766, 12), 238 => to_unsigned(1394, 12), 239 => to_unsigned(1448, 12), 240 => to_unsigned(794, 12), 241 => to_unsigned(4019, 12), 242 => to_unsigned(2555, 12), 243 => to_unsigned(1842, 12), 244 => to_unsigned(2109, 12), 245 => to_unsigned(1585, 12), 246 => to_unsigned(2527, 12), 247 => to_unsigned(575, 12), 248 => to_unsigned(3908, 12), 249 => to_unsigned(1268, 12), 250 => to_unsigned(658, 12), 251 => to_unsigned(596, 12), 252 => to_unsigned(3184, 12), 253 => to_unsigned(3485, 12), 254 => to_unsigned(3678, 12), 255 => to_unsigned(3276, 12), 256 => to_unsigned(3291, 12), 257 => to_unsigned(3669, 12), 258 => to_unsigned(3644, 12), 259 => to_unsigned(306, 12), 260 => to_unsigned(2256, 12), 261 => to_unsigned(1650, 12), 262 => to_unsigned(2226, 12), 263 => to_unsigned(3263, 12), 264 => to_unsigned(3401, 12), 265 => to_unsigned(3403, 12), 266 => to_unsigned(2918, 12), 267 => to_unsigned(932, 12), 268 => to_unsigned(2559, 12), 269 => to_unsigned(1579, 12), 270 => to_unsigned(3446, 12), 271 => to_unsigned(599, 12), 272 => to_unsigned(2818, 12), 273 => to_unsigned(126, 12), 274 => to_unsigned(1225, 12), 275 => to_unsigned(3289, 12), 276 => to_unsigned(2920, 12), 277 => to_unsigned(2920, 12), 278 => to_unsigned(1757, 12), 279 => to_unsigned(3293, 12), 280 => to_unsigned(2605, 12), 281 => to_unsigned(2137, 12), 282 => to_unsigned(1322, 12), 283 => to_unsigned(3975, 12), 284 => to_unsigned(3513, 12), 285 => to_unsigned(3641, 12), 286 => to_unsigned(1702, 12), 287 => to_unsigned(3835, 12), 288 => to_unsigned(484, 12), 289 => to_unsigned(1979, 12), 290 => to_unsigned(3654, 12), 291 => to_unsigned(1553, 12), 292 => to_unsigned(2861, 12), 293 => to_unsigned(378, 12), 294 => to_unsigned(331, 12), 295 => to_unsigned(3442, 12), 296 => to_unsigned(3583, 12), 297 => to_unsigned(2378, 12), 298 => to_unsigned(3954, 12), 299 => to_unsigned(4073, 12), 300 => to_unsigned(651, 12), 301 => to_unsigned(143, 12), 302 => to_unsigned(1233, 12), 303 => to_unsigned(2732, 12), 304 => to_unsigned(1879, 12), 305 => to_unsigned(3518, 12), 306 => to_unsigned(1313, 12), 307 => to_unsigned(905, 12), 308 => to_unsigned(456, 12), 309 => to_unsigned(1300, 12), 310 => to_unsigned(623, 12), 311 => to_unsigned(3884, 12), 312 => to_unsigned(3197, 12), 313 => to_unsigned(60, 12), 314 => to_unsigned(77, 12), 315 => to_unsigned(3499, 12), 316 => to_unsigned(598, 12), 317 => to_unsigned(122, 12), 318 => to_unsigned(3055, 12), 319 => to_unsigned(1717, 12), 320 => to_unsigned(31, 12), 321 => to_unsigned(1382, 12), 322 => to_unsigned(2696, 12), 323 => to_unsigned(2983, 12), 324 => to_unsigned(270, 12), 325 => to_unsigned(3389, 12), 326 => to_unsigned(455, 12), 327 => to_unsigned(3730, 12), 328 => to_unsigned(1117, 12), 329 => to_unsigned(1545, 12), 330 => to_unsigned(2434, 12), 331 => to_unsigned(2262, 12), 332 => to_unsigned(922, 12), 333 => to_unsigned(1810, 12), 334 => to_unsigned(1224, 12), 335 => to_unsigned(2836, 12), 336 => to_unsigned(3520, 12), 337 => to_unsigned(2811, 12), 338 => to_unsigned(2742, 12), 339 => to_unsigned(778, 12), 340 => to_unsigned(678, 12), 341 => to_unsigned(2142, 12), 342 => to_unsigned(948, 12), 343 => to_unsigned(676, 12), 344 => to_unsigned(3770, 12), 345 => to_unsigned(1136, 12), 346 => to_unsigned(1517, 12), 347 => to_unsigned(279, 12), 348 => to_unsigned(2621, 12), 349 => to_unsigned(1469, 12), 350 => to_unsigned(2013, 12), 351 => to_unsigned(158, 12), 352 => to_unsigned(3506, 12), 353 => to_unsigned(1217, 12), 354 => to_unsigned(27, 12), 355 => to_unsigned(2456, 12), 356 => to_unsigned(3118, 12), 357 => to_unsigned(2852, 12), 358 => to_unsigned(1203, 12), 359 => to_unsigned(3365, 12), 360 => to_unsigned(3736, 12), 361 => to_unsigned(585, 12), 362 => to_unsigned(2627, 12), 363 => to_unsigned(3273, 12), 364 => to_unsigned(2574, 12), 365 => to_unsigned(2975, 12), 366 => to_unsigned(4020, 12), 367 => to_unsigned(2427, 12), 368 => to_unsigned(2799, 12), 369 => to_unsigned(69, 12), 370 => to_unsigned(3619, 12), 371 => to_unsigned(90, 12), 372 => to_unsigned(684, 12), 373 => to_unsigned(589, 12), 374 => to_unsigned(3284, 12), 375 => to_unsigned(1498, 12), 376 => to_unsigned(1312, 12), 377 => to_unsigned(689, 12), 378 => to_unsigned(1141, 12), 379 => to_unsigned(2871, 12), 380 => to_unsigned(3498, 12), 381 => to_unsigned(2671, 12), 382 => to_unsigned(1122, 12), 383 => to_unsigned(1487, 12), 384 => to_unsigned(1236, 12), 385 => to_unsigned(3295, 12), 386 => to_unsigned(2307, 12), 387 => to_unsigned(2833, 12), 388 => to_unsigned(3224, 12), 389 => to_unsigned(1401, 12), 390 => to_unsigned(3811, 12), 391 => to_unsigned(454, 12), 392 => to_unsigned(612, 12), 393 => to_unsigned(2356, 12), 394 => to_unsigned(2157, 12), 395 => to_unsigned(3029, 12), 396 => to_unsigned(3970, 12), 397 => to_unsigned(3491, 12), 398 => to_unsigned(273, 12), 399 => to_unsigned(141, 12), 400 => to_unsigned(785, 12), 401 => to_unsigned(2552, 12), 402 => to_unsigned(2148, 12), 403 => to_unsigned(3891, 12), 404 => to_unsigned(3383, 12), 405 => to_unsigned(3589, 12), 406 => to_unsigned(4069, 12), 407 => to_unsigned(462, 12), 408 => to_unsigned(234, 12), 409 => to_unsigned(1828, 12), 410 => to_unsigned(1679, 12), 411 => to_unsigned(2630, 12), 412 => to_unsigned(3526, 12), 413 => to_unsigned(2682, 12), 414 => to_unsigned(1924, 12), 415 => to_unsigned(899, 12), 416 => to_unsigned(1262, 12), 417 => to_unsigned(1453, 12), 418 => to_unsigned(956, 12), 419 => to_unsigned(3102, 12), 420 => to_unsigned(4015, 12), 421 => to_unsigned(3361, 12), 422 => to_unsigned(3548, 12), 423 => to_unsigned(2873, 12), 424 => to_unsigned(1599, 12), 425 => to_unsigned(2879, 12), 426 => to_unsigned(2903, 12), 427 => to_unsigned(1078, 12), 428 => to_unsigned(3838, 12), 429 => to_unsigned(847, 12), 430 => to_unsigned(3355, 12), 431 => to_unsigned(3825, 12), 432 => to_unsigned(693, 12), 433 => to_unsigned(3357, 12), 434 => to_unsigned(2846, 12), 435 => to_unsigned(3727, 12), 436 => to_unsigned(3324, 12), 437 => to_unsigned(1111, 12), 438 => to_unsigned(2990, 12), 439 => to_unsigned(2416, 12), 440 => to_unsigned(2207, 12), 441 => to_unsigned(677, 12), 442 => to_unsigned(864, 12), 443 => to_unsigned(3839, 12), 444 => to_unsigned(3034, 12), 445 => to_unsigned(1746, 12), 446 => to_unsigned(3684, 12), 447 => to_unsigned(1589, 12), 448 => to_unsigned(2837, 12), 449 => to_unsigned(731, 12), 450 => to_unsigned(3534, 12), 451 => to_unsigned(2305, 12), 452 => to_unsigned(1251, 12), 453 => to_unsigned(591, 12), 454 => to_unsigned(2105, 12), 455 => to_unsigned(3423, 12), 456 => to_unsigned(918, 12), 457 => to_unsigned(1827, 12), 458 => to_unsigned(2909, 12), 459 => to_unsigned(1667, 12), 460 => to_unsigned(2483, 12), 461 => to_unsigned(379, 12), 462 => to_unsigned(54, 12), 463 => to_unsigned(1184, 12), 464 => to_unsigned(1783, 12), 465 => to_unsigned(949, 12), 466 => to_unsigned(3432, 12), 467 => to_unsigned(1625, 12), 468 => to_unsigned(1343, 12), 469 => to_unsigned(1778, 12), 470 => to_unsigned(2325, 12), 471 => to_unsigned(1651, 12), 472 => to_unsigned(3380, 12), 473 => to_unsigned(1154, 12), 474 => to_unsigned(1931, 12), 475 => to_unsigned(3822, 12), 476 => to_unsigned(965, 12), 477 => to_unsigned(1534, 12), 478 => to_unsigned(31, 12), 479 => to_unsigned(746, 12), 480 => to_unsigned(4083, 12), 481 => to_unsigned(1693, 12), 482 => to_unsigned(3517, 12), 483 => to_unsigned(1274, 12), 484 => to_unsigned(2950, 12), 485 => to_unsigned(1701, 12), 486 => to_unsigned(3072, 12), 487 => to_unsigned(3335, 12), 488 => to_unsigned(1694, 12), 489 => to_unsigned(1993, 12), 490 => to_unsigned(3938, 12), 491 => to_unsigned(1719, 12), 492 => to_unsigned(980, 12), 493 => to_unsigned(1745, 12), 494 => to_unsigned(1404, 12), 495 => to_unsigned(1813, 12), 496 => to_unsigned(1689, 12), 497 => to_unsigned(790, 12), 498 => to_unsigned(1964, 12), 499 => to_unsigned(3337, 12), 500 => to_unsigned(1261, 12), 501 => to_unsigned(1003, 12), 502 => to_unsigned(790, 12), 503 => to_unsigned(3509, 12), 504 => to_unsigned(633, 12), 505 => to_unsigned(638, 12), 506 => to_unsigned(3364, 12), 507 => to_unsigned(3544, 12), 508 => to_unsigned(826, 12), 509 => to_unsigned(3968, 12), 510 => to_unsigned(2393, 12), 511 => to_unsigned(2760, 12), 512 => to_unsigned(1718, 12), 513 => to_unsigned(1551, 12), 514 => to_unsigned(2912, 12), 515 => to_unsigned(496, 12), 516 => to_unsigned(203, 12), 517 => to_unsigned(1646, 12), 518 => to_unsigned(1788, 12), 519 => to_unsigned(3022, 12), 520 => to_unsigned(1468, 12), 521 => to_unsigned(2791, 12), 522 => to_unsigned(1706, 12), 523 => to_unsigned(880, 12), 524 => to_unsigned(422, 12), 525 => to_unsigned(1710, 12), 526 => to_unsigned(365, 12), 527 => to_unsigned(80, 12), 528 => to_unsigned(1746, 12), 529 => to_unsigned(3645, 12), 530 => to_unsigned(1564, 12), 531 => to_unsigned(704, 12), 532 => to_unsigned(1760, 12), 533 => to_unsigned(194, 12), 534 => to_unsigned(48, 12), 535 => to_unsigned(1599, 12), 536 => to_unsigned(914, 12), 537 => to_unsigned(1509, 12), 538 => to_unsigned(3759, 12), 539 => to_unsigned(1232, 12), 540 => to_unsigned(2981, 12), 541 => to_unsigned(90, 12), 542 => to_unsigned(2694, 12), 543 => to_unsigned(3251, 12), 544 => to_unsigned(587, 12), 545 => to_unsigned(3713, 12), 546 => to_unsigned(755, 12), 547 => to_unsigned(2945, 12), 548 => to_unsigned(2073, 12), 549 => to_unsigned(3564, 12), 550 => to_unsigned(3773, 12), 551 => to_unsigned(1597, 12), 552 => to_unsigned(2388, 12), 553 => to_unsigned(358, 12), 554 => to_unsigned(3660, 12), 555 => to_unsigned(2629, 12), 556 => to_unsigned(2790, 12), 557 => to_unsigned(947, 12), 558 => to_unsigned(1362, 12), 559 => to_unsigned(3992, 12), 560 => to_unsigned(4067, 12), 561 => to_unsigned(420, 12), 562 => to_unsigned(1704, 12), 563 => to_unsigned(2893, 12), 564 => to_unsigned(1710, 12), 565 => to_unsigned(3748, 12), 566 => to_unsigned(2203, 12), 567 => to_unsigned(659, 12), 568 => to_unsigned(449, 12), 569 => to_unsigned(3557, 12), 570 => to_unsigned(1319, 12), 571 => to_unsigned(3318, 12), 572 => to_unsigned(542, 12), 573 => to_unsigned(1243, 12), 574 => to_unsigned(2086, 12), 575 => to_unsigned(1520, 12), 576 => to_unsigned(758, 12), 577 => to_unsigned(754, 12), 578 => to_unsigned(74, 12), 579 => to_unsigned(1329, 12), 580 => to_unsigned(3843, 12), 581 => to_unsigned(2517, 12), 582 => to_unsigned(3586, 12), 583 => to_unsigned(2981, 12), 584 => to_unsigned(3204, 12), 585 => to_unsigned(3241, 12), 586 => to_unsigned(1604, 12), 587 => to_unsigned(1309, 12), 588 => to_unsigned(189, 12), 589 => to_unsigned(1501, 12), 590 => to_unsigned(3612, 12), 591 => to_unsigned(332, 12), 592 => to_unsigned(2067, 12), 593 => to_unsigned(2697, 12), 594 => to_unsigned(3533, 12), 595 => to_unsigned(3124, 12), 596 => to_unsigned(470, 12), 597 => to_unsigned(2342, 12), 598 => to_unsigned(804, 12), 599 => to_unsigned(1051, 12), 600 => to_unsigned(2862, 12), 601 => to_unsigned(2777, 12), 602 => to_unsigned(3663, 12), 603 => to_unsigned(3145, 12), 604 => to_unsigned(3687, 12), 605 => to_unsigned(2848, 12), 606 => to_unsigned(1348, 12), 607 => to_unsigned(3586, 12), 608 => to_unsigned(3747, 12), 609 => to_unsigned(3985, 12), 610 => to_unsigned(138, 12), 611 => to_unsigned(2686, 12), 612 => to_unsigned(1983, 12), 613 => to_unsigned(1480, 12), 614 => to_unsigned(1746, 12), 615 => to_unsigned(293, 12), 616 => to_unsigned(3054, 12), 617 => to_unsigned(1483, 12), 618 => to_unsigned(1439, 12), 619 => to_unsigned(4085, 12), 620 => to_unsigned(3685, 12), 621 => to_unsigned(993, 12), 622 => to_unsigned(3024, 12), 623 => to_unsigned(2679, 12), 624 => to_unsigned(4014, 12), 625 => to_unsigned(3705, 12), 626 => to_unsigned(2994, 12), 627 => to_unsigned(2979, 12), 628 => to_unsigned(3404, 12), 629 => to_unsigned(1476, 12), 630 => to_unsigned(2021, 12), 631 => to_unsigned(2919, 12), 632 => to_unsigned(1274, 12), 633 => to_unsigned(2785, 12), 634 => to_unsigned(1409, 12), 635 => to_unsigned(3328, 12), 636 => to_unsigned(2310, 12), 637 => to_unsigned(810, 12), 638 => to_unsigned(3112, 12), 639 => to_unsigned(2717, 12), 640 => to_unsigned(3639, 12), 641 => to_unsigned(3173, 12), 642 => to_unsigned(2945, 12), 643 => to_unsigned(1428, 12), 644 => to_unsigned(3459, 12), 645 => to_unsigned(3270, 12), 646 => to_unsigned(935, 12), 647 => to_unsigned(2934, 12), 648 => to_unsigned(3213, 12), 649 => to_unsigned(2837, 12), 650 => to_unsigned(424, 12), 651 => to_unsigned(3688, 12), 652 => to_unsigned(2118, 12), 653 => to_unsigned(2185, 12), 654 => to_unsigned(3561, 12), 655 => to_unsigned(1365, 12), 656 => to_unsigned(2684, 12), 657 => to_unsigned(4073, 12), 658 => to_unsigned(2906, 12), 659 => to_unsigned(283, 12), 660 => to_unsigned(2467, 12), 661 => to_unsigned(656, 12), 662 => to_unsigned(2469, 12), 663 => to_unsigned(2428, 12), 664 => to_unsigned(1859, 12), 665 => to_unsigned(2044, 12), 666 => to_unsigned(1532, 12), 667 => to_unsigned(3400, 12), 668 => to_unsigned(3171, 12), 669 => to_unsigned(593, 12), 670 => to_unsigned(1404, 12), 671 => to_unsigned(1850, 12), 672 => to_unsigned(1141, 12), 673 => to_unsigned(582, 12), 674 => to_unsigned(1032, 12), 675 => to_unsigned(1653, 12), 676 => to_unsigned(3044, 12), 677 => to_unsigned(4045, 12), 678 => to_unsigned(344, 12), 679 => to_unsigned(3832, 12), 680 => to_unsigned(3758, 12), 681 => to_unsigned(2866, 12), 682 => to_unsigned(2021, 12), 683 => to_unsigned(1148, 12), 684 => to_unsigned(93, 12), 685 => to_unsigned(1523, 12), 686 => to_unsigned(3979, 12), 687 => to_unsigned(3439, 12), 688 => to_unsigned(1564, 12), 689 => to_unsigned(2248, 12), 690 => to_unsigned(3961, 12), 691 => to_unsigned(751, 12), 692 => to_unsigned(277, 12), 693 => to_unsigned(4004, 12), 694 => to_unsigned(296, 12), 695 => to_unsigned(3489, 12), 696 => to_unsigned(2662, 12), 697 => to_unsigned(60, 12), 698 => to_unsigned(2929, 12), 699 => to_unsigned(2494, 12), 700 => to_unsigned(1155, 12), 701 => to_unsigned(3919, 12), 702 => to_unsigned(2301, 12), 703 => to_unsigned(2212, 12), 704 => to_unsigned(3289, 12), 705 => to_unsigned(1735, 12), 706 => to_unsigned(1618, 12), 707 => to_unsigned(2709, 12), 708 => to_unsigned(2751, 12), 709 => to_unsigned(126, 12), 710 => to_unsigned(4025, 12), 711 => to_unsigned(1027, 12), 712 => to_unsigned(3119, 12), 713 => to_unsigned(2770, 12), 714 => to_unsigned(3415, 12), 715 => to_unsigned(1636, 12), 716 => to_unsigned(3503, 12), 717 => to_unsigned(864, 12), 718 => to_unsigned(3991, 12), 719 => to_unsigned(186, 12), 720 => to_unsigned(3295, 12), 721 => to_unsigned(3565, 12), 722 => to_unsigned(1450, 12), 723 => to_unsigned(1501, 12), 724 => to_unsigned(2768, 12), 725 => to_unsigned(1380, 12), 726 => to_unsigned(1966, 12), 727 => to_unsigned(2500, 12), 728 => to_unsigned(518, 12), 729 => to_unsigned(177, 12), 730 => to_unsigned(2773, 12), 731 => to_unsigned(1136, 12), 732 => to_unsigned(4035, 12), 733 => to_unsigned(2179, 12), 734 => to_unsigned(2528, 12), 735 => to_unsigned(3006, 12), 736 => to_unsigned(2513, 12), 737 => to_unsigned(3093, 12), 738 => to_unsigned(365, 12), 739 => to_unsigned(134, 12), 740 => to_unsigned(2857, 12), 741 => to_unsigned(3028, 12), 742 => to_unsigned(1884, 12), 743 => to_unsigned(3584, 12), 744 => to_unsigned(133, 12), 745 => to_unsigned(2610, 12), 746 => to_unsigned(3101, 12), 747 => to_unsigned(3313, 12), 748 => to_unsigned(3139, 12), 749 => to_unsigned(3058, 12), 750 => to_unsigned(988, 12), 751 => to_unsigned(1003, 12), 752 => to_unsigned(3640, 12), 753 => to_unsigned(2195, 12), 754 => to_unsigned(386, 12), 755 => to_unsigned(1994, 12), 756 => to_unsigned(3090, 12), 757 => to_unsigned(3275, 12), 758 => to_unsigned(3634, 12), 759 => to_unsigned(3115, 12), 760 => to_unsigned(62, 12), 761 => to_unsigned(3712, 12), 762 => to_unsigned(3210, 12), 763 => to_unsigned(2735, 12), 764 => to_unsigned(912, 12), 765 => to_unsigned(2524, 12), 766 => to_unsigned(3883, 12), 767 => to_unsigned(3980, 12), 768 => to_unsigned(3293, 12), 769 => to_unsigned(465, 12), 770 => to_unsigned(906, 12), 771 => to_unsigned(2497, 12), 772 => to_unsigned(1669, 12), 773 => to_unsigned(679, 12), 774 => to_unsigned(732, 12), 775 => to_unsigned(1149, 12), 776 => to_unsigned(648, 12), 777 => to_unsigned(992, 12), 778 => to_unsigned(1832, 12), 779 => to_unsigned(1551, 12), 780 => to_unsigned(2305, 12), 781 => to_unsigned(4006, 12), 782 => to_unsigned(4001, 12), 783 => to_unsigned(1711, 12), 784 => to_unsigned(958, 12), 785 => to_unsigned(367, 12), 786 => to_unsigned(3767, 12), 787 => to_unsigned(3789, 12), 788 => to_unsigned(811, 12), 789 => to_unsigned(4089, 12), 790 => to_unsigned(3742, 12), 791 => to_unsigned(4041, 12), 792 => to_unsigned(3115, 12), 793 => to_unsigned(1524, 12), 794 => to_unsigned(285, 12), 795 => to_unsigned(646, 12), 796 => to_unsigned(1043, 12), 797 => to_unsigned(1814, 12), 798 => to_unsigned(790, 12), 799 => to_unsigned(680, 12), 800 => to_unsigned(3414, 12), 801 => to_unsigned(203, 12), 802 => to_unsigned(3061, 12), 803 => to_unsigned(1860, 12), 804 => to_unsigned(1294, 12), 805 => to_unsigned(2084, 12), 806 => to_unsigned(329, 12), 807 => to_unsigned(3597, 12), 808 => to_unsigned(1999, 12), 809 => to_unsigned(3722, 12), 810 => to_unsigned(2391, 12), 811 => to_unsigned(810, 12), 812 => to_unsigned(1660, 12), 813 => to_unsigned(723, 12), 814 => to_unsigned(3160, 12), 815 => to_unsigned(3801, 12), 816 => to_unsigned(4010, 12), 817 => to_unsigned(1988, 12), 818 => to_unsigned(1152, 12), 819 => to_unsigned(4028, 12), 820 => to_unsigned(3685, 12), 821 => to_unsigned(1111, 12), 822 => to_unsigned(3710, 12), 823 => to_unsigned(3910, 12), 824 => to_unsigned(1883, 12), 825 => to_unsigned(2294, 12), 826 => to_unsigned(3656, 12), 827 => to_unsigned(3271, 12), 828 => to_unsigned(45, 12), 829 => to_unsigned(2286, 12), 830 => to_unsigned(341, 12), 831 => to_unsigned(2186, 12), 832 => to_unsigned(3077, 12), 833 => to_unsigned(2152, 12), 834 => to_unsigned(1173, 12), 835 => to_unsigned(441, 12), 836 => to_unsigned(512, 12), 837 => to_unsigned(2428, 12), 838 => to_unsigned(1079, 12), 839 => to_unsigned(1726, 12), 840 => to_unsigned(3565, 12), 841 => to_unsigned(57, 12), 842 => to_unsigned(3114, 12), 843 => to_unsigned(1097, 12), 844 => to_unsigned(3515, 12), 845 => to_unsigned(1891, 12), 846 => to_unsigned(2388, 12), 847 => to_unsigned(2984, 12), 848 => to_unsigned(2049, 12), 849 => to_unsigned(3680, 12), 850 => to_unsigned(3124, 12), 851 => to_unsigned(2404, 12), 852 => to_unsigned(3196, 12), 853 => to_unsigned(1956, 12), 854 => to_unsigned(4054, 12), 855 => to_unsigned(593, 12), 856 => to_unsigned(3992, 12), 857 => to_unsigned(3946, 12), 858 => to_unsigned(1067, 12), 859 => to_unsigned(3242, 12), 860 => to_unsigned(2828, 12), 861 => to_unsigned(1831, 12), 862 => to_unsigned(3298, 12), 863 => to_unsigned(1119, 12), 864 => to_unsigned(1279, 12), 865 => to_unsigned(3925, 12), 866 => to_unsigned(2473, 12), 867 => to_unsigned(2880, 12), 868 => to_unsigned(287, 12), 869 => to_unsigned(1111, 12), 870 => to_unsigned(1885, 12), 871 => to_unsigned(1375, 12), 872 => to_unsigned(2114, 12), 873 => to_unsigned(3749, 12), 874 => to_unsigned(1326, 12), 875 => to_unsigned(16, 12), 876 => to_unsigned(1855, 12), 877 => to_unsigned(2040, 12), 878 => to_unsigned(3018, 12), 879 => to_unsigned(3354, 12), 880 => to_unsigned(1620, 12), 881 => to_unsigned(1941, 12), 882 => to_unsigned(2752, 12), 883 => to_unsigned(2983, 12), 884 => to_unsigned(1538, 12), 885 => to_unsigned(3877, 12), 886 => to_unsigned(3918, 12), 887 => to_unsigned(602, 12), 888 => to_unsigned(2507, 12), 889 => to_unsigned(2705, 12), 890 => to_unsigned(1796, 12), 891 => to_unsigned(3193, 12), 892 => to_unsigned(1704, 12), 893 => to_unsigned(898, 12), 894 => to_unsigned(254, 12), 895 => to_unsigned(2332, 12), 896 => to_unsigned(2688, 12), 897 => to_unsigned(2739, 12), 898 => to_unsigned(837, 12), 899 => to_unsigned(3507, 12), 900 => to_unsigned(3326, 12), 901 => to_unsigned(2220, 12), 902 => to_unsigned(2335, 12), 903 => to_unsigned(3248, 12), 904 => to_unsigned(1919, 12), 905 => to_unsigned(1594, 12), 906 => to_unsigned(921, 12), 907 => to_unsigned(2098, 12), 908 => to_unsigned(2583, 12), 909 => to_unsigned(774, 12), 910 => to_unsigned(3498, 12), 911 => to_unsigned(2863, 12), 912 => to_unsigned(2316, 12), 913 => to_unsigned(1079, 12), 914 => to_unsigned(3625, 12), 915 => to_unsigned(1258, 12), 916 => to_unsigned(692, 12), 917 => to_unsigned(1066, 12), 918 => to_unsigned(3739, 12), 919 => to_unsigned(484, 12), 920 => to_unsigned(1068, 12), 921 => to_unsigned(4030, 12), 922 => to_unsigned(2039, 12), 923 => to_unsigned(928, 12), 924 => to_unsigned(2539, 12), 925 => to_unsigned(3798, 12), 926 => to_unsigned(3585, 12), 927 => to_unsigned(3679, 12), 928 => to_unsigned(1864, 12), 929 => to_unsigned(915, 12), 930 => to_unsigned(1172, 12), 931 => to_unsigned(2878, 12), 932 => to_unsigned(2048, 12), 933 => to_unsigned(2411, 12), 934 => to_unsigned(1207, 12), 935 => to_unsigned(1553, 12), 936 => to_unsigned(787, 12), 937 => to_unsigned(3781, 12), 938 => to_unsigned(2658, 12), 939 => to_unsigned(3356, 12), 940 => to_unsigned(4026, 12), 941 => to_unsigned(797, 12), 942 => to_unsigned(2535, 12), 943 => to_unsigned(3149, 12), 944 => to_unsigned(685, 12), 945 => to_unsigned(3704, 12), 946 => to_unsigned(1887, 12), 947 => to_unsigned(3823, 12), 948 => to_unsigned(506, 12), 949 => to_unsigned(1719, 12), 950 => to_unsigned(154, 12), 951 => to_unsigned(1832, 12), 952 => to_unsigned(1690, 12), 953 => to_unsigned(1365, 12), 954 => to_unsigned(1088, 12), 955 => to_unsigned(1104, 12), 956 => to_unsigned(3225, 12), 957 => to_unsigned(2590, 12), 958 => to_unsigned(3290, 12), 959 => to_unsigned(2243, 12), 960 => to_unsigned(4036, 12), 961 => to_unsigned(1413, 12), 962 => to_unsigned(2914, 12), 963 => to_unsigned(558, 12), 964 => to_unsigned(456, 12), 965 => to_unsigned(2122, 12), 966 => to_unsigned(366, 12), 967 => to_unsigned(3746, 12), 968 => to_unsigned(880, 12), 969 => to_unsigned(3177, 12), 970 => to_unsigned(2418, 12), 971 => to_unsigned(638, 12), 972 => to_unsigned(973, 12), 973 => to_unsigned(316, 12), 974 => to_unsigned(2386, 12), 975 => to_unsigned(2236, 12), 976 => to_unsigned(4042, 12), 977 => to_unsigned(830, 12), 978 => to_unsigned(268, 12), 979 => to_unsigned(3817, 12), 980 => to_unsigned(1187, 12), 981 => to_unsigned(3769, 12), 982 => to_unsigned(2056, 12), 983 => to_unsigned(3186, 12), 984 => to_unsigned(413, 12), 985 => to_unsigned(182, 12), 986 => to_unsigned(388, 12), 987 => to_unsigned(3754, 12), 988 => to_unsigned(1245, 12), 989 => to_unsigned(944, 12), 990 => to_unsigned(1675, 12), 991 => to_unsigned(55, 12), 992 => to_unsigned(2230, 12), 993 => to_unsigned(3726, 12), 994 => to_unsigned(2786, 12), 995 => to_unsigned(2919, 12), 996 => to_unsigned(2688, 12), 997 => to_unsigned(3176, 12), 998 => to_unsigned(844, 12), 999 => to_unsigned(1021, 12), 1000 => to_unsigned(3732, 12), 1001 => to_unsigned(2360, 12), 1002 => to_unsigned(3101, 12), 1003 => to_unsigned(2638, 12), 1004 => to_unsigned(1772, 12), 1005 => to_unsigned(3222, 12), 1006 => to_unsigned(84, 12), 1007 => to_unsigned(2689, 12), 1008 => to_unsigned(3503, 12), 1009 => to_unsigned(1598, 12), 1010 => to_unsigned(2339, 12), 1011 => to_unsigned(3449, 12), 1012 => to_unsigned(794, 12), 1013 => to_unsigned(1525, 12), 1014 => to_unsigned(53, 12), 1015 => to_unsigned(809, 12), 1016 => to_unsigned(2547, 12), 1017 => to_unsigned(843, 12), 1018 => to_unsigned(1292, 12), 1019 => to_unsigned(2663, 12), 1020 => to_unsigned(3789, 12), 1021 => to_unsigned(2159, 12), 1022 => to_unsigned(580, 12), 1023 => to_unsigned(3971, 12), 1024 => to_unsigned(839, 12), 1025 => to_unsigned(1258, 12), 1026 => to_unsigned(2891, 12), 1027 => to_unsigned(3565, 12), 1028 => to_unsigned(171, 12), 1029 => to_unsigned(2248, 12), 1030 => to_unsigned(2586, 12), 1031 => to_unsigned(2240, 12), 1032 => to_unsigned(2695, 12), 1033 => to_unsigned(4032, 12), 1034 => to_unsigned(1270, 12), 1035 => to_unsigned(1156, 12), 1036 => to_unsigned(1124, 12), 1037 => to_unsigned(2607, 12), 1038 => to_unsigned(1502, 12), 1039 => to_unsigned(2229, 12), 1040 => to_unsigned(4044, 12), 1041 => to_unsigned(2062, 12), 1042 => to_unsigned(3776, 12), 1043 => to_unsigned(2095, 12), 1044 => to_unsigned(1489, 12), 1045 => to_unsigned(1493, 12), 1046 => to_unsigned(4045, 12), 1047 => to_unsigned(3838, 12), 1048 => to_unsigned(936, 12), 1049 => to_unsigned(3355, 12), 1050 => to_unsigned(1403, 12), 1051 => to_unsigned(3253, 12), 1052 => to_unsigned(382, 12), 1053 => to_unsigned(1976, 12), 1054 => to_unsigned(739, 12), 1055 => to_unsigned(2394, 12), 1056 => to_unsigned(3350, 12), 1057 => to_unsigned(344, 12), 1058 => to_unsigned(2841, 12), 1059 => to_unsigned(3483, 12), 1060 => to_unsigned(2768, 12), 1061 => to_unsigned(1349, 12), 1062 => to_unsigned(1361, 12), 1063 => to_unsigned(1891, 12), 1064 => to_unsigned(3552, 12), 1065 => to_unsigned(1143, 12), 1066 => to_unsigned(1683, 12), 1067 => to_unsigned(3552, 12), 1068 => to_unsigned(3229, 12), 1069 => to_unsigned(402, 12), 1070 => to_unsigned(1686, 12), 1071 => to_unsigned(496, 12), 1072 => to_unsigned(2117, 12), 1073 => to_unsigned(2195, 12), 1074 => to_unsigned(1757, 12), 1075 => to_unsigned(1708, 12), 1076 => to_unsigned(2214, 12), 1077 => to_unsigned(1131, 12), 1078 => to_unsigned(891, 12), 1079 => to_unsigned(3126, 12), 1080 => to_unsigned(3527, 12), 1081 => to_unsigned(3613, 12), 1082 => to_unsigned(1010, 12), 1083 => to_unsigned(3462, 12), 1084 => to_unsigned(394, 12), 1085 => to_unsigned(3812, 12), 1086 => to_unsigned(2990, 12), 1087 => to_unsigned(1655, 12), 1088 => to_unsigned(3440, 12), 1089 => to_unsigned(2762, 12), 1090 => to_unsigned(2901, 12), 1091 => to_unsigned(277, 12), 1092 => to_unsigned(3582, 12), 1093 => to_unsigned(4067, 12), 1094 => to_unsigned(925, 12), 1095 => to_unsigned(1058, 12), 1096 => to_unsigned(2204, 12), 1097 => to_unsigned(1793, 12), 1098 => to_unsigned(3760, 12), 1099 => to_unsigned(1849, 12), 1100 => to_unsigned(717, 12), 1101 => to_unsigned(1191, 12), 1102 => to_unsigned(1085, 12), 1103 => to_unsigned(4, 12), 1104 => to_unsigned(322, 12), 1105 => to_unsigned(585, 12), 1106 => to_unsigned(556, 12), 1107 => to_unsigned(1707, 12), 1108 => to_unsigned(594, 12), 1109 => to_unsigned(2948, 12), 1110 => to_unsigned(3452, 12), 1111 => to_unsigned(1768, 12), 1112 => to_unsigned(2032, 12), 1113 => to_unsigned(481, 12), 1114 => to_unsigned(228, 12), 1115 => to_unsigned(2170, 12), 1116 => to_unsigned(684, 12), 1117 => to_unsigned(2788, 12), 1118 => to_unsigned(4019, 12), 1119 => to_unsigned(1393, 12), 1120 => to_unsigned(1381, 12), 1121 => to_unsigned(614, 12), 1122 => to_unsigned(1295, 12), 1123 => to_unsigned(703, 12), 1124 => to_unsigned(3761, 12), 1125 => to_unsigned(3006, 12), 1126 => to_unsigned(1548, 12), 1127 => to_unsigned(2216, 12), 1128 => to_unsigned(4052, 12), 1129 => to_unsigned(3088, 12), 1130 => to_unsigned(1873, 12), 1131 => to_unsigned(730, 12), 1132 => to_unsigned(3941, 12), 1133 => to_unsigned(2222, 12), 1134 => to_unsigned(1513, 12), 1135 => to_unsigned(1655, 12), 1136 => to_unsigned(556, 12), 1137 => to_unsigned(2667, 12), 1138 => to_unsigned(3691, 12), 1139 => to_unsigned(431, 12), 1140 => to_unsigned(2528, 12), 1141 => to_unsigned(277, 12), 1142 => to_unsigned(3696, 12), 1143 => to_unsigned(162, 12), 1144 => to_unsigned(2889, 12), 1145 => to_unsigned(3325, 12), 1146 => to_unsigned(3180, 12), 1147 => to_unsigned(40, 12), 1148 => to_unsigned(797, 12), 1149 => to_unsigned(3420, 12), 1150 => to_unsigned(1671, 12), 1151 => to_unsigned(727, 12), 1152 => to_unsigned(2754, 12), 1153 => to_unsigned(2442, 12), 1154 => to_unsigned(2585, 12), 1155 => to_unsigned(2645, 12), 1156 => to_unsigned(1320, 12), 1157 => to_unsigned(1542, 12), 1158 => to_unsigned(2514, 12), 1159 => to_unsigned(3216, 12), 1160 => to_unsigned(2187, 12), 1161 => to_unsigned(685, 12), 1162 => to_unsigned(3736, 12), 1163 => to_unsigned(790, 12), 1164 => to_unsigned(955, 12), 1165 => to_unsigned(2115, 12), 1166 => to_unsigned(1003, 12), 1167 => to_unsigned(94, 12), 1168 => to_unsigned(1965, 12), 1169 => to_unsigned(2152, 12), 1170 => to_unsigned(1799, 12), 1171 => to_unsigned(3842, 12), 1172 => to_unsigned(1821, 12), 1173 => to_unsigned(4040, 12), 1174 => to_unsigned(3889, 12), 1175 => to_unsigned(3704, 12), 1176 => to_unsigned(1949, 12), 1177 => to_unsigned(770, 12), 1178 => to_unsigned(3334, 12), 1179 => to_unsigned(3518, 12), 1180 => to_unsigned(1588, 12), 1181 => to_unsigned(90, 12), 1182 => to_unsigned(2817, 12), 1183 => to_unsigned(381, 12), 1184 => to_unsigned(3679, 12), 1185 => to_unsigned(1768, 12), 1186 => to_unsigned(1835, 12), 1187 => to_unsigned(2666, 12), 1188 => to_unsigned(317, 12), 1189 => to_unsigned(367, 12), 1190 => to_unsigned(3917, 12), 1191 => to_unsigned(430, 12), 1192 => to_unsigned(3573, 12), 1193 => to_unsigned(1736, 12), 1194 => to_unsigned(837, 12), 1195 => to_unsigned(2891, 12), 1196 => to_unsigned(1311, 12), 1197 => to_unsigned(1570, 12), 1198 => to_unsigned(2624, 12), 1199 => to_unsigned(3582, 12), 1200 => to_unsigned(1292, 12), 1201 => to_unsigned(2476, 12), 1202 => to_unsigned(1876, 12), 1203 => to_unsigned(372, 12), 1204 => to_unsigned(3214, 12), 1205 => to_unsigned(1634, 12), 1206 => to_unsigned(1053, 12), 1207 => to_unsigned(861, 12), 1208 => to_unsigned(2870, 12), 1209 => to_unsigned(1309, 12), 1210 => to_unsigned(3969, 12), 1211 => to_unsigned(210, 12), 1212 => to_unsigned(539, 12), 1213 => to_unsigned(3273, 12), 1214 => to_unsigned(2603, 12), 1215 => to_unsigned(1524, 12), 1216 => to_unsigned(1532, 12), 1217 => to_unsigned(2136, 12), 1218 => to_unsigned(3432, 12), 1219 => to_unsigned(413, 12), 1220 => to_unsigned(2316, 12), 1221 => to_unsigned(1185, 12), 1222 => to_unsigned(2506, 12), 1223 => to_unsigned(63, 12), 1224 => to_unsigned(945, 12), 1225 => to_unsigned(1676, 12), 1226 => to_unsigned(2182, 12), 1227 => to_unsigned(3526, 12), 1228 => to_unsigned(2042, 12), 1229 => to_unsigned(1054, 12), 1230 => to_unsigned(618, 12), 1231 => to_unsigned(3653, 12), 1232 => to_unsigned(2916, 12), 1233 => to_unsigned(3101, 12), 1234 => to_unsigned(3610, 12), 1235 => to_unsigned(1468, 12), 1236 => to_unsigned(797, 12), 1237 => to_unsigned(2066, 12), 1238 => to_unsigned(4092, 12), 1239 => to_unsigned(1607, 12), 1240 => to_unsigned(2708, 12), 1241 => to_unsigned(600, 12), 1242 => to_unsigned(3616, 12), 1243 => to_unsigned(191, 12), 1244 => to_unsigned(734, 12), 1245 => to_unsigned(4059, 12), 1246 => to_unsigned(3096, 12), 1247 => to_unsigned(1276, 12), 1248 => to_unsigned(2691, 12), 1249 => to_unsigned(2693, 12), 1250 => to_unsigned(2445, 12), 1251 => to_unsigned(1259, 12), 1252 => to_unsigned(2373, 12), 1253 => to_unsigned(1425, 12), 1254 => to_unsigned(856, 12), 1255 => to_unsigned(1619, 12), 1256 => to_unsigned(1456, 12), 1257 => to_unsigned(1625, 12), 1258 => to_unsigned(1401, 12), 1259 => to_unsigned(1156, 12), 1260 => to_unsigned(145, 12), 1261 => to_unsigned(510, 12), 1262 => to_unsigned(2593, 12), 1263 => to_unsigned(1816, 12), 1264 => to_unsigned(2404, 12), 1265 => to_unsigned(740, 12), 1266 => to_unsigned(805, 12), 1267 => to_unsigned(2591, 12), 1268 => to_unsigned(212, 12), 1269 => to_unsigned(564, 12), 1270 => to_unsigned(1491, 12), 1271 => to_unsigned(3730, 12), 1272 => to_unsigned(1742, 12), 1273 => to_unsigned(668, 12), 1274 => to_unsigned(1906, 12), 1275 => to_unsigned(1498, 12), 1276 => to_unsigned(3704, 12), 1277 => to_unsigned(2426, 12), 1278 => to_unsigned(719, 12), 1279 => to_unsigned(2792, 12), 1280 => to_unsigned(2049, 12), 1281 => to_unsigned(3789, 12), 1282 => to_unsigned(1918, 12), 1283 => to_unsigned(2590, 12), 1284 => to_unsigned(2427, 12), 1285 => to_unsigned(3025, 12), 1286 => to_unsigned(1332, 12), 1287 => to_unsigned(191, 12), 1288 => to_unsigned(1189, 12), 1289 => to_unsigned(2726, 12), 1290 => to_unsigned(1566, 12), 1291 => to_unsigned(42, 12), 1292 => to_unsigned(2033, 12), 1293 => to_unsigned(1380, 12), 1294 => to_unsigned(1802, 12), 1295 => to_unsigned(1000, 12), 1296 => to_unsigned(3537, 12), 1297 => to_unsigned(1838, 12), 1298 => to_unsigned(1400, 12), 1299 => to_unsigned(4021, 12), 1300 => to_unsigned(1527, 12), 1301 => to_unsigned(1296, 12), 1302 => to_unsigned(570, 12), 1303 => to_unsigned(1940, 12), 1304 => to_unsigned(2862, 12), 1305 => to_unsigned(206, 12), 1306 => to_unsigned(2016, 12), 1307 => to_unsigned(1932, 12), 1308 => to_unsigned(1483, 12), 1309 => to_unsigned(3204, 12), 1310 => to_unsigned(2065, 12), 1311 => to_unsigned(3603, 12), 1312 => to_unsigned(1582, 12), 1313 => to_unsigned(1043, 12), 1314 => to_unsigned(2569, 12), 1315 => to_unsigned(264, 12), 1316 => to_unsigned(2538, 12), 1317 => to_unsigned(20, 12), 1318 => to_unsigned(2663, 12), 1319 => to_unsigned(1710, 12), 1320 => to_unsigned(2543, 12), 1321 => to_unsigned(2170, 12), 1322 => to_unsigned(1008, 12), 1323 => to_unsigned(982, 12), 1324 => to_unsigned(3206, 12), 1325 => to_unsigned(2163, 12), 1326 => to_unsigned(799, 12), 1327 => to_unsigned(3161, 12), 1328 => to_unsigned(3302, 12), 1329 => to_unsigned(4066, 12), 1330 => to_unsigned(1593, 12), 1331 => to_unsigned(1737, 12), 1332 => to_unsigned(4049, 12), 1333 => to_unsigned(1043, 12), 1334 => to_unsigned(3988, 12), 1335 => to_unsigned(1468, 12), 1336 => to_unsigned(3791, 12), 1337 => to_unsigned(3341, 12), 1338 => to_unsigned(2808, 12), 1339 => to_unsigned(1328, 12), 1340 => to_unsigned(195, 12), 1341 => to_unsigned(1798, 12), 1342 => to_unsigned(2827, 12), 1343 => to_unsigned(3194, 12), 1344 => to_unsigned(47, 12), 1345 => to_unsigned(3599, 12), 1346 => to_unsigned(1103, 12), 1347 => to_unsigned(584, 12), 1348 => to_unsigned(3877, 12), 1349 => to_unsigned(2866, 12), 1350 => to_unsigned(3281, 12), 1351 => to_unsigned(1180, 12), 1352 => to_unsigned(3542, 12), 1353 => to_unsigned(929, 12), 1354 => to_unsigned(636, 12), 1355 => to_unsigned(4013, 12), 1356 => to_unsigned(709, 12), 1357 => to_unsigned(2114, 12), 1358 => to_unsigned(2903, 12), 1359 => to_unsigned(3007, 12), 1360 => to_unsigned(2976, 12), 1361 => to_unsigned(468, 12), 1362 => to_unsigned(3582, 12), 1363 => to_unsigned(2839, 12), 1364 => to_unsigned(270, 12), 1365 => to_unsigned(71, 12), 1366 => to_unsigned(709, 12), 1367 => to_unsigned(1012, 12), 1368 => to_unsigned(1203, 12), 1369 => to_unsigned(679, 12), 1370 => to_unsigned(1417, 12), 1371 => to_unsigned(34, 12), 1372 => to_unsigned(1971, 12), 1373 => to_unsigned(3519, 12), 1374 => to_unsigned(1658, 12), 1375 => to_unsigned(1254, 12), 1376 => to_unsigned(3641, 12), 1377 => to_unsigned(2015, 12), 1378 => to_unsigned(1179, 12), 1379 => to_unsigned(3513, 12), 1380 => to_unsigned(1624, 12), 1381 => to_unsigned(1189, 12), 1382 => to_unsigned(303, 12), 1383 => to_unsigned(3830, 12), 1384 => to_unsigned(3262, 12), 1385 => to_unsigned(1324, 12), 1386 => to_unsigned(1043, 12), 1387 => to_unsigned(1137, 12), 1388 => to_unsigned(2798, 12), 1389 => to_unsigned(3956, 12), 1390 => to_unsigned(3588, 12), 1391 => to_unsigned(1928, 12), 1392 => to_unsigned(2992, 12), 1393 => to_unsigned(3837, 12), 1394 => to_unsigned(303, 12), 1395 => to_unsigned(1652, 12), 1396 => to_unsigned(1320, 12), 1397 => to_unsigned(3850, 12), 1398 => to_unsigned(2594, 12), 1399 => to_unsigned(3770, 12), 1400 => to_unsigned(438, 12), 1401 => to_unsigned(3117, 12), 1402 => to_unsigned(2572, 12), 1403 => to_unsigned(3646, 12), 1404 => to_unsigned(3330, 12), 1405 => to_unsigned(158, 12), 1406 => to_unsigned(4015, 12), 1407 => to_unsigned(967, 12), 1408 => to_unsigned(526, 12), 1409 => to_unsigned(1668, 12), 1410 => to_unsigned(75, 12), 1411 => to_unsigned(3448, 12), 1412 => to_unsigned(3417, 12), 1413 => to_unsigned(1785, 12), 1414 => to_unsigned(29, 12), 1415 => to_unsigned(1587, 12), 1416 => to_unsigned(2576, 12), 1417 => to_unsigned(2309, 12), 1418 => to_unsigned(714, 12), 1419 => to_unsigned(638, 12), 1420 => to_unsigned(957, 12), 1421 => to_unsigned(1309, 12), 1422 => to_unsigned(1545, 12), 1423 => to_unsigned(644, 12), 1424 => to_unsigned(3425, 12), 1425 => to_unsigned(2798, 12), 1426 => to_unsigned(270, 12), 1427 => to_unsigned(1875, 12), 1428 => to_unsigned(2650, 12), 1429 => to_unsigned(1616, 12), 1430 => to_unsigned(220, 12), 1431 => to_unsigned(3440, 12), 1432 => to_unsigned(1252, 12), 1433 => to_unsigned(2526, 12), 1434 => to_unsigned(2505, 12), 1435 => to_unsigned(1312, 12), 1436 => to_unsigned(2000, 12), 1437 => to_unsigned(280, 12), 1438 => to_unsigned(1110, 12), 1439 => to_unsigned(870, 12), 1440 => to_unsigned(1487, 12), 1441 => to_unsigned(163, 12), 1442 => to_unsigned(3632, 12), 1443 => to_unsigned(2704, 12), 1444 => to_unsigned(1269, 12), 1445 => to_unsigned(1803, 12), 1446 => to_unsigned(1076, 12), 1447 => to_unsigned(3542, 12), 1448 => to_unsigned(1233, 12), 1449 => to_unsigned(2614, 12), 1450 => to_unsigned(1234, 12), 1451 => to_unsigned(1252, 12), 1452 => to_unsigned(1758, 12), 1453 => to_unsigned(952, 12), 1454 => to_unsigned(3583, 12), 1455 => to_unsigned(1785, 12), 1456 => to_unsigned(22, 12), 1457 => to_unsigned(2216, 12), 1458 => to_unsigned(912, 12), 1459 => to_unsigned(396, 12), 1460 => to_unsigned(3239, 12), 1461 => to_unsigned(278, 12), 1462 => to_unsigned(3014, 12), 1463 => to_unsigned(3285, 12), 1464 => to_unsigned(2018, 12), 1465 => to_unsigned(1752, 12), 1466 => to_unsigned(1018, 12), 1467 => to_unsigned(3017, 12), 1468 => to_unsigned(1911, 12), 1469 => to_unsigned(378, 12), 1470 => to_unsigned(3519, 12), 1471 => to_unsigned(1603, 12), 1472 => to_unsigned(2100, 12), 1473 => to_unsigned(3662, 12), 1474 => to_unsigned(913, 12), 1475 => to_unsigned(3990, 12), 1476 => to_unsigned(3374, 12), 1477 => to_unsigned(543, 12), 1478 => to_unsigned(1585, 12), 1479 => to_unsigned(3869, 12), 1480 => to_unsigned(777, 12), 1481 => to_unsigned(3164, 12), 1482 => to_unsigned(1972, 12), 1483 => to_unsigned(1, 12), 1484 => to_unsigned(2197, 12), 1485 => to_unsigned(227, 12), 1486 => to_unsigned(1057, 12), 1487 => to_unsigned(2402, 12), 1488 => to_unsigned(2443, 12), 1489 => to_unsigned(3704, 12), 1490 => to_unsigned(1733, 12), 1491 => to_unsigned(1194, 12), 1492 => to_unsigned(1075, 12), 1493 => to_unsigned(1165, 12), 1494 => to_unsigned(3238, 12), 1495 => to_unsigned(303, 12), 1496 => to_unsigned(3086, 12), 1497 => to_unsigned(159, 12), 1498 => to_unsigned(2109, 12), 1499 => to_unsigned(4060, 12), 1500 => to_unsigned(220, 12), 1501 => to_unsigned(2777, 12), 1502 => to_unsigned(2291, 12), 1503 => to_unsigned(3573, 12), 1504 => to_unsigned(834, 12), 1505 => to_unsigned(3325, 12), 1506 => to_unsigned(3283, 12), 1507 => to_unsigned(3117, 12), 1508 => to_unsigned(298, 12), 1509 => to_unsigned(3222, 12), 1510 => to_unsigned(2203, 12), 1511 => to_unsigned(907, 12), 1512 => to_unsigned(2425, 12), 1513 => to_unsigned(3638, 12), 1514 => to_unsigned(925, 12), 1515 => to_unsigned(1648, 12), 1516 => to_unsigned(619, 12), 1517 => to_unsigned(2381, 12), 1518 => to_unsigned(1189, 12), 1519 => to_unsigned(3252, 12), 1520 => to_unsigned(222, 12), 1521 => to_unsigned(2659, 12), 1522 => to_unsigned(81, 12), 1523 => to_unsigned(1568, 12), 1524 => to_unsigned(686, 12), 1525 => to_unsigned(1595, 12), 1526 => to_unsigned(902, 12), 1527 => to_unsigned(921, 12), 1528 => to_unsigned(473, 12), 1529 => to_unsigned(1223, 12), 1530 => to_unsigned(3687, 12), 1531 => to_unsigned(3487, 12), 1532 => to_unsigned(103, 12), 1533 => to_unsigned(2701, 12), 1534 => to_unsigned(1715, 12), 1535 => to_unsigned(3096, 12), 1536 => to_unsigned(3281, 12), 1537 => to_unsigned(1527, 12), 1538 => to_unsigned(1722, 12), 1539 => to_unsigned(1885, 12), 1540 => to_unsigned(3606, 12), 1541 => to_unsigned(3484, 12), 1542 => to_unsigned(1896, 12), 1543 => to_unsigned(1844, 12), 1544 => to_unsigned(1486, 12), 1545 => to_unsigned(3432, 12), 1546 => to_unsigned(2969, 12), 1547 => to_unsigned(2287, 12), 1548 => to_unsigned(3563, 12), 1549 => to_unsigned(2324, 12), 1550 => to_unsigned(963, 12), 1551 => to_unsigned(1227, 12), 1552 => to_unsigned(253, 12), 1553 => to_unsigned(1421, 12), 1554 => to_unsigned(3072, 12), 1555 => to_unsigned(1509, 12), 1556 => to_unsigned(2834, 12), 1557 => to_unsigned(2345, 12), 1558 => to_unsigned(3840, 12), 1559 => to_unsigned(3148, 12), 1560 => to_unsigned(1185, 12), 1561 => to_unsigned(1822, 12), 1562 => to_unsigned(1667, 12), 1563 => to_unsigned(2467, 12), 1564 => to_unsigned(1050, 12), 1565 => to_unsigned(2430, 12), 1566 => to_unsigned(2896, 12), 1567 => to_unsigned(3628, 12), 1568 => to_unsigned(1966, 12), 1569 => to_unsigned(2691, 12), 1570 => to_unsigned(2153, 12), 1571 => to_unsigned(1979, 12), 1572 => to_unsigned(960, 12), 1573 => to_unsigned(641, 12), 1574 => to_unsigned(3335, 12), 1575 => to_unsigned(2654, 12), 1576 => to_unsigned(3416, 12), 1577 => to_unsigned(2463, 12), 1578 => to_unsigned(3779, 12), 1579 => to_unsigned(112, 12), 1580 => to_unsigned(2998, 12), 1581 => to_unsigned(763, 12), 1582 => to_unsigned(1648, 12), 1583 => to_unsigned(610, 12), 1584 => to_unsigned(2630, 12), 1585 => to_unsigned(2824, 12), 1586 => to_unsigned(3456, 12), 1587 => to_unsigned(919, 12), 1588 => to_unsigned(24, 12), 1589 => to_unsigned(2014, 12), 1590 => to_unsigned(3175, 12), 1591 => to_unsigned(1754, 12), 1592 => to_unsigned(2650, 12), 1593 => to_unsigned(3109, 12), 1594 => to_unsigned(3116, 12), 1595 => to_unsigned(1867, 12), 1596 => to_unsigned(142, 12), 1597 => to_unsigned(701, 12), 1598 => to_unsigned(1567, 12), 1599 => to_unsigned(3181, 12), 1600 => to_unsigned(1801, 12), 1601 => to_unsigned(2032, 12), 1602 => to_unsigned(2190, 12), 1603 => to_unsigned(3306, 12), 1604 => to_unsigned(2250, 12), 1605 => to_unsigned(3787, 12), 1606 => to_unsigned(927, 12), 1607 => to_unsigned(1821, 12), 1608 => to_unsigned(3506, 12), 1609 => to_unsigned(2061, 12), 1610 => to_unsigned(3859, 12), 1611 => to_unsigned(608, 12), 1612 => to_unsigned(3699, 12), 1613 => to_unsigned(2992, 12), 1614 => to_unsigned(414, 12), 1615 => to_unsigned(613, 12), 1616 => to_unsigned(2264, 12), 1617 => to_unsigned(2686, 12), 1618 => to_unsigned(3471, 12), 1619 => to_unsigned(1064, 12), 1620 => to_unsigned(2315, 12), 1621 => to_unsigned(2532, 12), 1622 => to_unsigned(639, 12), 1623 => to_unsigned(75, 12), 1624 => to_unsigned(73, 12), 1625 => to_unsigned(1472, 12), 1626 => to_unsigned(2905, 12), 1627 => to_unsigned(2257, 12), 1628 => to_unsigned(576, 12), 1629 => to_unsigned(2215, 12), 1630 => to_unsigned(1910, 12), 1631 => to_unsigned(3130, 12), 1632 => to_unsigned(1647, 12), 1633 => to_unsigned(1735, 12), 1634 => to_unsigned(1071, 12), 1635 => to_unsigned(1669, 12), 1636 => to_unsigned(1988, 12), 1637 => to_unsigned(4008, 12), 1638 => to_unsigned(2520, 12), 1639 => to_unsigned(2074, 12), 1640 => to_unsigned(3054, 12), 1641 => to_unsigned(1234, 12), 1642 => to_unsigned(105, 12), 1643 => to_unsigned(588, 12), 1644 => to_unsigned(1225, 12), 1645 => to_unsigned(3986, 12), 1646 => to_unsigned(2825, 12), 1647 => to_unsigned(4068, 12), 1648 => to_unsigned(1977, 12), 1649 => to_unsigned(2049, 12), 1650 => to_unsigned(2743, 12), 1651 => to_unsigned(1582, 12), 1652 => to_unsigned(59, 12), 1653 => to_unsigned(2731, 12), 1654 => to_unsigned(568, 12), 1655 => to_unsigned(308, 12), 1656 => to_unsigned(837, 12), 1657 => to_unsigned(3227, 12), 1658 => to_unsigned(2717, 12), 1659 => to_unsigned(298, 12), 1660 => to_unsigned(2008, 12), 1661 => to_unsigned(636, 12), 1662 => to_unsigned(1305, 12), 1663 => to_unsigned(365, 12), 1664 => to_unsigned(3381, 12), 1665 => to_unsigned(754, 12), 1666 => to_unsigned(1903, 12), 1667 => to_unsigned(2642, 12), 1668 => to_unsigned(2853, 12), 1669 => to_unsigned(1812, 12), 1670 => to_unsigned(3550, 12), 1671 => to_unsigned(3511, 12), 1672 => to_unsigned(1729, 12), 1673 => to_unsigned(1294, 12), 1674 => to_unsigned(2974, 12), 1675 => to_unsigned(1370, 12), 1676 => to_unsigned(1511, 12), 1677 => to_unsigned(104, 12), 1678 => to_unsigned(68, 12), 1679 => to_unsigned(696, 12), 1680 => to_unsigned(2965, 12), 1681 => to_unsigned(1120, 12), 1682 => to_unsigned(3831, 12), 1683 => to_unsigned(2501, 12), 1684 => to_unsigned(701, 12), 1685 => to_unsigned(4018, 12), 1686 => to_unsigned(1568, 12), 1687 => to_unsigned(1970, 12), 1688 => to_unsigned(1985, 12), 1689 => to_unsigned(417, 12), 1690 => to_unsigned(1470, 12), 1691 => to_unsigned(3353, 12), 1692 => to_unsigned(2802, 12), 1693 => to_unsigned(3773, 12), 1694 => to_unsigned(1633, 12), 1695 => to_unsigned(1429, 12), 1696 => to_unsigned(997, 12), 1697 => to_unsigned(950, 12), 1698 => to_unsigned(1916, 12), 1699 => to_unsigned(1577, 12), 1700 => to_unsigned(3874, 12), 1701 => to_unsigned(1427, 12), 1702 => to_unsigned(4072, 12), 1703 => to_unsigned(3298, 12), 1704 => to_unsigned(1966, 12), 1705 => to_unsigned(2203, 12), 1706 => to_unsigned(3980, 12), 1707 => to_unsigned(242, 12), 1708 => to_unsigned(2084, 12), 1709 => to_unsigned(2117, 12), 1710 => to_unsigned(163, 12), 1711 => to_unsigned(3333, 12), 1712 => to_unsigned(3042, 12), 1713 => to_unsigned(2078, 12), 1714 => to_unsigned(2369, 12), 1715 => to_unsigned(992, 12), 1716 => to_unsigned(1155, 12), 1717 => to_unsigned(1586, 12), 1718 => to_unsigned(950, 12), 1719 => to_unsigned(966, 12), 1720 => to_unsigned(983, 12), 1721 => to_unsigned(3745, 12), 1722 => to_unsigned(1707, 12), 1723 => to_unsigned(2065, 12), 1724 => to_unsigned(1844, 12), 1725 => to_unsigned(470, 12), 1726 => to_unsigned(2205, 12), 1727 => to_unsigned(377, 12), 1728 => to_unsigned(346, 12), 1729 => to_unsigned(3275, 12), 1730 => to_unsigned(751, 12), 1731 => to_unsigned(599, 12), 1732 => to_unsigned(3516, 12), 1733 => to_unsigned(488, 12), 1734 => to_unsigned(3498, 12), 1735 => to_unsigned(480, 12), 1736 => to_unsigned(1524, 12), 1737 => to_unsigned(450, 12), 1738 => to_unsigned(1401, 12), 1739 => to_unsigned(3150, 12), 1740 => to_unsigned(2317, 12), 1741 => to_unsigned(2479, 12), 1742 => to_unsigned(1422, 12), 1743 => to_unsigned(451, 12), 1744 => to_unsigned(878, 12), 1745 => to_unsigned(1579, 12), 1746 => to_unsigned(3707, 12), 1747 => to_unsigned(399, 12), 1748 => to_unsigned(2388, 12), 1749 => to_unsigned(1041, 12), 1750 => to_unsigned(1669, 12), 1751 => to_unsigned(807, 12), 1752 => to_unsigned(1968, 12), 1753 => to_unsigned(1389, 12), 1754 => to_unsigned(3009, 12), 1755 => to_unsigned(3729, 12), 1756 => to_unsigned(1488, 12), 1757 => to_unsigned(2309, 12), 1758 => to_unsigned(1194, 12), 1759 => to_unsigned(2890, 12), 1760 => to_unsigned(3163, 12), 1761 => to_unsigned(2582, 12), 1762 => to_unsigned(362, 12), 1763 => to_unsigned(1455, 12), 1764 => to_unsigned(2895, 12), 1765 => to_unsigned(2959, 12), 1766 => to_unsigned(2701, 12), 1767 => to_unsigned(1157, 12), 1768 => to_unsigned(2841, 12), 1769 => to_unsigned(2956, 12), 1770 => to_unsigned(660, 12), 1771 => to_unsigned(1744, 12), 1772 => to_unsigned(1307, 12), 1773 => to_unsigned(894, 12), 1774 => to_unsigned(2076, 12), 1775 => to_unsigned(1985, 12), 1776 => to_unsigned(859, 12), 1777 => to_unsigned(790, 12), 1778 => to_unsigned(624, 12), 1779 => to_unsigned(1265, 12), 1780 => to_unsigned(3226, 12), 1781 => to_unsigned(1200, 12), 1782 => to_unsigned(1962, 12), 1783 => to_unsigned(1795, 12), 1784 => to_unsigned(1685, 12), 1785 => to_unsigned(3665, 12), 1786 => to_unsigned(3443, 12), 1787 => to_unsigned(767, 12), 1788 => to_unsigned(221, 12), 1789 => to_unsigned(1344, 12), 1790 => to_unsigned(3588, 12), 1791 => to_unsigned(2791, 12), 1792 => to_unsigned(600, 12), 1793 => to_unsigned(3564, 12), 1794 => to_unsigned(3551, 12), 1795 => to_unsigned(547, 12), 1796 => to_unsigned(573, 12), 1797 => to_unsigned(3185, 12), 1798 => to_unsigned(694, 12), 1799 => to_unsigned(3522, 12), 1800 => to_unsigned(2137, 12), 1801 => to_unsigned(670, 12), 1802 => to_unsigned(2001, 12), 1803 => to_unsigned(2736, 12), 1804 => to_unsigned(264, 12), 1805 => to_unsigned(144, 12), 1806 => to_unsigned(3192, 12), 1807 => to_unsigned(2206, 12), 1808 => to_unsigned(3267, 12), 1809 => to_unsigned(1390, 12), 1810 => to_unsigned(3863, 12), 1811 => to_unsigned(3680, 12), 1812 => to_unsigned(3119, 12), 1813 => to_unsigned(267, 12), 1814 => to_unsigned(1325, 12), 1815 => to_unsigned(91, 12), 1816 => to_unsigned(3236, 12), 1817 => to_unsigned(1279, 12), 1818 => to_unsigned(2332, 12), 1819 => to_unsigned(1833, 12), 1820 => to_unsigned(1755, 12), 1821 => to_unsigned(775, 12), 1822 => to_unsigned(1980, 12), 1823 => to_unsigned(3893, 12), 1824 => to_unsigned(1400, 12), 1825 => to_unsigned(1645, 12), 1826 => to_unsigned(2168, 12), 1827 => to_unsigned(991, 12), 1828 => to_unsigned(82, 12), 1829 => to_unsigned(1441, 12), 1830 => to_unsigned(1966, 12), 1831 => to_unsigned(3857, 12), 1832 => to_unsigned(3052, 12), 1833 => to_unsigned(3973, 12), 1834 => to_unsigned(3421, 12), 1835 => to_unsigned(1382, 12), 1836 => to_unsigned(3113, 12), 1837 => to_unsigned(3514, 12), 1838 => to_unsigned(1483, 12), 1839 => to_unsigned(1637, 12), 1840 => to_unsigned(3816, 12), 1841 => to_unsigned(3976, 12), 1842 => to_unsigned(3948, 12), 1843 => to_unsigned(1508, 12), 1844 => to_unsigned(474, 12), 1845 => to_unsigned(985, 12), 1846 => to_unsigned(1692, 12), 1847 => to_unsigned(858, 12), 1848 => to_unsigned(1822, 12), 1849 => to_unsigned(730, 12), 1850 => to_unsigned(3954, 12), 1851 => to_unsigned(1408, 12), 1852 => to_unsigned(2600, 12), 1853 => to_unsigned(1145, 12), 1854 => to_unsigned(1049, 12), 1855 => to_unsigned(2727, 12), 1856 => to_unsigned(3718, 12), 1857 => to_unsigned(643, 12), 1858 => to_unsigned(556, 12), 1859 => to_unsigned(587, 12), 1860 => to_unsigned(1702, 12), 1861 => to_unsigned(3242, 12), 1862 => to_unsigned(2549, 12), 1863 => to_unsigned(582, 12), 1864 => to_unsigned(3424, 12), 1865 => to_unsigned(1086, 12), 1866 => to_unsigned(2262, 12), 1867 => to_unsigned(2455, 12), 1868 => to_unsigned(3844, 12), 1869 => to_unsigned(3138, 12), 1870 => to_unsigned(940, 12), 1871 => to_unsigned(871, 12), 1872 => to_unsigned(185, 12), 1873 => to_unsigned(1343, 12), 1874 => to_unsigned(2510, 12), 1875 => to_unsigned(795, 12), 1876 => to_unsigned(3713, 12), 1877 => to_unsigned(2157, 12), 1878 => to_unsigned(1871, 12), 1879 => to_unsigned(2350, 12), 1880 => to_unsigned(1463, 12), 1881 => to_unsigned(2031, 12), 1882 => to_unsigned(3860, 12), 1883 => to_unsigned(2952, 12), 1884 => to_unsigned(3176, 12), 1885 => to_unsigned(3707, 12), 1886 => to_unsigned(1296, 12), 1887 => to_unsigned(1685, 12), 1888 => to_unsigned(2422, 12), 1889 => to_unsigned(1058, 12), 1890 => to_unsigned(805, 12), 1891 => to_unsigned(3032, 12), 1892 => to_unsigned(3971, 12), 1893 => to_unsigned(214, 12), 1894 => to_unsigned(3967, 12), 1895 => to_unsigned(2914, 12), 1896 => to_unsigned(3406, 12), 1897 => to_unsigned(1515, 12), 1898 => to_unsigned(267, 12), 1899 => to_unsigned(1408, 12), 1900 => to_unsigned(925, 12), 1901 => to_unsigned(3316, 12), 1902 => to_unsigned(3277, 12), 1903 => to_unsigned(1971, 12), 1904 => to_unsigned(1302, 12), 1905 => to_unsigned(358, 12), 1906 => to_unsigned(666, 12), 1907 => to_unsigned(2938, 12), 1908 => to_unsigned(3893, 12), 1909 => to_unsigned(1138, 12), 1910 => to_unsigned(3485, 12), 1911 => to_unsigned(1703, 12), 1912 => to_unsigned(1207, 12), 1913 => to_unsigned(1138, 12), 1914 => to_unsigned(1543, 12), 1915 => to_unsigned(2755, 12), 1916 => to_unsigned(1964, 12), 1917 => to_unsigned(2516, 12), 1918 => to_unsigned(2399, 12), 1919 => to_unsigned(2287, 12), 1920 => to_unsigned(1031, 12), 1921 => to_unsigned(2936, 12), 1922 => to_unsigned(1230, 12), 1923 => to_unsigned(2061, 12), 1924 => to_unsigned(3689, 12), 1925 => to_unsigned(734, 12), 1926 => to_unsigned(1521, 12), 1927 => to_unsigned(1858, 12), 1928 => to_unsigned(3961, 12), 1929 => to_unsigned(2426, 12), 1930 => to_unsigned(2310, 12), 1931 => to_unsigned(2267, 12), 1932 => to_unsigned(519, 12), 1933 => to_unsigned(745, 12), 1934 => to_unsigned(133, 12), 1935 => to_unsigned(3427, 12), 1936 => to_unsigned(44, 12), 1937 => to_unsigned(3686, 12), 1938 => to_unsigned(971, 12), 1939 => to_unsigned(501, 12), 1940 => to_unsigned(1956, 12), 1941 => to_unsigned(2721, 12), 1942 => to_unsigned(1899, 12), 1943 => to_unsigned(2485, 12), 1944 => to_unsigned(2906, 12), 1945 => to_unsigned(1817, 12), 1946 => to_unsigned(908, 12), 1947 => to_unsigned(2012, 12), 1948 => to_unsigned(951, 12), 1949 => to_unsigned(3528, 12), 1950 => to_unsigned(2604, 12), 1951 => to_unsigned(2891, 12), 1952 => to_unsigned(3050, 12), 1953 => to_unsigned(513, 12), 1954 => to_unsigned(1852, 12), 1955 => to_unsigned(1706, 12), 1956 => to_unsigned(1461, 12), 1957 => to_unsigned(2578, 12), 1958 => to_unsigned(2371, 12), 1959 => to_unsigned(1154, 12), 1960 => to_unsigned(2041, 12), 1961 => to_unsigned(3110, 12), 1962 => to_unsigned(1928, 12), 1963 => to_unsigned(470, 12), 1964 => to_unsigned(3683, 12), 1965 => to_unsigned(3268, 12), 1966 => to_unsigned(2730, 12), 1967 => to_unsigned(1231, 12), 1968 => to_unsigned(3998, 12), 1969 => to_unsigned(2833, 12), 1970 => to_unsigned(702, 12), 1971 => to_unsigned(1381, 12), 1972 => to_unsigned(3268, 12), 1973 => to_unsigned(790, 12), 1974 => to_unsigned(1651, 12), 1975 => to_unsigned(3502, 12), 1976 => to_unsigned(3826, 12), 1977 => to_unsigned(1158, 12), 1978 => to_unsigned(1689, 12), 1979 => to_unsigned(982, 12), 1980 => to_unsigned(1651, 12), 1981 => to_unsigned(3256, 12), 1982 => to_unsigned(3683, 12), 1983 => to_unsigned(3900, 12), 1984 => to_unsigned(3013, 12), 1985 => to_unsigned(2236, 12), 1986 => to_unsigned(298, 12), 1987 => to_unsigned(986, 12), 1988 => to_unsigned(1286, 12), 1989 => to_unsigned(3556, 12), 1990 => to_unsigned(3114, 12), 1991 => to_unsigned(3363, 12), 1992 => to_unsigned(2740, 12), 1993 => to_unsigned(3608, 12), 1994 => to_unsigned(3600, 12), 1995 => to_unsigned(1871, 12), 1996 => to_unsigned(2899, 12), 1997 => to_unsigned(2717, 12), 1998 => to_unsigned(2241, 12), 1999 => to_unsigned(3486, 12), 2000 => to_unsigned(324, 12), 2001 => to_unsigned(4074, 12), 2002 => to_unsigned(3705, 12), 2003 => to_unsigned(2360, 12), 2004 => to_unsigned(2144, 12), 2005 => to_unsigned(2744, 12), 2006 => to_unsigned(2579, 12), 2007 => to_unsigned(2136, 12), 2008 => to_unsigned(1008, 12), 2009 => to_unsigned(3513, 12), 2010 => to_unsigned(1714, 12), 2011 => to_unsigned(755, 12), 2012 => to_unsigned(370, 12), 2013 => to_unsigned(1459, 12), 2014 => to_unsigned(1771, 12), 2015 => to_unsigned(2, 12), 2016 => to_unsigned(173, 12), 2017 => to_unsigned(285, 12), 2018 => to_unsigned(2829, 12), 2019 => to_unsigned(2818, 12), 2020 => to_unsigned(300, 12), 2021 => to_unsigned(112, 12), 2022 => to_unsigned(1409, 12), 2023 => to_unsigned(2736, 12), 2024 => to_unsigned(3727, 12), 2025 => to_unsigned(3140, 12), 2026 => to_unsigned(2275, 12), 2027 => to_unsigned(50, 12), 2028 => to_unsigned(3663, 12), 2029 => to_unsigned(2750, 12), 2030 => to_unsigned(3990, 12), 2031 => to_unsigned(148, 12), 2032 => to_unsigned(3553, 12), 2033 => to_unsigned(2594, 12), 2034 => to_unsigned(3266, 12), 2035 => to_unsigned(799, 12), 2036 => to_unsigned(638, 12), 2037 => to_unsigned(2435, 12), 2038 => to_unsigned(2309, 12), 2039 => to_unsigned(2261, 12), 2040 => to_unsigned(3693, 12), 2041 => to_unsigned(575, 12), 2042 => to_unsigned(3967, 12), 2043 => to_unsigned(1708, 12), 2044 => to_unsigned(1834, 12), 2045 => to_unsigned(1675, 12), 2046 => to_unsigned(3329, 12), 2047 => to_unsigned(595, 12)),
            9 => (0 => to_unsigned(1621, 12), 1 => to_unsigned(1898, 12), 2 => to_unsigned(3608, 12), 3 => to_unsigned(3857, 12), 4 => to_unsigned(3815, 12), 5 => to_unsigned(1507, 12), 6 => to_unsigned(4082, 12), 7 => to_unsigned(2091, 12), 8 => to_unsigned(2296, 12), 9 => to_unsigned(2572, 12), 10 => to_unsigned(1275, 12), 11 => to_unsigned(429, 12), 12 => to_unsigned(1453, 12), 13 => to_unsigned(3263, 12), 14 => to_unsigned(2945, 12), 15 => to_unsigned(3673, 12), 16 => to_unsigned(1532, 12), 17 => to_unsigned(1114, 12), 18 => to_unsigned(2015, 12), 19 => to_unsigned(2664, 12), 20 => to_unsigned(831, 12), 21 => to_unsigned(2944, 12), 22 => to_unsigned(3210, 12), 23 => to_unsigned(3761, 12), 24 => to_unsigned(679, 12), 25 => to_unsigned(3221, 12), 26 => to_unsigned(3020, 12), 27 => to_unsigned(1583, 12), 28 => to_unsigned(2146, 12), 29 => to_unsigned(396, 12), 30 => to_unsigned(2295, 12), 31 => to_unsigned(1707, 12), 32 => to_unsigned(3495, 12), 33 => to_unsigned(3411, 12), 34 => to_unsigned(1070, 12), 35 => to_unsigned(3630, 12), 36 => to_unsigned(2022, 12), 37 => to_unsigned(1336, 12), 38 => to_unsigned(833, 12), 39 => to_unsigned(3652, 12), 40 => to_unsigned(1456, 12), 41 => to_unsigned(3170, 12), 42 => to_unsigned(3682, 12), 43 => to_unsigned(1880, 12), 44 => to_unsigned(680, 12), 45 => to_unsigned(2388, 12), 46 => to_unsigned(648, 12), 47 => to_unsigned(1054, 12), 48 => to_unsigned(2963, 12), 49 => to_unsigned(1052, 12), 50 => to_unsigned(3431, 12), 51 => to_unsigned(3373, 12), 52 => to_unsigned(3670, 12), 53 => to_unsigned(392, 12), 54 => to_unsigned(1934, 12), 55 => to_unsigned(3849, 12), 56 => to_unsigned(767, 12), 57 => to_unsigned(2285, 12), 58 => to_unsigned(2326, 12), 59 => to_unsigned(309, 12), 60 => to_unsigned(949, 12), 61 => to_unsigned(2446, 12), 62 => to_unsigned(3983, 12), 63 => to_unsigned(2866, 12), 64 => to_unsigned(4091, 12), 65 => to_unsigned(1840, 12), 66 => to_unsigned(579, 12), 67 => to_unsigned(1090, 12), 68 => to_unsigned(2694, 12), 69 => to_unsigned(3230, 12), 70 => to_unsigned(3361, 12), 71 => to_unsigned(886, 12), 72 => to_unsigned(3869, 12), 73 => to_unsigned(880, 12), 74 => to_unsigned(1267, 12), 75 => to_unsigned(3668, 12), 76 => to_unsigned(2379, 12), 77 => to_unsigned(2139, 12), 78 => to_unsigned(1396, 12), 79 => to_unsigned(3688, 12), 80 => to_unsigned(576, 12), 81 => to_unsigned(3624, 12), 82 => to_unsigned(3930, 12), 83 => to_unsigned(2519, 12), 84 => to_unsigned(932, 12), 85 => to_unsigned(2905, 12), 86 => to_unsigned(3165, 12), 87 => to_unsigned(2135, 12), 88 => to_unsigned(700, 12), 89 => to_unsigned(3014, 12), 90 => to_unsigned(1564, 12), 91 => to_unsigned(228, 12), 92 => to_unsigned(3707, 12), 93 => to_unsigned(138, 12), 94 => to_unsigned(796, 12), 95 => to_unsigned(2691, 12), 96 => to_unsigned(2228, 12), 97 => to_unsigned(602, 12), 98 => to_unsigned(3839, 12), 99 => to_unsigned(1819, 12), 100 => to_unsigned(2679, 12), 101 => to_unsigned(2774, 12), 102 => to_unsigned(725, 12), 103 => to_unsigned(2457, 12), 104 => to_unsigned(3201, 12), 105 => to_unsigned(3838, 12), 106 => to_unsigned(3951, 12), 107 => to_unsigned(58, 12), 108 => to_unsigned(1572, 12), 109 => to_unsigned(3008, 12), 110 => to_unsigned(2269, 12), 111 => to_unsigned(2045, 12), 112 => to_unsigned(223, 12), 113 => to_unsigned(1644, 12), 114 => to_unsigned(3350, 12), 115 => to_unsigned(1261, 12), 116 => to_unsigned(1739, 12), 117 => to_unsigned(641, 12), 118 => to_unsigned(1333, 12), 119 => to_unsigned(256, 12), 120 => to_unsigned(3599, 12), 121 => to_unsigned(69, 12), 122 => to_unsigned(1835, 12), 123 => to_unsigned(3232, 12), 124 => to_unsigned(2167, 12), 125 => to_unsigned(484, 12), 126 => to_unsigned(4093, 12), 127 => to_unsigned(3802, 12), 128 => to_unsigned(528, 12), 129 => to_unsigned(2840, 12), 130 => to_unsigned(546, 12), 131 => to_unsigned(3965, 12), 132 => to_unsigned(2024, 12), 133 => to_unsigned(3652, 12), 134 => to_unsigned(1853, 12), 135 => to_unsigned(600, 12), 136 => to_unsigned(3953, 12), 137 => to_unsigned(2484, 12), 138 => to_unsigned(3523, 12), 139 => to_unsigned(3591, 12), 140 => to_unsigned(1271, 12), 141 => to_unsigned(2777, 12), 142 => to_unsigned(3744, 12), 143 => to_unsigned(2228, 12), 144 => to_unsigned(3106, 12), 145 => to_unsigned(3545, 12), 146 => to_unsigned(3150, 12), 147 => to_unsigned(2316, 12), 148 => to_unsigned(1667, 12), 149 => to_unsigned(1742, 12), 150 => to_unsigned(1727, 12), 151 => to_unsigned(3117, 12), 152 => to_unsigned(3825, 12), 153 => to_unsigned(1277, 12), 154 => to_unsigned(329, 12), 155 => to_unsigned(502, 12), 156 => to_unsigned(3851, 12), 157 => to_unsigned(569, 12), 158 => to_unsigned(3743, 12), 159 => to_unsigned(3842, 12), 160 => to_unsigned(2903, 12), 161 => to_unsigned(842, 12), 162 => to_unsigned(1623, 12), 163 => to_unsigned(655, 12), 164 => to_unsigned(1684, 12), 165 => to_unsigned(200, 12), 166 => to_unsigned(823, 12), 167 => to_unsigned(7, 12), 168 => to_unsigned(642, 12), 169 => to_unsigned(486, 12), 170 => to_unsigned(3821, 12), 171 => to_unsigned(1950, 12), 172 => to_unsigned(563, 12), 173 => to_unsigned(1265, 12), 174 => to_unsigned(628, 12), 175 => to_unsigned(2894, 12), 176 => to_unsigned(2812, 12), 177 => to_unsigned(289, 12), 178 => to_unsigned(112, 12), 179 => to_unsigned(3850, 12), 180 => to_unsigned(283, 12), 181 => to_unsigned(2272, 12), 182 => to_unsigned(921, 12), 183 => to_unsigned(868, 12), 184 => to_unsigned(2335, 12), 185 => to_unsigned(3811, 12), 186 => to_unsigned(3187, 12), 187 => to_unsigned(1678, 12), 188 => to_unsigned(2292, 12), 189 => to_unsigned(1546, 12), 190 => to_unsigned(1880, 12), 191 => to_unsigned(1636, 12), 192 => to_unsigned(1501, 12), 193 => to_unsigned(7, 12), 194 => to_unsigned(2481, 12), 195 => to_unsigned(3167, 12), 196 => to_unsigned(1395, 12), 197 => to_unsigned(3408, 12), 198 => to_unsigned(2685, 12), 199 => to_unsigned(339, 12), 200 => to_unsigned(3336, 12), 201 => to_unsigned(614, 12), 202 => to_unsigned(371, 12), 203 => to_unsigned(3367, 12), 204 => to_unsigned(998, 12), 205 => to_unsigned(1196, 12), 206 => to_unsigned(3302, 12), 207 => to_unsigned(2160, 12), 208 => to_unsigned(378, 12), 209 => to_unsigned(623, 12), 210 => to_unsigned(2049, 12), 211 => to_unsigned(409, 12), 212 => to_unsigned(64, 12), 213 => to_unsigned(85, 12), 214 => to_unsigned(3244, 12), 215 => to_unsigned(2825, 12), 216 => to_unsigned(114, 12), 217 => to_unsigned(1120, 12), 218 => to_unsigned(2798, 12), 219 => to_unsigned(985, 12), 220 => to_unsigned(1667, 12), 221 => to_unsigned(3953, 12), 222 => to_unsigned(1546, 12), 223 => to_unsigned(1356, 12), 224 => to_unsigned(1098, 12), 225 => to_unsigned(2661, 12), 226 => to_unsigned(2478, 12), 227 => to_unsigned(3372, 12), 228 => to_unsigned(2608, 12), 229 => to_unsigned(2683, 12), 230 => to_unsigned(2127, 12), 231 => to_unsigned(150, 12), 232 => to_unsigned(1513, 12), 233 => to_unsigned(3208, 12), 234 => to_unsigned(3044, 12), 235 => to_unsigned(2024, 12), 236 => to_unsigned(1080, 12), 237 => to_unsigned(362, 12), 238 => to_unsigned(1729, 12), 239 => to_unsigned(3557, 12), 240 => to_unsigned(1202, 12), 241 => to_unsigned(660, 12), 242 => to_unsigned(24, 12), 243 => to_unsigned(1652, 12), 244 => to_unsigned(3033, 12), 245 => to_unsigned(1985, 12), 246 => to_unsigned(2119, 12), 247 => to_unsigned(2128, 12), 248 => to_unsigned(2240, 12), 249 => to_unsigned(1780, 12), 250 => to_unsigned(2184, 12), 251 => to_unsigned(2898, 12), 252 => to_unsigned(1572, 12), 253 => to_unsigned(2582, 12), 254 => to_unsigned(3302, 12), 255 => to_unsigned(2550, 12), 256 => to_unsigned(2130, 12), 257 => to_unsigned(2365, 12), 258 => to_unsigned(564, 12), 259 => to_unsigned(630, 12), 260 => to_unsigned(1370, 12), 261 => to_unsigned(565, 12), 262 => to_unsigned(2954, 12), 263 => to_unsigned(3594, 12), 264 => to_unsigned(1972, 12), 265 => to_unsigned(3387, 12), 266 => to_unsigned(111, 12), 267 => to_unsigned(2860, 12), 268 => to_unsigned(3888, 12), 269 => to_unsigned(2387, 12), 270 => to_unsigned(1786, 12), 271 => to_unsigned(1450, 12), 272 => to_unsigned(528, 12), 273 => to_unsigned(2279, 12), 274 => to_unsigned(381, 12), 275 => to_unsigned(3630, 12), 276 => to_unsigned(1572, 12), 277 => to_unsigned(1518, 12), 278 => to_unsigned(460, 12), 279 => to_unsigned(219, 12), 280 => to_unsigned(1891, 12), 281 => to_unsigned(3088, 12), 282 => to_unsigned(2439, 12), 283 => to_unsigned(1161, 12), 284 => to_unsigned(746, 12), 285 => to_unsigned(825, 12), 286 => to_unsigned(3781, 12), 287 => to_unsigned(2310, 12), 288 => to_unsigned(547, 12), 289 => to_unsigned(624, 12), 290 => to_unsigned(2704, 12), 291 => to_unsigned(583, 12), 292 => to_unsigned(1886, 12), 293 => to_unsigned(3693, 12), 294 => to_unsigned(2368, 12), 295 => to_unsigned(3639, 12), 296 => to_unsigned(1479, 12), 297 => to_unsigned(771, 12), 298 => to_unsigned(2095, 12), 299 => to_unsigned(899, 12), 300 => to_unsigned(2200, 12), 301 => to_unsigned(3585, 12), 302 => to_unsigned(1157, 12), 303 => to_unsigned(676, 12), 304 => to_unsigned(2710, 12), 305 => to_unsigned(2265, 12), 306 => to_unsigned(2693, 12), 307 => to_unsigned(821, 12), 308 => to_unsigned(910, 12), 309 => to_unsigned(1151, 12), 310 => to_unsigned(2255, 12), 311 => to_unsigned(2213, 12), 312 => to_unsigned(1586, 12), 313 => to_unsigned(1346, 12), 314 => to_unsigned(3037, 12), 315 => to_unsigned(819, 12), 316 => to_unsigned(186, 12), 317 => to_unsigned(2370, 12), 318 => to_unsigned(3143, 12), 319 => to_unsigned(3967, 12), 320 => to_unsigned(3655, 12), 321 => to_unsigned(3984, 12), 322 => to_unsigned(1044, 12), 323 => to_unsigned(4071, 12), 324 => to_unsigned(1618, 12), 325 => to_unsigned(685, 12), 326 => to_unsigned(1385, 12), 327 => to_unsigned(2038, 12), 328 => to_unsigned(3674, 12), 329 => to_unsigned(3430, 12), 330 => to_unsigned(1306, 12), 331 => to_unsigned(3278, 12), 332 => to_unsigned(346, 12), 333 => to_unsigned(3324, 12), 334 => to_unsigned(2532, 12), 335 => to_unsigned(1793, 12), 336 => to_unsigned(588, 12), 337 => to_unsigned(266, 12), 338 => to_unsigned(1681, 12), 339 => to_unsigned(2061, 12), 340 => to_unsigned(2959, 12), 341 => to_unsigned(3249, 12), 342 => to_unsigned(3790, 12), 343 => to_unsigned(2851, 12), 344 => to_unsigned(130, 12), 345 => to_unsigned(468, 12), 346 => to_unsigned(1805, 12), 347 => to_unsigned(2791, 12), 348 => to_unsigned(2696, 12), 349 => to_unsigned(3087, 12), 350 => to_unsigned(3604, 12), 351 => to_unsigned(4095, 12), 352 => to_unsigned(2196, 12), 353 => to_unsigned(2962, 12), 354 => to_unsigned(519, 12), 355 => to_unsigned(3038, 12), 356 => to_unsigned(603, 12), 357 => to_unsigned(1272, 12), 358 => to_unsigned(1227, 12), 359 => to_unsigned(2562, 12), 360 => to_unsigned(1664, 12), 361 => to_unsigned(1327, 12), 362 => to_unsigned(3008, 12), 363 => to_unsigned(3933, 12), 364 => to_unsigned(2346, 12), 365 => to_unsigned(2038, 12), 366 => to_unsigned(4082, 12), 367 => to_unsigned(2531, 12), 368 => to_unsigned(1706, 12), 369 => to_unsigned(3612, 12), 370 => to_unsigned(3066, 12), 371 => to_unsigned(82, 12), 372 => to_unsigned(677, 12), 373 => to_unsigned(2057, 12), 374 => to_unsigned(393, 12), 375 => to_unsigned(1696, 12), 376 => to_unsigned(237, 12), 377 => to_unsigned(3999, 12), 378 => to_unsigned(2103, 12), 379 => to_unsigned(1272, 12), 380 => to_unsigned(3014, 12), 381 => to_unsigned(2127, 12), 382 => to_unsigned(981, 12), 383 => to_unsigned(2277, 12), 384 => to_unsigned(348, 12), 385 => to_unsigned(1579, 12), 386 => to_unsigned(1978, 12), 387 => to_unsigned(2756, 12), 388 => to_unsigned(838, 12), 389 => to_unsigned(3006, 12), 390 => to_unsigned(3318, 12), 391 => to_unsigned(1375, 12), 392 => to_unsigned(3014, 12), 393 => to_unsigned(575, 12), 394 => to_unsigned(1642, 12), 395 => to_unsigned(1124, 12), 396 => to_unsigned(2159, 12), 397 => to_unsigned(2024, 12), 398 => to_unsigned(112, 12), 399 => to_unsigned(2290, 12), 400 => to_unsigned(3995, 12), 401 => to_unsigned(360, 12), 402 => to_unsigned(1339, 12), 403 => to_unsigned(943, 12), 404 => to_unsigned(1879, 12), 405 => to_unsigned(2651, 12), 406 => to_unsigned(1434, 12), 407 => to_unsigned(1437, 12), 408 => to_unsigned(3329, 12), 409 => to_unsigned(2765, 12), 410 => to_unsigned(2726, 12), 411 => to_unsigned(3791, 12), 412 => to_unsigned(3322, 12), 413 => to_unsigned(1884, 12), 414 => to_unsigned(3559, 12), 415 => to_unsigned(1245, 12), 416 => to_unsigned(2467, 12), 417 => to_unsigned(3532, 12), 418 => to_unsigned(1688, 12), 419 => to_unsigned(289, 12), 420 => to_unsigned(2927, 12), 421 => to_unsigned(2282, 12), 422 => to_unsigned(898, 12), 423 => to_unsigned(3688, 12), 424 => to_unsigned(3390, 12), 425 => to_unsigned(1901, 12), 426 => to_unsigned(63, 12), 427 => to_unsigned(693, 12), 428 => to_unsigned(2480, 12), 429 => to_unsigned(2988, 12), 430 => to_unsigned(165, 12), 431 => to_unsigned(3088, 12), 432 => to_unsigned(295, 12), 433 => to_unsigned(3408, 12), 434 => to_unsigned(3758, 12), 435 => to_unsigned(1850, 12), 436 => to_unsigned(1316, 12), 437 => to_unsigned(1793, 12), 438 => to_unsigned(93, 12), 439 => to_unsigned(85, 12), 440 => to_unsigned(461, 12), 441 => to_unsigned(1345, 12), 442 => to_unsigned(1184, 12), 443 => to_unsigned(3872, 12), 444 => to_unsigned(2314, 12), 445 => to_unsigned(3230, 12), 446 => to_unsigned(447, 12), 447 => to_unsigned(3619, 12), 448 => to_unsigned(3406, 12), 449 => to_unsigned(2259, 12), 450 => to_unsigned(386, 12), 451 => to_unsigned(547, 12), 452 => to_unsigned(3894, 12), 453 => to_unsigned(2608, 12), 454 => to_unsigned(2751, 12), 455 => to_unsigned(1961, 12), 456 => to_unsigned(2341, 12), 457 => to_unsigned(2462, 12), 458 => to_unsigned(161, 12), 459 => to_unsigned(525, 12), 460 => to_unsigned(2581, 12), 461 => to_unsigned(1653, 12), 462 => to_unsigned(414, 12), 463 => to_unsigned(3596, 12), 464 => to_unsigned(2483, 12), 465 => to_unsigned(3290, 12), 466 => to_unsigned(3151, 12), 467 => to_unsigned(3101, 12), 468 => to_unsigned(2119, 12), 469 => to_unsigned(2605, 12), 470 => to_unsigned(2287, 12), 471 => to_unsigned(719, 12), 472 => to_unsigned(1418, 12), 473 => to_unsigned(3944, 12), 474 => to_unsigned(1271, 12), 475 => to_unsigned(639, 12), 476 => to_unsigned(2200, 12), 477 => to_unsigned(1105, 12), 478 => to_unsigned(987, 12), 479 => to_unsigned(1195, 12), 480 => to_unsigned(323, 12), 481 => to_unsigned(268, 12), 482 => to_unsigned(2484, 12), 483 => to_unsigned(1194, 12), 484 => to_unsigned(3961, 12), 485 => to_unsigned(4049, 12), 486 => to_unsigned(2851, 12), 487 => to_unsigned(4003, 12), 488 => to_unsigned(1431, 12), 489 => to_unsigned(1138, 12), 490 => to_unsigned(4092, 12), 491 => to_unsigned(51, 12), 492 => to_unsigned(1912, 12), 493 => to_unsigned(2877, 12), 494 => to_unsigned(92, 12), 495 => to_unsigned(2884, 12), 496 => to_unsigned(2994, 12), 497 => to_unsigned(1903, 12), 498 => to_unsigned(422, 12), 499 => to_unsigned(2245, 12), 500 => to_unsigned(463, 12), 501 => to_unsigned(2446, 12), 502 => to_unsigned(2918, 12), 503 => to_unsigned(1079, 12), 504 => to_unsigned(2133, 12), 505 => to_unsigned(3532, 12), 506 => to_unsigned(3645, 12), 507 => to_unsigned(3755, 12), 508 => to_unsigned(4048, 12), 509 => to_unsigned(3432, 12), 510 => to_unsigned(1107, 12), 511 => to_unsigned(890, 12), 512 => to_unsigned(435, 12), 513 => to_unsigned(1816, 12), 514 => to_unsigned(4049, 12), 515 => to_unsigned(3891, 12), 516 => to_unsigned(1723, 12), 517 => to_unsigned(2731, 12), 518 => to_unsigned(201, 12), 519 => to_unsigned(2693, 12), 520 => to_unsigned(3058, 12), 521 => to_unsigned(3555, 12), 522 => to_unsigned(3865, 12), 523 => to_unsigned(3529, 12), 524 => to_unsigned(3780, 12), 525 => to_unsigned(3665, 12), 526 => to_unsigned(93, 12), 527 => to_unsigned(1226, 12), 528 => to_unsigned(981, 12), 529 => to_unsigned(2545, 12), 530 => to_unsigned(29, 12), 531 => to_unsigned(2344, 12), 532 => to_unsigned(185, 12), 533 => to_unsigned(665, 12), 534 => to_unsigned(1321, 12), 535 => to_unsigned(1604, 12), 536 => to_unsigned(1089, 12), 537 => to_unsigned(698, 12), 538 => to_unsigned(1702, 12), 539 => to_unsigned(1516, 12), 540 => to_unsigned(130, 12), 541 => to_unsigned(1504, 12), 542 => to_unsigned(434, 12), 543 => to_unsigned(2689, 12), 544 => to_unsigned(2934, 12), 545 => to_unsigned(3502, 12), 546 => to_unsigned(4086, 12), 547 => to_unsigned(3953, 12), 548 => to_unsigned(625, 12), 549 => to_unsigned(398, 12), 550 => to_unsigned(401, 12), 551 => to_unsigned(1858, 12), 552 => to_unsigned(131, 12), 553 => to_unsigned(1679, 12), 554 => to_unsigned(1991, 12), 555 => to_unsigned(3541, 12), 556 => to_unsigned(683, 12), 557 => to_unsigned(3143, 12), 558 => to_unsigned(1076, 12), 559 => to_unsigned(3473, 12), 560 => to_unsigned(539, 12), 561 => to_unsigned(2728, 12), 562 => to_unsigned(788, 12), 563 => to_unsigned(2239, 12), 564 => to_unsigned(2293, 12), 565 => to_unsigned(400, 12), 566 => to_unsigned(3697, 12), 567 => to_unsigned(491, 12), 568 => to_unsigned(1309, 12), 569 => to_unsigned(3689, 12), 570 => to_unsigned(2524, 12), 571 => to_unsigned(711, 12), 572 => to_unsigned(69, 12), 573 => to_unsigned(519, 12), 574 => to_unsigned(634, 12), 575 => to_unsigned(4018, 12), 576 => to_unsigned(872, 12), 577 => to_unsigned(2213, 12), 578 => to_unsigned(2009, 12), 579 => to_unsigned(3776, 12), 580 => to_unsigned(2266, 12), 581 => to_unsigned(1136, 12), 582 => to_unsigned(1709, 12), 583 => to_unsigned(3595, 12), 584 => to_unsigned(592, 12), 585 => to_unsigned(3604, 12), 586 => to_unsigned(1684, 12), 587 => to_unsigned(3356, 12), 588 => to_unsigned(1463, 12), 589 => to_unsigned(3057, 12), 590 => to_unsigned(3474, 12), 591 => to_unsigned(2377, 12), 592 => to_unsigned(1506, 12), 593 => to_unsigned(1347, 12), 594 => to_unsigned(2689, 12), 595 => to_unsigned(1605, 12), 596 => to_unsigned(1379, 12), 597 => to_unsigned(403, 12), 598 => to_unsigned(1884, 12), 599 => to_unsigned(531, 12), 600 => to_unsigned(3628, 12), 601 => to_unsigned(2098, 12), 602 => to_unsigned(3331, 12), 603 => to_unsigned(275, 12), 604 => to_unsigned(1461, 12), 605 => to_unsigned(501, 12), 606 => to_unsigned(522, 12), 607 => to_unsigned(3953, 12), 608 => to_unsigned(612, 12), 609 => to_unsigned(483, 12), 610 => to_unsigned(1853, 12), 611 => to_unsigned(2642, 12), 612 => to_unsigned(2321, 12), 613 => to_unsigned(2922, 12), 614 => to_unsigned(2493, 12), 615 => to_unsigned(950, 12), 616 => to_unsigned(1717, 12), 617 => to_unsigned(3932, 12), 618 => to_unsigned(2660, 12), 619 => to_unsigned(2703, 12), 620 => to_unsigned(933, 12), 621 => to_unsigned(3890, 12), 622 => to_unsigned(758, 12), 623 => to_unsigned(4006, 12), 624 => to_unsigned(3467, 12), 625 => to_unsigned(1743, 12), 626 => to_unsigned(234, 12), 627 => to_unsigned(2870, 12), 628 => to_unsigned(3893, 12), 629 => to_unsigned(2760, 12), 630 => to_unsigned(4029, 12), 631 => to_unsigned(3947, 12), 632 => to_unsigned(2649, 12), 633 => to_unsigned(3535, 12), 634 => to_unsigned(2639, 12), 635 => to_unsigned(2368, 12), 636 => to_unsigned(175, 12), 637 => to_unsigned(1973, 12), 638 => to_unsigned(1914, 12), 639 => to_unsigned(3816, 12), 640 => to_unsigned(3284, 12), 641 => to_unsigned(493, 12), 642 => to_unsigned(1487, 12), 643 => to_unsigned(1961, 12), 644 => to_unsigned(2857, 12), 645 => to_unsigned(1561, 12), 646 => to_unsigned(1484, 12), 647 => to_unsigned(2512, 12), 648 => to_unsigned(2514, 12), 649 => to_unsigned(3373, 12), 650 => to_unsigned(91, 12), 651 => to_unsigned(2073, 12), 652 => to_unsigned(2158, 12), 653 => to_unsigned(1679, 12), 654 => to_unsigned(1588, 12), 655 => to_unsigned(1316, 12), 656 => to_unsigned(3916, 12), 657 => to_unsigned(2382, 12), 658 => to_unsigned(1527, 12), 659 => to_unsigned(1865, 12), 660 => to_unsigned(2972, 12), 661 => to_unsigned(1832, 12), 662 => to_unsigned(3369, 12), 663 => to_unsigned(2013, 12), 664 => to_unsigned(3629, 12), 665 => to_unsigned(1546, 12), 666 => to_unsigned(2846, 12), 667 => to_unsigned(3592, 12), 668 => to_unsigned(3814, 12), 669 => to_unsigned(1156, 12), 670 => to_unsigned(4083, 12), 671 => to_unsigned(3534, 12), 672 => to_unsigned(104, 12), 673 => to_unsigned(3480, 12), 674 => to_unsigned(2919, 12), 675 => to_unsigned(712, 12), 676 => to_unsigned(341, 12), 677 => to_unsigned(2193, 12), 678 => to_unsigned(3178, 12), 679 => to_unsigned(3207, 12), 680 => to_unsigned(905, 12), 681 => to_unsigned(872, 12), 682 => to_unsigned(4053, 12), 683 => to_unsigned(2945, 12), 684 => to_unsigned(415, 12), 685 => to_unsigned(2457, 12), 686 => to_unsigned(824, 12), 687 => to_unsigned(1705, 12), 688 => to_unsigned(2742, 12), 689 => to_unsigned(220, 12), 690 => to_unsigned(3717, 12), 691 => to_unsigned(225, 12), 692 => to_unsigned(1671, 12), 693 => to_unsigned(624, 12), 694 => to_unsigned(4011, 12), 695 => to_unsigned(3052, 12), 696 => to_unsigned(1577, 12), 697 => to_unsigned(204, 12), 698 => to_unsigned(2818, 12), 699 => to_unsigned(918, 12), 700 => to_unsigned(3170, 12), 701 => to_unsigned(1906, 12), 702 => to_unsigned(2694, 12), 703 => to_unsigned(1018, 12), 704 => to_unsigned(1624, 12), 705 => to_unsigned(1836, 12), 706 => to_unsigned(2580, 12), 707 => to_unsigned(602, 12), 708 => to_unsigned(1075, 12), 709 => to_unsigned(891, 12), 710 => to_unsigned(1777, 12), 711 => to_unsigned(2678, 12), 712 => to_unsigned(171, 12), 713 => to_unsigned(3523, 12), 714 => to_unsigned(3855, 12), 715 => to_unsigned(2349, 12), 716 => to_unsigned(3810, 12), 717 => to_unsigned(2780, 12), 718 => to_unsigned(3764, 12), 719 => to_unsigned(1634, 12), 720 => to_unsigned(1881, 12), 721 => to_unsigned(2432, 12), 722 => to_unsigned(1587, 12), 723 => to_unsigned(507, 12), 724 => to_unsigned(2938, 12), 725 => to_unsigned(1670, 12), 726 => to_unsigned(2478, 12), 727 => to_unsigned(4018, 12), 728 => to_unsigned(2418, 12), 729 => to_unsigned(2712, 12), 730 => to_unsigned(386, 12), 731 => to_unsigned(2217, 12), 732 => to_unsigned(3398, 12), 733 => to_unsigned(2358, 12), 734 => to_unsigned(1631, 12), 735 => to_unsigned(2717, 12), 736 => to_unsigned(1439, 12), 737 => to_unsigned(488, 12), 738 => to_unsigned(2638, 12), 739 => to_unsigned(3756, 12), 740 => to_unsigned(3767, 12), 741 => to_unsigned(2502, 12), 742 => to_unsigned(119, 12), 743 => to_unsigned(1418, 12), 744 => to_unsigned(3716, 12), 745 => to_unsigned(2493, 12), 746 => to_unsigned(431, 12), 747 => to_unsigned(577, 12), 748 => to_unsigned(2855, 12), 749 => to_unsigned(2074, 12), 750 => to_unsigned(1667, 12), 751 => to_unsigned(1253, 12), 752 => to_unsigned(186, 12), 753 => to_unsigned(608, 12), 754 => to_unsigned(3985, 12), 755 => to_unsigned(2935, 12), 756 => to_unsigned(90, 12), 757 => to_unsigned(1802, 12), 758 => to_unsigned(2457, 12), 759 => to_unsigned(3615, 12), 760 => to_unsigned(1193, 12), 761 => to_unsigned(4032, 12), 762 => to_unsigned(2853, 12), 763 => to_unsigned(1782, 12), 764 => to_unsigned(741, 12), 765 => to_unsigned(3360, 12), 766 => to_unsigned(1420, 12), 767 => to_unsigned(2156, 12), 768 => to_unsigned(364, 12), 769 => to_unsigned(552, 12), 770 => to_unsigned(3104, 12), 771 => to_unsigned(2615, 12), 772 => to_unsigned(2733, 12), 773 => to_unsigned(3317, 12), 774 => to_unsigned(1816, 12), 775 => to_unsigned(1513, 12), 776 => to_unsigned(2466, 12), 777 => to_unsigned(3879, 12), 778 => to_unsigned(1950, 12), 779 => to_unsigned(2870, 12), 780 => to_unsigned(3379, 12), 781 => to_unsigned(687, 12), 782 => to_unsigned(749, 12), 783 => to_unsigned(1059, 12), 784 => to_unsigned(3649, 12), 785 => to_unsigned(3180, 12), 786 => to_unsigned(2427, 12), 787 => to_unsigned(2690, 12), 788 => to_unsigned(1530, 12), 789 => to_unsigned(979, 12), 790 => to_unsigned(729, 12), 791 => to_unsigned(2809, 12), 792 => to_unsigned(3081, 12), 793 => to_unsigned(904, 12), 794 => to_unsigned(4028, 12), 795 => to_unsigned(2530, 12), 796 => to_unsigned(1661, 12), 797 => to_unsigned(1839, 12), 798 => to_unsigned(3702, 12), 799 => to_unsigned(2561, 12), 800 => to_unsigned(1156, 12), 801 => to_unsigned(1349, 12), 802 => to_unsigned(3224, 12), 803 => to_unsigned(1957, 12), 804 => to_unsigned(2949, 12), 805 => to_unsigned(3123, 12), 806 => to_unsigned(839, 12), 807 => to_unsigned(1514, 12), 808 => to_unsigned(1784, 12), 809 => to_unsigned(3612, 12), 810 => to_unsigned(1653, 12), 811 => to_unsigned(579, 12), 812 => to_unsigned(2814, 12), 813 => to_unsigned(1421, 12), 814 => to_unsigned(2725, 12), 815 => to_unsigned(192, 12), 816 => to_unsigned(1163, 12), 817 => to_unsigned(629, 12), 818 => to_unsigned(2388, 12), 819 => to_unsigned(316, 12), 820 => to_unsigned(2619, 12), 821 => to_unsigned(1377, 12), 822 => to_unsigned(1181, 12), 823 => to_unsigned(854, 12), 824 => to_unsigned(474, 12), 825 => to_unsigned(1351, 12), 826 => to_unsigned(2529, 12), 827 => to_unsigned(166, 12), 828 => to_unsigned(3684, 12), 829 => to_unsigned(3089, 12), 830 => to_unsigned(3849, 12), 831 => to_unsigned(621, 12), 832 => to_unsigned(793, 12), 833 => to_unsigned(677, 12), 834 => to_unsigned(1916, 12), 835 => to_unsigned(2129, 12), 836 => to_unsigned(1563, 12), 837 => to_unsigned(2522, 12), 838 => to_unsigned(2138, 12), 839 => to_unsigned(3534, 12), 840 => to_unsigned(3254, 12), 841 => to_unsigned(2014, 12), 842 => to_unsigned(2599, 12), 843 => to_unsigned(2739, 12), 844 => to_unsigned(241, 12), 845 => to_unsigned(2918, 12), 846 => to_unsigned(2023, 12), 847 => to_unsigned(3324, 12), 848 => to_unsigned(1733, 12), 849 => to_unsigned(1912, 12), 850 => to_unsigned(2729, 12), 851 => to_unsigned(2941, 12), 852 => to_unsigned(2307, 12), 853 => to_unsigned(3644, 12), 854 => to_unsigned(78, 12), 855 => to_unsigned(2842, 12), 856 => to_unsigned(342, 12), 857 => to_unsigned(1144, 12), 858 => to_unsigned(1013, 12), 859 => to_unsigned(2738, 12), 860 => to_unsigned(339, 12), 861 => to_unsigned(1070, 12), 862 => to_unsigned(3018, 12), 863 => to_unsigned(749, 12), 864 => to_unsigned(854, 12), 865 => to_unsigned(2674, 12), 866 => to_unsigned(2380, 12), 867 => to_unsigned(1363, 12), 868 => to_unsigned(3869, 12), 869 => to_unsigned(2401, 12), 870 => to_unsigned(1528, 12), 871 => to_unsigned(752, 12), 872 => to_unsigned(2371, 12), 873 => to_unsigned(218, 12), 874 => to_unsigned(988, 12), 875 => to_unsigned(3631, 12), 876 => to_unsigned(739, 12), 877 => to_unsigned(2979, 12), 878 => to_unsigned(1203, 12), 879 => to_unsigned(201, 12), 880 => to_unsigned(604, 12), 881 => to_unsigned(3157, 12), 882 => to_unsigned(2488, 12), 883 => to_unsigned(3086, 12), 884 => to_unsigned(2383, 12), 885 => to_unsigned(1272, 12), 886 => to_unsigned(2206, 12), 887 => to_unsigned(499, 12), 888 => to_unsigned(3837, 12), 889 => to_unsigned(3249, 12), 890 => to_unsigned(3208, 12), 891 => to_unsigned(496, 12), 892 => to_unsigned(2875, 12), 893 => to_unsigned(3220, 12), 894 => to_unsigned(1754, 12), 895 => to_unsigned(3637, 12), 896 => to_unsigned(1147, 12), 897 => to_unsigned(3086, 12), 898 => to_unsigned(1180, 12), 899 => to_unsigned(4008, 12), 900 => to_unsigned(3036, 12), 901 => to_unsigned(2259, 12), 902 => to_unsigned(2292, 12), 903 => to_unsigned(1955, 12), 904 => to_unsigned(3587, 12), 905 => to_unsigned(1651, 12), 906 => to_unsigned(1357, 12), 907 => to_unsigned(2384, 12), 908 => to_unsigned(2597, 12), 909 => to_unsigned(3147, 12), 910 => to_unsigned(1998, 12), 911 => to_unsigned(1098, 12), 912 => to_unsigned(3254, 12), 913 => to_unsigned(3161, 12), 914 => to_unsigned(163, 12), 915 => to_unsigned(1497, 12), 916 => to_unsigned(3246, 12), 917 => to_unsigned(161, 12), 918 => to_unsigned(201, 12), 919 => to_unsigned(2906, 12), 920 => to_unsigned(586, 12), 921 => to_unsigned(346, 12), 922 => to_unsigned(3334, 12), 923 => to_unsigned(1385, 12), 924 => to_unsigned(1663, 12), 925 => to_unsigned(1828, 12), 926 => to_unsigned(3869, 12), 927 => to_unsigned(2451, 12), 928 => to_unsigned(579, 12), 929 => to_unsigned(2868, 12), 930 => to_unsigned(2722, 12), 931 => to_unsigned(3176, 12), 932 => to_unsigned(2418, 12), 933 => to_unsigned(3304, 12), 934 => to_unsigned(1023, 12), 935 => to_unsigned(3778, 12), 936 => to_unsigned(1011, 12), 937 => to_unsigned(455, 12), 938 => to_unsigned(1757, 12), 939 => to_unsigned(242, 12), 940 => to_unsigned(1937, 12), 941 => to_unsigned(2992, 12), 942 => to_unsigned(183, 12), 943 => to_unsigned(3241, 12), 944 => to_unsigned(54, 12), 945 => to_unsigned(1885, 12), 946 => to_unsigned(3862, 12), 947 => to_unsigned(2465, 12), 948 => to_unsigned(1485, 12), 949 => to_unsigned(1425, 12), 950 => to_unsigned(263, 12), 951 => to_unsigned(2862, 12), 952 => to_unsigned(1700, 12), 953 => to_unsigned(2756, 12), 954 => to_unsigned(539, 12), 955 => to_unsigned(1812, 12), 956 => to_unsigned(1514, 12), 957 => to_unsigned(2694, 12), 958 => to_unsigned(2161, 12), 959 => to_unsigned(3147, 12), 960 => to_unsigned(1966, 12), 961 => to_unsigned(3479, 12), 962 => to_unsigned(1481, 12), 963 => to_unsigned(1784, 12), 964 => to_unsigned(1141, 12), 965 => to_unsigned(1502, 12), 966 => to_unsigned(1849, 12), 967 => to_unsigned(1575, 12), 968 => to_unsigned(3087, 12), 969 => to_unsigned(1292, 12), 970 => to_unsigned(2586, 12), 971 => to_unsigned(760, 12), 972 => to_unsigned(2181, 12), 973 => to_unsigned(2942, 12), 974 => to_unsigned(1381, 12), 975 => to_unsigned(3653, 12), 976 => to_unsigned(1592, 12), 977 => to_unsigned(338, 12), 978 => to_unsigned(3469, 12), 979 => to_unsigned(309, 12), 980 => to_unsigned(3198, 12), 981 => to_unsigned(2240, 12), 982 => to_unsigned(2037, 12), 983 => to_unsigned(1810, 12), 984 => to_unsigned(2363, 12), 985 => to_unsigned(3966, 12), 986 => to_unsigned(3612, 12), 987 => to_unsigned(102, 12), 988 => to_unsigned(1157, 12), 989 => to_unsigned(3027, 12), 990 => to_unsigned(81, 12), 991 => to_unsigned(685, 12), 992 => to_unsigned(430, 12), 993 => to_unsigned(2108, 12), 994 => to_unsigned(3046, 12), 995 => to_unsigned(2969, 12), 996 => to_unsigned(3869, 12), 997 => to_unsigned(654, 12), 998 => to_unsigned(3834, 12), 999 => to_unsigned(3779, 12), 1000 => to_unsigned(482, 12), 1001 => to_unsigned(305, 12), 1002 => to_unsigned(3011, 12), 1003 => to_unsigned(1447, 12), 1004 => to_unsigned(4043, 12), 1005 => to_unsigned(1064, 12), 1006 => to_unsigned(681, 12), 1007 => to_unsigned(1749, 12), 1008 => to_unsigned(1052, 12), 1009 => to_unsigned(344, 12), 1010 => to_unsigned(2630, 12), 1011 => to_unsigned(3594, 12), 1012 => to_unsigned(1873, 12), 1013 => to_unsigned(2113, 12), 1014 => to_unsigned(1298, 12), 1015 => to_unsigned(2383, 12), 1016 => to_unsigned(867, 12), 1017 => to_unsigned(508, 12), 1018 => to_unsigned(3532, 12), 1019 => to_unsigned(741, 12), 1020 => to_unsigned(1468, 12), 1021 => to_unsigned(1667, 12), 1022 => to_unsigned(437, 12), 1023 => to_unsigned(261, 12), 1024 => to_unsigned(3006, 12), 1025 => to_unsigned(2234, 12), 1026 => to_unsigned(977, 12), 1027 => to_unsigned(3147, 12), 1028 => to_unsigned(3134, 12), 1029 => to_unsigned(1660, 12), 1030 => to_unsigned(1203, 12), 1031 => to_unsigned(4013, 12), 1032 => to_unsigned(916, 12), 1033 => to_unsigned(1223, 12), 1034 => to_unsigned(2558, 12), 1035 => to_unsigned(1595, 12), 1036 => to_unsigned(3162, 12), 1037 => to_unsigned(3617, 12), 1038 => to_unsigned(2403, 12), 1039 => to_unsigned(3803, 12), 1040 => to_unsigned(1882, 12), 1041 => to_unsigned(38, 12), 1042 => to_unsigned(3429, 12), 1043 => to_unsigned(1562, 12), 1044 => to_unsigned(474, 12), 1045 => to_unsigned(2606, 12), 1046 => to_unsigned(4054, 12), 1047 => to_unsigned(2048, 12), 1048 => to_unsigned(2900, 12), 1049 => to_unsigned(3829, 12), 1050 => to_unsigned(1092, 12), 1051 => to_unsigned(1615, 12), 1052 => to_unsigned(764, 12), 1053 => to_unsigned(838, 12), 1054 => to_unsigned(1883, 12), 1055 => to_unsigned(3711, 12), 1056 => to_unsigned(2965, 12), 1057 => to_unsigned(347, 12), 1058 => to_unsigned(1198, 12), 1059 => to_unsigned(3982, 12), 1060 => to_unsigned(3671, 12), 1061 => to_unsigned(397, 12), 1062 => to_unsigned(2428, 12), 1063 => to_unsigned(2943, 12), 1064 => to_unsigned(2977, 12), 1065 => to_unsigned(1662, 12), 1066 => to_unsigned(3722, 12), 1067 => to_unsigned(2996, 12), 1068 => to_unsigned(3164, 12), 1069 => to_unsigned(51, 12), 1070 => to_unsigned(4079, 12), 1071 => to_unsigned(2424, 12), 1072 => to_unsigned(3117, 12), 1073 => to_unsigned(3418, 12), 1074 => to_unsigned(1824, 12), 1075 => to_unsigned(4093, 12), 1076 => to_unsigned(1685, 12), 1077 => to_unsigned(651, 12), 1078 => to_unsigned(3411, 12), 1079 => to_unsigned(1131, 12), 1080 => to_unsigned(889, 12), 1081 => to_unsigned(2068, 12), 1082 => to_unsigned(3239, 12), 1083 => to_unsigned(3273, 12), 1084 => to_unsigned(490, 12), 1085 => to_unsigned(3478, 12), 1086 => to_unsigned(2916, 12), 1087 => to_unsigned(3292, 12), 1088 => to_unsigned(629, 12), 1089 => to_unsigned(3728, 12), 1090 => to_unsigned(3299, 12), 1091 => to_unsigned(240, 12), 1092 => to_unsigned(3328, 12), 1093 => to_unsigned(2265, 12), 1094 => to_unsigned(996, 12), 1095 => to_unsigned(2223, 12), 1096 => to_unsigned(2616, 12), 1097 => to_unsigned(3406, 12), 1098 => to_unsigned(2261, 12), 1099 => to_unsigned(1660, 12), 1100 => to_unsigned(1081, 12), 1101 => to_unsigned(3807, 12), 1102 => to_unsigned(2378, 12), 1103 => to_unsigned(2785, 12), 1104 => to_unsigned(1465, 12), 1105 => to_unsigned(36, 12), 1106 => to_unsigned(927, 12), 1107 => to_unsigned(2088, 12), 1108 => to_unsigned(375, 12), 1109 => to_unsigned(2182, 12), 1110 => to_unsigned(3862, 12), 1111 => to_unsigned(3875, 12), 1112 => to_unsigned(3729, 12), 1113 => to_unsigned(1734, 12), 1114 => to_unsigned(259, 12), 1115 => to_unsigned(2217, 12), 1116 => to_unsigned(907, 12), 1117 => to_unsigned(2571, 12), 1118 => to_unsigned(401, 12), 1119 => to_unsigned(250, 12), 1120 => to_unsigned(1847, 12), 1121 => to_unsigned(3321, 12), 1122 => to_unsigned(3816, 12), 1123 => to_unsigned(2882, 12), 1124 => to_unsigned(2714, 12), 1125 => to_unsigned(1415, 12), 1126 => to_unsigned(2770, 12), 1127 => to_unsigned(2033, 12), 1128 => to_unsigned(1969, 12), 1129 => to_unsigned(3139, 12), 1130 => to_unsigned(3335, 12), 1131 => to_unsigned(3836, 12), 1132 => to_unsigned(3055, 12), 1133 => to_unsigned(3639, 12), 1134 => to_unsigned(2731, 12), 1135 => to_unsigned(1982, 12), 1136 => to_unsigned(3726, 12), 1137 => to_unsigned(3657, 12), 1138 => to_unsigned(3565, 12), 1139 => to_unsigned(531, 12), 1140 => to_unsigned(3825, 12), 1141 => to_unsigned(1243, 12), 1142 => to_unsigned(1672, 12), 1143 => to_unsigned(1484, 12), 1144 => to_unsigned(498, 12), 1145 => to_unsigned(661, 12), 1146 => to_unsigned(638, 12), 1147 => to_unsigned(2513, 12), 1148 => to_unsigned(315, 12), 1149 => to_unsigned(2817, 12), 1150 => to_unsigned(1113, 12), 1151 => to_unsigned(763, 12), 1152 => to_unsigned(100, 12), 1153 => to_unsigned(3927, 12), 1154 => to_unsigned(59, 12), 1155 => to_unsigned(2884, 12), 1156 => to_unsigned(1594, 12), 1157 => to_unsigned(1055, 12), 1158 => to_unsigned(1508, 12), 1159 => to_unsigned(2712, 12), 1160 => to_unsigned(424, 12), 1161 => to_unsigned(1682, 12), 1162 => to_unsigned(1367, 12), 1163 => to_unsigned(32, 12), 1164 => to_unsigned(2552, 12), 1165 => to_unsigned(1281, 12), 1166 => to_unsigned(2279, 12), 1167 => to_unsigned(3549, 12), 1168 => to_unsigned(1457, 12), 1169 => to_unsigned(1563, 12), 1170 => to_unsigned(975, 12), 1171 => to_unsigned(1597, 12), 1172 => to_unsigned(2628, 12), 1173 => to_unsigned(2210, 12), 1174 => to_unsigned(2756, 12), 1175 => to_unsigned(2756, 12), 1176 => to_unsigned(4032, 12), 1177 => to_unsigned(3821, 12), 1178 => to_unsigned(3580, 12), 1179 => to_unsigned(1437, 12), 1180 => to_unsigned(2838, 12), 1181 => to_unsigned(2742, 12), 1182 => to_unsigned(3103, 12), 1183 => to_unsigned(1040, 12), 1184 => to_unsigned(772, 12), 1185 => to_unsigned(644, 12), 1186 => to_unsigned(2487, 12), 1187 => to_unsigned(3679, 12), 1188 => to_unsigned(2398, 12), 1189 => to_unsigned(3181, 12), 1190 => to_unsigned(3895, 12), 1191 => to_unsigned(3527, 12), 1192 => to_unsigned(962, 12), 1193 => to_unsigned(395, 12), 1194 => to_unsigned(1890, 12), 1195 => to_unsigned(2014, 12), 1196 => to_unsigned(758, 12), 1197 => to_unsigned(1191, 12), 1198 => to_unsigned(2225, 12), 1199 => to_unsigned(3710, 12), 1200 => to_unsigned(1378, 12), 1201 => to_unsigned(4005, 12), 1202 => to_unsigned(3086, 12), 1203 => to_unsigned(2365, 12), 1204 => to_unsigned(1789, 12), 1205 => to_unsigned(1926, 12), 1206 => to_unsigned(1272, 12), 1207 => to_unsigned(1345, 12), 1208 => to_unsigned(2032, 12), 1209 => to_unsigned(1379, 12), 1210 => to_unsigned(2765, 12), 1211 => to_unsigned(1795, 12), 1212 => to_unsigned(1059, 12), 1213 => to_unsigned(2522, 12), 1214 => to_unsigned(4078, 12), 1215 => to_unsigned(2198, 12), 1216 => to_unsigned(3391, 12), 1217 => to_unsigned(3723, 12), 1218 => to_unsigned(2846, 12), 1219 => to_unsigned(2663, 12), 1220 => to_unsigned(3778, 12), 1221 => to_unsigned(2941, 12), 1222 => to_unsigned(1306, 12), 1223 => to_unsigned(320, 12), 1224 => to_unsigned(1484, 12), 1225 => to_unsigned(3336, 12), 1226 => to_unsigned(2167, 12), 1227 => to_unsigned(1217, 12), 1228 => to_unsigned(379, 12), 1229 => to_unsigned(639, 12), 1230 => to_unsigned(3503, 12), 1231 => to_unsigned(1308, 12), 1232 => to_unsigned(2229, 12), 1233 => to_unsigned(4021, 12), 1234 => to_unsigned(1655, 12), 1235 => to_unsigned(1407, 12), 1236 => to_unsigned(2712, 12), 1237 => to_unsigned(3715, 12), 1238 => to_unsigned(3871, 12), 1239 => to_unsigned(3737, 12), 1240 => to_unsigned(1586, 12), 1241 => to_unsigned(2261, 12), 1242 => to_unsigned(2489, 12), 1243 => to_unsigned(1762, 12), 1244 => to_unsigned(3662, 12), 1245 => to_unsigned(215, 12), 1246 => to_unsigned(1717, 12), 1247 => to_unsigned(3381, 12), 1248 => to_unsigned(45, 12), 1249 => to_unsigned(116, 12), 1250 => to_unsigned(3776, 12), 1251 => to_unsigned(1457, 12), 1252 => to_unsigned(1412, 12), 1253 => to_unsigned(3695, 12), 1254 => to_unsigned(3750, 12), 1255 => to_unsigned(2544, 12), 1256 => to_unsigned(1663, 12), 1257 => to_unsigned(2903, 12), 1258 => to_unsigned(748, 12), 1259 => to_unsigned(2164, 12), 1260 => to_unsigned(1755, 12), 1261 => to_unsigned(1262, 12), 1262 => to_unsigned(2896, 12), 1263 => to_unsigned(3073, 12), 1264 => to_unsigned(1379, 12), 1265 => to_unsigned(3523, 12), 1266 => to_unsigned(852, 12), 1267 => to_unsigned(3426, 12), 1268 => to_unsigned(3079, 12), 1269 => to_unsigned(1511, 12), 1270 => to_unsigned(2668, 12), 1271 => to_unsigned(246, 12), 1272 => to_unsigned(3280, 12), 1273 => to_unsigned(3042, 12), 1274 => to_unsigned(526, 12), 1275 => to_unsigned(2242, 12), 1276 => to_unsigned(1556, 12), 1277 => to_unsigned(3989, 12), 1278 => to_unsigned(37, 12), 1279 => to_unsigned(839, 12), 1280 => to_unsigned(153, 12), 1281 => to_unsigned(3392, 12), 1282 => to_unsigned(2498, 12), 1283 => to_unsigned(2483, 12), 1284 => to_unsigned(3156, 12), 1285 => to_unsigned(3032, 12), 1286 => to_unsigned(3366, 12), 1287 => to_unsigned(3920, 12), 1288 => to_unsigned(2898, 12), 1289 => to_unsigned(3353, 12), 1290 => to_unsigned(880, 12), 1291 => to_unsigned(3196, 12), 1292 => to_unsigned(1131, 12), 1293 => to_unsigned(1659, 12), 1294 => to_unsigned(549, 12), 1295 => to_unsigned(926, 12), 1296 => to_unsigned(36, 12), 1297 => to_unsigned(2759, 12), 1298 => to_unsigned(2117, 12), 1299 => to_unsigned(3, 12), 1300 => to_unsigned(972, 12), 1301 => to_unsigned(25, 12), 1302 => to_unsigned(1621, 12), 1303 => to_unsigned(2353, 12), 1304 => to_unsigned(3257, 12), 1305 => to_unsigned(386, 12), 1306 => to_unsigned(75, 12), 1307 => to_unsigned(3165, 12), 1308 => to_unsigned(2615, 12), 1309 => to_unsigned(1217, 12), 1310 => to_unsigned(1844, 12), 1311 => to_unsigned(2139, 12), 1312 => to_unsigned(1718, 12), 1313 => to_unsigned(3532, 12), 1314 => to_unsigned(2143, 12), 1315 => to_unsigned(2895, 12), 1316 => to_unsigned(2974, 12), 1317 => to_unsigned(2583, 12), 1318 => to_unsigned(3260, 12), 1319 => to_unsigned(1532, 12), 1320 => to_unsigned(2915, 12), 1321 => to_unsigned(1285, 12), 1322 => to_unsigned(3928, 12), 1323 => to_unsigned(1577, 12), 1324 => to_unsigned(2384, 12), 1325 => to_unsigned(3790, 12), 1326 => to_unsigned(3075, 12), 1327 => to_unsigned(3835, 12), 1328 => to_unsigned(3559, 12), 1329 => to_unsigned(1062, 12), 1330 => to_unsigned(3565, 12), 1331 => to_unsigned(1861, 12), 1332 => to_unsigned(1245, 12), 1333 => to_unsigned(1746, 12), 1334 => to_unsigned(2267, 12), 1335 => to_unsigned(2684, 12), 1336 => to_unsigned(868, 12), 1337 => to_unsigned(318, 12), 1338 => to_unsigned(1155, 12), 1339 => to_unsigned(3804, 12), 1340 => to_unsigned(1295, 12), 1341 => to_unsigned(127, 12), 1342 => to_unsigned(1148, 12), 1343 => to_unsigned(3, 12), 1344 => to_unsigned(1485, 12), 1345 => to_unsigned(2967, 12), 1346 => to_unsigned(630, 12), 1347 => to_unsigned(3751, 12), 1348 => to_unsigned(421, 12), 1349 => to_unsigned(896, 12), 1350 => to_unsigned(1633, 12), 1351 => to_unsigned(490, 12), 1352 => to_unsigned(1059, 12), 1353 => to_unsigned(832, 12), 1354 => to_unsigned(1582, 12), 1355 => to_unsigned(1906, 12), 1356 => to_unsigned(2433, 12), 1357 => to_unsigned(3453, 12), 1358 => to_unsigned(1198, 12), 1359 => to_unsigned(3048, 12), 1360 => to_unsigned(3636, 12), 1361 => to_unsigned(3644, 12), 1362 => to_unsigned(1440, 12), 1363 => to_unsigned(2599, 12), 1364 => to_unsigned(3966, 12), 1365 => to_unsigned(2765, 12), 1366 => to_unsigned(3329, 12), 1367 => to_unsigned(2179, 12), 1368 => to_unsigned(272, 12), 1369 => to_unsigned(2229, 12), 1370 => to_unsigned(91, 12), 1371 => to_unsigned(1966, 12), 1372 => to_unsigned(2563, 12), 1373 => to_unsigned(788, 12), 1374 => to_unsigned(4056, 12), 1375 => to_unsigned(1054, 12), 1376 => to_unsigned(3809, 12), 1377 => to_unsigned(1135, 12), 1378 => to_unsigned(1201, 12), 1379 => to_unsigned(2835, 12), 1380 => to_unsigned(2797, 12), 1381 => to_unsigned(2950, 12), 1382 => to_unsigned(3555, 12), 1383 => to_unsigned(45, 12), 1384 => to_unsigned(3046, 12), 1385 => to_unsigned(1602, 12), 1386 => to_unsigned(3773, 12), 1387 => to_unsigned(2174, 12), 1388 => to_unsigned(2174, 12), 1389 => to_unsigned(1735, 12), 1390 => to_unsigned(498, 12), 1391 => to_unsigned(1057, 12), 1392 => to_unsigned(1808, 12), 1393 => to_unsigned(3180, 12), 1394 => to_unsigned(808, 12), 1395 => to_unsigned(3228, 12), 1396 => to_unsigned(576, 12), 1397 => to_unsigned(220, 12), 1398 => to_unsigned(3789, 12), 1399 => to_unsigned(998, 12), 1400 => to_unsigned(4005, 12), 1401 => to_unsigned(2036, 12), 1402 => to_unsigned(1304, 12), 1403 => to_unsigned(1403, 12), 1404 => to_unsigned(2604, 12), 1405 => to_unsigned(14, 12), 1406 => to_unsigned(1437, 12), 1407 => to_unsigned(3401, 12), 1408 => to_unsigned(2579, 12), 1409 => to_unsigned(1629, 12), 1410 => to_unsigned(2080, 12), 1411 => to_unsigned(1098, 12), 1412 => to_unsigned(884, 12), 1413 => to_unsigned(965, 12), 1414 => to_unsigned(58, 12), 1415 => to_unsigned(207, 12), 1416 => to_unsigned(3698, 12), 1417 => to_unsigned(1850, 12), 1418 => to_unsigned(3254, 12), 1419 => to_unsigned(843, 12), 1420 => to_unsigned(3009, 12), 1421 => to_unsigned(2827, 12), 1422 => to_unsigned(3129, 12), 1423 => to_unsigned(2055, 12), 1424 => to_unsigned(522, 12), 1425 => to_unsigned(1997, 12), 1426 => to_unsigned(3124, 12), 1427 => to_unsigned(1817, 12), 1428 => to_unsigned(399, 12), 1429 => to_unsigned(1551, 12), 1430 => to_unsigned(3965, 12), 1431 => to_unsigned(1849, 12), 1432 => to_unsigned(3918, 12), 1433 => to_unsigned(3133, 12), 1434 => to_unsigned(3515, 12), 1435 => to_unsigned(2734, 12), 1436 => to_unsigned(3990, 12), 1437 => to_unsigned(3462, 12), 1438 => to_unsigned(3281, 12), 1439 => to_unsigned(1179, 12), 1440 => to_unsigned(3642, 12), 1441 => to_unsigned(1855, 12), 1442 => to_unsigned(1191, 12), 1443 => to_unsigned(1179, 12), 1444 => to_unsigned(1389, 12), 1445 => to_unsigned(49, 12), 1446 => to_unsigned(2064, 12), 1447 => to_unsigned(398, 12), 1448 => to_unsigned(3411, 12), 1449 => to_unsigned(1638, 12), 1450 => to_unsigned(3991, 12), 1451 => to_unsigned(1187, 12), 1452 => to_unsigned(925, 12), 1453 => to_unsigned(2605, 12), 1454 => to_unsigned(25, 12), 1455 => to_unsigned(433, 12), 1456 => to_unsigned(557, 12), 1457 => to_unsigned(244, 12), 1458 => to_unsigned(3486, 12), 1459 => to_unsigned(3836, 12), 1460 => to_unsigned(2440, 12), 1461 => to_unsigned(1284, 12), 1462 => to_unsigned(3271, 12), 1463 => to_unsigned(2187, 12), 1464 => to_unsigned(1503, 12), 1465 => to_unsigned(3502, 12), 1466 => to_unsigned(3888, 12), 1467 => to_unsigned(1003, 12), 1468 => to_unsigned(3006, 12), 1469 => to_unsigned(2086, 12), 1470 => to_unsigned(1180, 12), 1471 => to_unsigned(251, 12), 1472 => to_unsigned(3695, 12), 1473 => to_unsigned(2042, 12), 1474 => to_unsigned(369, 12), 1475 => to_unsigned(2456, 12), 1476 => to_unsigned(3257, 12), 1477 => to_unsigned(2032, 12), 1478 => to_unsigned(604, 12), 1479 => to_unsigned(2110, 12), 1480 => to_unsigned(1782, 12), 1481 => to_unsigned(129, 12), 1482 => to_unsigned(2593, 12), 1483 => to_unsigned(208, 12), 1484 => to_unsigned(1049, 12), 1485 => to_unsigned(1356, 12), 1486 => to_unsigned(249, 12), 1487 => to_unsigned(3582, 12), 1488 => to_unsigned(4027, 12), 1489 => to_unsigned(460, 12), 1490 => to_unsigned(3428, 12), 1491 => to_unsigned(2069, 12), 1492 => to_unsigned(1675, 12), 1493 => to_unsigned(1668, 12), 1494 => to_unsigned(932, 12), 1495 => to_unsigned(2019, 12), 1496 => to_unsigned(3015, 12), 1497 => to_unsigned(3505, 12), 1498 => to_unsigned(518, 12), 1499 => to_unsigned(2453, 12), 1500 => to_unsigned(2196, 12), 1501 => to_unsigned(3905, 12), 1502 => to_unsigned(3634, 12), 1503 => to_unsigned(2026, 12), 1504 => to_unsigned(3945, 12), 1505 => to_unsigned(3871, 12), 1506 => to_unsigned(1956, 12), 1507 => to_unsigned(2346, 12), 1508 => to_unsigned(3885, 12), 1509 => to_unsigned(1396, 12), 1510 => to_unsigned(3082, 12), 1511 => to_unsigned(1119, 12), 1512 => to_unsigned(2390, 12), 1513 => to_unsigned(2086, 12), 1514 => to_unsigned(3936, 12), 1515 => to_unsigned(2225, 12), 1516 => to_unsigned(1220, 12), 1517 => to_unsigned(3045, 12), 1518 => to_unsigned(1960, 12), 1519 => to_unsigned(2095, 12), 1520 => to_unsigned(3549, 12), 1521 => to_unsigned(3126, 12), 1522 => to_unsigned(3825, 12), 1523 => to_unsigned(1202, 12), 1524 => to_unsigned(368, 12), 1525 => to_unsigned(973, 12), 1526 => to_unsigned(3800, 12), 1527 => to_unsigned(1729, 12), 1528 => to_unsigned(1328, 12), 1529 => to_unsigned(3465, 12), 1530 => to_unsigned(943, 12), 1531 => to_unsigned(904, 12), 1532 => to_unsigned(149, 12), 1533 => to_unsigned(3963, 12), 1534 => to_unsigned(1310, 12), 1535 => to_unsigned(2076, 12), 1536 => to_unsigned(893, 12), 1537 => to_unsigned(3400, 12), 1538 => to_unsigned(636, 12), 1539 => to_unsigned(3709, 12), 1540 => to_unsigned(2151, 12), 1541 => to_unsigned(2597, 12), 1542 => to_unsigned(3322, 12), 1543 => to_unsigned(3262, 12), 1544 => to_unsigned(3221, 12), 1545 => to_unsigned(1988, 12), 1546 => to_unsigned(3525, 12), 1547 => to_unsigned(3284, 12), 1548 => to_unsigned(2531, 12), 1549 => to_unsigned(262, 12), 1550 => to_unsigned(248, 12), 1551 => to_unsigned(982, 12), 1552 => to_unsigned(652, 12), 1553 => to_unsigned(863, 12), 1554 => to_unsigned(4061, 12), 1555 => to_unsigned(3022, 12), 1556 => to_unsigned(3802, 12), 1557 => to_unsigned(3123, 12), 1558 => to_unsigned(2136, 12), 1559 => to_unsigned(349, 12), 1560 => to_unsigned(1212, 12), 1561 => to_unsigned(1497, 12), 1562 => to_unsigned(3324, 12), 1563 => to_unsigned(589, 12), 1564 => to_unsigned(3971, 12), 1565 => to_unsigned(64, 12), 1566 => to_unsigned(2935, 12), 1567 => to_unsigned(642, 12), 1568 => to_unsigned(2871, 12), 1569 => to_unsigned(1704, 12), 1570 => to_unsigned(469, 12), 1571 => to_unsigned(3207, 12), 1572 => to_unsigned(2726, 12), 1573 => to_unsigned(25, 12), 1574 => to_unsigned(2246, 12), 1575 => to_unsigned(2399, 12), 1576 => to_unsigned(4000, 12), 1577 => to_unsigned(685, 12), 1578 => to_unsigned(1037, 12), 1579 => to_unsigned(2538, 12), 1580 => to_unsigned(1877, 12), 1581 => to_unsigned(223, 12), 1582 => to_unsigned(3319, 12), 1583 => to_unsigned(2749, 12), 1584 => to_unsigned(3993, 12), 1585 => to_unsigned(236, 12), 1586 => to_unsigned(77, 12), 1587 => to_unsigned(437, 12), 1588 => to_unsigned(1837, 12), 1589 => to_unsigned(1859, 12), 1590 => to_unsigned(1837, 12), 1591 => to_unsigned(3825, 12), 1592 => to_unsigned(1253, 12), 1593 => to_unsigned(1521, 12), 1594 => to_unsigned(2668, 12), 1595 => to_unsigned(3405, 12), 1596 => to_unsigned(2855, 12), 1597 => to_unsigned(90, 12), 1598 => to_unsigned(2468, 12), 1599 => to_unsigned(3405, 12), 1600 => to_unsigned(2193, 12), 1601 => to_unsigned(1054, 12), 1602 => to_unsigned(3571, 12), 1603 => to_unsigned(1508, 12), 1604 => to_unsigned(999, 12), 1605 => to_unsigned(1395, 12), 1606 => to_unsigned(3874, 12), 1607 => to_unsigned(1740, 12), 1608 => to_unsigned(1156, 12), 1609 => to_unsigned(214, 12), 1610 => to_unsigned(1105, 12), 1611 => to_unsigned(2487, 12), 1612 => to_unsigned(2408, 12), 1613 => to_unsigned(186, 12), 1614 => to_unsigned(99, 12), 1615 => to_unsigned(200, 12), 1616 => to_unsigned(2393, 12), 1617 => to_unsigned(1740, 12), 1618 => to_unsigned(2331, 12), 1619 => to_unsigned(3995, 12), 1620 => to_unsigned(2413, 12), 1621 => to_unsigned(1046, 12), 1622 => to_unsigned(394, 12), 1623 => to_unsigned(3927, 12), 1624 => to_unsigned(495, 12), 1625 => to_unsigned(3483, 12), 1626 => to_unsigned(2777, 12), 1627 => to_unsigned(1955, 12), 1628 => to_unsigned(2130, 12), 1629 => to_unsigned(1664, 12), 1630 => to_unsigned(2268, 12), 1631 => to_unsigned(323, 12), 1632 => to_unsigned(437, 12), 1633 => to_unsigned(297, 12), 1634 => to_unsigned(3323, 12), 1635 => to_unsigned(3198, 12), 1636 => to_unsigned(3227, 12), 1637 => to_unsigned(1839, 12), 1638 => to_unsigned(260, 12), 1639 => to_unsigned(2194, 12), 1640 => to_unsigned(134, 12), 1641 => to_unsigned(2765, 12), 1642 => to_unsigned(1490, 12), 1643 => to_unsigned(2731, 12), 1644 => to_unsigned(3336, 12), 1645 => to_unsigned(2393, 12), 1646 => to_unsigned(3089, 12), 1647 => to_unsigned(51, 12), 1648 => to_unsigned(3792, 12), 1649 => to_unsigned(2900, 12), 1650 => to_unsigned(337, 12), 1651 => to_unsigned(4045, 12), 1652 => to_unsigned(2304, 12), 1653 => to_unsigned(466, 12), 1654 => to_unsigned(1445, 12), 1655 => to_unsigned(2462, 12), 1656 => to_unsigned(1876, 12), 1657 => to_unsigned(3177, 12), 1658 => to_unsigned(436, 12), 1659 => to_unsigned(3975, 12), 1660 => to_unsigned(1095, 12), 1661 => to_unsigned(3772, 12), 1662 => to_unsigned(2823, 12), 1663 => to_unsigned(2254, 12), 1664 => to_unsigned(902, 12), 1665 => to_unsigned(808, 12), 1666 => to_unsigned(2511, 12), 1667 => to_unsigned(3462, 12), 1668 => to_unsigned(1861, 12), 1669 => to_unsigned(902, 12), 1670 => to_unsigned(727, 12), 1671 => to_unsigned(1302, 12), 1672 => to_unsigned(306, 12), 1673 => to_unsigned(1756, 12), 1674 => to_unsigned(1099, 12), 1675 => to_unsigned(2984, 12), 1676 => to_unsigned(903, 12), 1677 => to_unsigned(547, 12), 1678 => to_unsigned(2706, 12), 1679 => to_unsigned(4016, 12), 1680 => to_unsigned(3838, 12), 1681 => to_unsigned(1807, 12), 1682 => to_unsigned(3211, 12), 1683 => to_unsigned(1490, 12), 1684 => to_unsigned(1220, 12), 1685 => to_unsigned(3960, 12), 1686 => to_unsigned(2779, 12), 1687 => to_unsigned(628, 12), 1688 => to_unsigned(2113, 12), 1689 => to_unsigned(1991, 12), 1690 => to_unsigned(1043, 12), 1691 => to_unsigned(1483, 12), 1692 => to_unsigned(710, 12), 1693 => to_unsigned(3552, 12), 1694 => to_unsigned(2629, 12), 1695 => to_unsigned(3885, 12), 1696 => to_unsigned(1703, 12), 1697 => to_unsigned(116, 12), 1698 => to_unsigned(1875, 12), 1699 => to_unsigned(2814, 12), 1700 => to_unsigned(68, 12), 1701 => to_unsigned(405, 12), 1702 => to_unsigned(1692, 12), 1703 => to_unsigned(2225, 12), 1704 => to_unsigned(1944, 12), 1705 => to_unsigned(2918, 12), 1706 => to_unsigned(2187, 12), 1707 => to_unsigned(1909, 12), 1708 => to_unsigned(467, 12), 1709 => to_unsigned(1761, 12), 1710 => to_unsigned(1068, 12), 1711 => to_unsigned(3303, 12), 1712 => to_unsigned(2511, 12), 1713 => to_unsigned(3726, 12), 1714 => to_unsigned(1427, 12), 1715 => to_unsigned(3368, 12), 1716 => to_unsigned(2020, 12), 1717 => to_unsigned(1869, 12), 1718 => to_unsigned(1724, 12), 1719 => to_unsigned(1000, 12), 1720 => to_unsigned(2298, 12), 1721 => to_unsigned(361, 12), 1722 => to_unsigned(2098, 12), 1723 => to_unsigned(308, 12), 1724 => to_unsigned(1917, 12), 1725 => to_unsigned(2906, 12), 1726 => to_unsigned(440, 12), 1727 => to_unsigned(351, 12), 1728 => to_unsigned(4018, 12), 1729 => to_unsigned(2727, 12), 1730 => to_unsigned(1191, 12), 1731 => to_unsigned(1979, 12), 1732 => to_unsigned(427, 12), 1733 => to_unsigned(2213, 12), 1734 => to_unsigned(775, 12), 1735 => to_unsigned(3512, 12), 1736 => to_unsigned(3148, 12), 1737 => to_unsigned(3498, 12), 1738 => to_unsigned(1633, 12), 1739 => to_unsigned(1104, 12), 1740 => to_unsigned(530, 12), 1741 => to_unsigned(2530, 12), 1742 => to_unsigned(433, 12), 1743 => to_unsigned(2886, 12), 1744 => to_unsigned(2649, 12), 1745 => to_unsigned(2815, 12), 1746 => to_unsigned(459, 12), 1747 => to_unsigned(3669, 12), 1748 => to_unsigned(2787, 12), 1749 => to_unsigned(1209, 12), 1750 => to_unsigned(1235, 12), 1751 => to_unsigned(2157, 12), 1752 => to_unsigned(3483, 12), 1753 => to_unsigned(198, 12), 1754 => to_unsigned(3907, 12), 1755 => to_unsigned(512, 12), 1756 => to_unsigned(629, 12), 1757 => to_unsigned(3339, 12), 1758 => to_unsigned(2756, 12), 1759 => to_unsigned(3775, 12), 1760 => to_unsigned(2714, 12), 1761 => to_unsigned(613, 12), 1762 => to_unsigned(1612, 12), 1763 => to_unsigned(3574, 12), 1764 => to_unsigned(3967, 12), 1765 => to_unsigned(3010, 12), 1766 => to_unsigned(2801, 12), 1767 => to_unsigned(4022, 12), 1768 => to_unsigned(2990, 12), 1769 => to_unsigned(1335, 12), 1770 => to_unsigned(246, 12), 1771 => to_unsigned(3511, 12), 1772 => to_unsigned(3199, 12), 1773 => to_unsigned(438, 12), 1774 => to_unsigned(2665, 12), 1775 => to_unsigned(2775, 12), 1776 => to_unsigned(1294, 12), 1777 => to_unsigned(2661, 12), 1778 => to_unsigned(2160, 12), 1779 => to_unsigned(3998, 12), 1780 => to_unsigned(2566, 12), 1781 => to_unsigned(1421, 12), 1782 => to_unsigned(2835, 12), 1783 => to_unsigned(2985, 12), 1784 => to_unsigned(2667, 12), 1785 => to_unsigned(2751, 12), 1786 => to_unsigned(3221, 12), 1787 => to_unsigned(3525, 12), 1788 => to_unsigned(2083, 12), 1789 => to_unsigned(2447, 12), 1790 => to_unsigned(1770, 12), 1791 => to_unsigned(870, 12), 1792 => to_unsigned(3238, 12), 1793 => to_unsigned(547, 12), 1794 => to_unsigned(2054, 12), 1795 => to_unsigned(2236, 12), 1796 => to_unsigned(3221, 12), 1797 => to_unsigned(250, 12), 1798 => to_unsigned(2093, 12), 1799 => to_unsigned(717, 12), 1800 => to_unsigned(983, 12), 1801 => to_unsigned(351, 12), 1802 => to_unsigned(3633, 12), 1803 => to_unsigned(2589, 12), 1804 => to_unsigned(2664, 12), 1805 => to_unsigned(737, 12), 1806 => to_unsigned(2877, 12), 1807 => to_unsigned(1567, 12), 1808 => to_unsigned(3304, 12), 1809 => to_unsigned(474, 12), 1810 => to_unsigned(1825, 12), 1811 => to_unsigned(3285, 12), 1812 => to_unsigned(1424, 12), 1813 => to_unsigned(2568, 12), 1814 => to_unsigned(3440, 12), 1815 => to_unsigned(3583, 12), 1816 => to_unsigned(204, 12), 1817 => to_unsigned(807, 12), 1818 => to_unsigned(3506, 12), 1819 => to_unsigned(908, 12), 1820 => to_unsigned(1224, 12), 1821 => to_unsigned(3739, 12), 1822 => to_unsigned(224, 12), 1823 => to_unsigned(170, 12), 1824 => to_unsigned(2884, 12), 1825 => to_unsigned(3500, 12), 1826 => to_unsigned(1121, 12), 1827 => to_unsigned(2538, 12), 1828 => to_unsigned(3140, 12), 1829 => to_unsigned(1855, 12), 1830 => to_unsigned(2602, 12), 1831 => to_unsigned(2545, 12), 1832 => to_unsigned(918, 12), 1833 => to_unsigned(3408, 12), 1834 => to_unsigned(2104, 12), 1835 => to_unsigned(3664, 12), 1836 => to_unsigned(987, 12), 1837 => to_unsigned(2892, 12), 1838 => to_unsigned(1042, 12), 1839 => to_unsigned(650, 12), 1840 => to_unsigned(415, 12), 1841 => to_unsigned(1017, 12), 1842 => to_unsigned(1340, 12), 1843 => to_unsigned(483, 12), 1844 => to_unsigned(519, 12), 1845 => to_unsigned(1958, 12), 1846 => to_unsigned(2138, 12), 1847 => to_unsigned(449, 12), 1848 => to_unsigned(3537, 12), 1849 => to_unsigned(1801, 12), 1850 => to_unsigned(3882, 12), 1851 => to_unsigned(1731, 12), 1852 => to_unsigned(3544, 12), 1853 => to_unsigned(1127, 12), 1854 => to_unsigned(3719, 12), 1855 => to_unsigned(387, 12), 1856 => to_unsigned(273, 12), 1857 => to_unsigned(1809, 12), 1858 => to_unsigned(2912, 12), 1859 => to_unsigned(2692, 12), 1860 => to_unsigned(3299, 12), 1861 => to_unsigned(2059, 12), 1862 => to_unsigned(463, 12), 1863 => to_unsigned(2904, 12), 1864 => to_unsigned(2914, 12), 1865 => to_unsigned(864, 12), 1866 => to_unsigned(3336, 12), 1867 => to_unsigned(4040, 12), 1868 => to_unsigned(4063, 12), 1869 => to_unsigned(2926, 12), 1870 => to_unsigned(3687, 12), 1871 => to_unsigned(3292, 12), 1872 => to_unsigned(500, 12), 1873 => to_unsigned(2369, 12), 1874 => to_unsigned(98, 12), 1875 => to_unsigned(638, 12), 1876 => to_unsigned(2502, 12), 1877 => to_unsigned(419, 12), 1878 => to_unsigned(3296, 12), 1879 => to_unsigned(3785, 12), 1880 => to_unsigned(82, 12), 1881 => to_unsigned(2163, 12), 1882 => to_unsigned(1246, 12), 1883 => to_unsigned(853, 12), 1884 => to_unsigned(1860, 12), 1885 => to_unsigned(1742, 12), 1886 => to_unsigned(1586, 12), 1887 => to_unsigned(3222, 12), 1888 => to_unsigned(3402, 12), 1889 => to_unsigned(2838, 12), 1890 => to_unsigned(2318, 12), 1891 => to_unsigned(1126, 12), 1892 => to_unsigned(2924, 12), 1893 => to_unsigned(1366, 12), 1894 => to_unsigned(1443, 12), 1895 => to_unsigned(334, 12), 1896 => to_unsigned(1390, 12), 1897 => to_unsigned(101, 12), 1898 => to_unsigned(1005, 12), 1899 => to_unsigned(1733, 12), 1900 => to_unsigned(1520, 12), 1901 => to_unsigned(3928, 12), 1902 => to_unsigned(2189, 12), 1903 => to_unsigned(3064, 12), 1904 => to_unsigned(259, 12), 1905 => to_unsigned(2473, 12), 1906 => to_unsigned(690, 12), 1907 => to_unsigned(58, 12), 1908 => to_unsigned(2602, 12), 1909 => to_unsigned(9, 12), 1910 => to_unsigned(3582, 12), 1911 => to_unsigned(2994, 12), 1912 => to_unsigned(2464, 12), 1913 => to_unsigned(2984, 12), 1914 => to_unsigned(705, 12), 1915 => to_unsigned(3455, 12), 1916 => to_unsigned(1378, 12), 1917 => to_unsigned(1477, 12), 1918 => to_unsigned(2359, 12), 1919 => to_unsigned(813, 12), 1920 => to_unsigned(1059, 12), 1921 => to_unsigned(1173, 12), 1922 => to_unsigned(948, 12), 1923 => to_unsigned(2645, 12), 1924 => to_unsigned(1179, 12), 1925 => to_unsigned(3341, 12), 1926 => to_unsigned(3636, 12), 1927 => to_unsigned(635, 12), 1928 => to_unsigned(380, 12), 1929 => to_unsigned(1736, 12), 1930 => to_unsigned(861, 12), 1931 => to_unsigned(574, 12), 1932 => to_unsigned(1685, 12), 1933 => to_unsigned(1978, 12), 1934 => to_unsigned(563, 12), 1935 => to_unsigned(1257, 12), 1936 => to_unsigned(3943, 12), 1937 => to_unsigned(3073, 12), 1938 => to_unsigned(1065, 12), 1939 => to_unsigned(246, 12), 1940 => to_unsigned(2936, 12), 1941 => to_unsigned(1354, 12), 1942 => to_unsigned(454, 12), 1943 => to_unsigned(3651, 12), 1944 => to_unsigned(1551, 12), 1945 => to_unsigned(1001, 12), 1946 => to_unsigned(3440, 12), 1947 => to_unsigned(3522, 12), 1948 => to_unsigned(1332, 12), 1949 => to_unsigned(3801, 12), 1950 => to_unsigned(2112, 12), 1951 => to_unsigned(2090, 12), 1952 => to_unsigned(691, 12), 1953 => to_unsigned(3204, 12), 1954 => to_unsigned(1707, 12), 1955 => to_unsigned(2720, 12), 1956 => to_unsigned(528, 12), 1957 => to_unsigned(4094, 12), 1958 => to_unsigned(3086, 12), 1959 => to_unsigned(2649, 12), 1960 => to_unsigned(1238, 12), 1961 => to_unsigned(3438, 12), 1962 => to_unsigned(3453, 12), 1963 => to_unsigned(3988, 12), 1964 => to_unsigned(381, 12), 1965 => to_unsigned(697, 12), 1966 => to_unsigned(2715, 12), 1967 => to_unsigned(2307, 12), 1968 => to_unsigned(1206, 12), 1969 => to_unsigned(2613, 12), 1970 => to_unsigned(1297, 12), 1971 => to_unsigned(465, 12), 1972 => to_unsigned(2742, 12), 1973 => to_unsigned(517, 12), 1974 => to_unsigned(395, 12), 1975 => to_unsigned(3935, 12), 1976 => to_unsigned(2111, 12), 1977 => to_unsigned(5, 12), 1978 => to_unsigned(755, 12), 1979 => to_unsigned(2278, 12), 1980 => to_unsigned(36, 12), 1981 => to_unsigned(2353, 12), 1982 => to_unsigned(1620, 12), 1983 => to_unsigned(3980, 12), 1984 => to_unsigned(460, 12), 1985 => to_unsigned(2972, 12), 1986 => to_unsigned(2371, 12), 1987 => to_unsigned(1615, 12), 1988 => to_unsigned(318, 12), 1989 => to_unsigned(3133, 12), 1990 => to_unsigned(2984, 12), 1991 => to_unsigned(198, 12), 1992 => to_unsigned(315, 12), 1993 => to_unsigned(1368, 12), 1994 => to_unsigned(2363, 12), 1995 => to_unsigned(3898, 12), 1996 => to_unsigned(3418, 12), 1997 => to_unsigned(3682, 12), 1998 => to_unsigned(2961, 12), 1999 => to_unsigned(3910, 12), 2000 => to_unsigned(1623, 12), 2001 => to_unsigned(3299, 12), 2002 => to_unsigned(2830, 12), 2003 => to_unsigned(2167, 12), 2004 => to_unsigned(3526, 12), 2005 => to_unsigned(3364, 12), 2006 => to_unsigned(783, 12), 2007 => to_unsigned(3182, 12), 2008 => to_unsigned(1818, 12), 2009 => to_unsigned(2686, 12), 2010 => to_unsigned(2840, 12), 2011 => to_unsigned(3970, 12), 2012 => to_unsigned(1983, 12), 2013 => to_unsigned(2982, 12), 2014 => to_unsigned(3866, 12), 2015 => to_unsigned(458, 12), 2016 => to_unsigned(1790, 12), 2017 => to_unsigned(2479, 12), 2018 => to_unsigned(934, 12), 2019 => to_unsigned(4080, 12), 2020 => to_unsigned(2780, 12), 2021 => to_unsigned(84, 12), 2022 => to_unsigned(632, 12), 2023 => to_unsigned(2472, 12), 2024 => to_unsigned(3824, 12), 2025 => to_unsigned(248, 12), 2026 => to_unsigned(2971, 12), 2027 => to_unsigned(3997, 12), 2028 => to_unsigned(3731, 12), 2029 => to_unsigned(3689, 12), 2030 => to_unsigned(1304, 12), 2031 => to_unsigned(3414, 12), 2032 => to_unsigned(2315, 12), 2033 => to_unsigned(2891, 12), 2034 => to_unsigned(1066, 12), 2035 => to_unsigned(255, 12), 2036 => to_unsigned(1373, 12), 2037 => to_unsigned(960, 12), 2038 => to_unsigned(604, 12), 2039 => to_unsigned(1100, 12), 2040 => to_unsigned(2347, 12), 2041 => to_unsigned(3291, 12), 2042 => to_unsigned(605, 12), 2043 => to_unsigned(755, 12), 2044 => to_unsigned(1736, 12), 2045 => to_unsigned(895, 12), 2046 => to_unsigned(1437, 12), 2047 => to_unsigned(999, 12))
        ),
        2 => (
            0 => (0 => to_unsigned(3976, 12), 1 => to_unsigned(350, 12), 2 => to_unsigned(1255, 12), 3 => to_unsigned(1889, 12), 4 => to_unsigned(2699, 12), 5 => to_unsigned(324, 12), 6 => to_unsigned(2195, 12), 7 => to_unsigned(2927, 12), 8 => to_unsigned(3702, 12), 9 => to_unsigned(3445, 12), 10 => to_unsigned(1979, 12), 11 => to_unsigned(2218, 12), 12 => to_unsigned(1732, 12), 13 => to_unsigned(886, 12), 14 => to_unsigned(3826, 12), 15 => to_unsigned(3915, 12), 16 => to_unsigned(2391, 12), 17 => to_unsigned(2199, 12), 18 => to_unsigned(579, 12), 19 => to_unsigned(3892, 12), 20 => to_unsigned(210, 12), 21 => to_unsigned(1394, 12), 22 => to_unsigned(51, 12), 23 => to_unsigned(3023, 12), 24 => to_unsigned(2247, 12), 25 => to_unsigned(1348, 12), 26 => to_unsigned(2513, 12), 27 => to_unsigned(3999, 12), 28 => to_unsigned(2009, 12), 29 => to_unsigned(3113, 12), 30 => to_unsigned(3929, 12), 31 => to_unsigned(1830, 12), 32 => to_unsigned(3659, 12), 33 => to_unsigned(1467, 12), 34 => to_unsigned(879, 12), 35 => to_unsigned(2515, 12), 36 => to_unsigned(2799, 12), 37 => to_unsigned(3665, 12), 38 => to_unsigned(662, 12), 39 => to_unsigned(1416, 12), 40 => to_unsigned(3009, 12), 41 => to_unsigned(622, 12), 42 => to_unsigned(1033, 12), 43 => to_unsigned(3125, 12), 44 => to_unsigned(3907, 12), 45 => to_unsigned(165, 12), 46 => to_unsigned(3929, 12), 47 => to_unsigned(2780, 12), 48 => to_unsigned(3673, 12), 49 => to_unsigned(2670, 12), 50 => to_unsigned(1343, 12), 51 => to_unsigned(1389, 12), 52 => to_unsigned(767, 12), 53 => to_unsigned(1882, 12), 54 => to_unsigned(213, 12), 55 => to_unsigned(2719, 12), 56 => to_unsigned(1298, 12), 57 => to_unsigned(357, 12), 58 => to_unsigned(3561, 12), 59 => to_unsigned(1893, 12), 60 => to_unsigned(807, 12), 61 => to_unsigned(1994, 12), 62 => to_unsigned(662, 12), 63 => to_unsigned(1349, 12), 64 => to_unsigned(3908, 12), 65 => to_unsigned(97, 12), 66 => to_unsigned(505, 12), 67 => to_unsigned(2792, 12), 68 => to_unsigned(3562, 12), 69 => to_unsigned(3421, 12), 70 => to_unsigned(3372, 12), 71 => to_unsigned(1206, 12), 72 => to_unsigned(2196, 12), 73 => to_unsigned(1989, 12), 74 => to_unsigned(3194, 12), 75 => to_unsigned(111, 12), 76 => to_unsigned(2703, 12), 77 => to_unsigned(1904, 12), 78 => to_unsigned(2852, 12), 79 => to_unsigned(1053, 12), 80 => to_unsigned(245, 12), 81 => to_unsigned(1742, 12), 82 => to_unsigned(3311, 12), 83 => to_unsigned(3761, 12), 84 => to_unsigned(169, 12), 85 => to_unsigned(2164, 12), 86 => to_unsigned(1632, 12), 87 => to_unsigned(2800, 12), 88 => to_unsigned(730, 12), 89 => to_unsigned(870, 12), 90 => to_unsigned(2678, 12), 91 => to_unsigned(379, 12), 92 => to_unsigned(3776, 12), 93 => to_unsigned(2713, 12), 94 => to_unsigned(1050, 12), 95 => to_unsigned(1039, 12), 96 => to_unsigned(646, 12), 97 => to_unsigned(2340, 12), 98 => to_unsigned(237, 12), 99 => to_unsigned(3087, 12), 100 => to_unsigned(2311, 12), 101 => to_unsigned(3876, 12), 102 => to_unsigned(1223, 12), 103 => to_unsigned(2141, 12), 104 => to_unsigned(3832, 12), 105 => to_unsigned(1633, 12), 106 => to_unsigned(1606, 12), 107 => to_unsigned(1558, 12), 108 => to_unsigned(3097, 12), 109 => to_unsigned(1123, 12), 110 => to_unsigned(550, 12), 111 => to_unsigned(3657, 12), 112 => to_unsigned(2505, 12), 113 => to_unsigned(3392, 12), 114 => to_unsigned(2592, 12), 115 => to_unsigned(109, 12), 116 => to_unsigned(172, 12), 117 => to_unsigned(1701, 12), 118 => to_unsigned(2140, 12), 119 => to_unsigned(3402, 12), 120 => to_unsigned(1046, 12), 121 => to_unsigned(2248, 12), 122 => to_unsigned(2885, 12), 123 => to_unsigned(1489, 12), 124 => to_unsigned(1811, 12), 125 => to_unsigned(2104, 12), 126 => to_unsigned(2459, 12), 127 => to_unsigned(1586, 12), 128 => to_unsigned(1148, 12), 129 => to_unsigned(4052, 12), 130 => to_unsigned(1358, 12), 131 => to_unsigned(2774, 12), 132 => to_unsigned(4054, 12), 133 => to_unsigned(1933, 12), 134 => to_unsigned(1158, 12), 135 => to_unsigned(1662, 12), 136 => to_unsigned(3295, 12), 137 => to_unsigned(3487, 12), 138 => to_unsigned(264, 12), 139 => to_unsigned(202, 12), 140 => to_unsigned(3472, 12), 141 => to_unsigned(2245, 12), 142 => to_unsigned(2000, 12), 143 => to_unsigned(1402, 12), 144 => to_unsigned(2504, 12), 145 => to_unsigned(1866, 12), 146 => to_unsigned(2881, 12), 147 => to_unsigned(646, 12), 148 => to_unsigned(3724, 12), 149 => to_unsigned(3648, 12), 150 => to_unsigned(324, 12), 151 => to_unsigned(2495, 12), 152 => to_unsigned(3257, 12), 153 => to_unsigned(4029, 12), 154 => to_unsigned(2367, 12), 155 => to_unsigned(1189, 12), 156 => to_unsigned(4089, 12), 157 => to_unsigned(2306, 12), 158 => to_unsigned(506, 12), 159 => to_unsigned(1451, 12), 160 => to_unsigned(2527, 12), 161 => to_unsigned(2437, 12), 162 => to_unsigned(57, 12), 163 => to_unsigned(3474, 12), 164 => to_unsigned(1671, 12), 165 => to_unsigned(233, 12), 166 => to_unsigned(2146, 12), 167 => to_unsigned(2355, 12), 168 => to_unsigned(3277, 12), 169 => to_unsigned(3261, 12), 170 => to_unsigned(2102, 12), 171 => to_unsigned(3091, 12), 172 => to_unsigned(1763, 12), 173 => to_unsigned(3859, 12), 174 => to_unsigned(1490, 12), 175 => to_unsigned(761, 12), 176 => to_unsigned(2927, 12), 177 => to_unsigned(1002, 12), 178 => to_unsigned(3828, 12), 179 => to_unsigned(2015, 12), 180 => to_unsigned(2682, 12), 181 => to_unsigned(527, 12), 182 => to_unsigned(981, 12), 183 => to_unsigned(2865, 12), 184 => to_unsigned(3731, 12), 185 => to_unsigned(507, 12), 186 => to_unsigned(3774, 12), 187 => to_unsigned(3604, 12), 188 => to_unsigned(126, 12), 189 => to_unsigned(803, 12), 190 => to_unsigned(689, 12), 191 => to_unsigned(906, 12), 192 => to_unsigned(2925, 12), 193 => to_unsigned(1703, 12), 194 => to_unsigned(1036, 12), 195 => to_unsigned(397, 12), 196 => to_unsigned(3988, 12), 197 => to_unsigned(245, 12), 198 => to_unsigned(2238, 12), 199 => to_unsigned(3643, 12), 200 => to_unsigned(2226, 12), 201 => to_unsigned(1470, 12), 202 => to_unsigned(3909, 12), 203 => to_unsigned(3924, 12), 204 => to_unsigned(3899, 12), 205 => to_unsigned(2909, 12), 206 => to_unsigned(4013, 12), 207 => to_unsigned(2502, 12), 208 => to_unsigned(3258, 12), 209 => to_unsigned(3929, 12), 210 => to_unsigned(1444, 12), 211 => to_unsigned(685, 12), 212 => to_unsigned(3523, 12), 213 => to_unsigned(3349, 12), 214 => to_unsigned(1862, 12), 215 => to_unsigned(1862, 12), 216 => to_unsigned(860, 12), 217 => to_unsigned(553, 12), 218 => to_unsigned(934, 12), 219 => to_unsigned(904, 12), 220 => to_unsigned(1748, 12), 221 => to_unsigned(784, 12), 222 => to_unsigned(3571, 12), 223 => to_unsigned(2688, 12), 224 => to_unsigned(2797, 12), 225 => to_unsigned(2343, 12), 226 => to_unsigned(1643, 12), 227 => to_unsigned(453, 12), 228 => to_unsigned(3798, 12), 229 => to_unsigned(2510, 12), 230 => to_unsigned(678, 12), 231 => to_unsigned(1420, 12), 232 => to_unsigned(1261, 12), 233 => to_unsigned(3693, 12), 234 => to_unsigned(1743, 12), 235 => to_unsigned(2364, 12), 236 => to_unsigned(1967, 12), 237 => to_unsigned(3158, 12), 238 => to_unsigned(1283, 12), 239 => to_unsigned(3638, 12), 240 => to_unsigned(2111, 12), 241 => to_unsigned(914, 12), 242 => to_unsigned(2601, 12), 243 => to_unsigned(2571, 12), 244 => to_unsigned(2548, 12), 245 => to_unsigned(10, 12), 246 => to_unsigned(3217, 12), 247 => to_unsigned(4046, 12), 248 => to_unsigned(2745, 12), 249 => to_unsigned(2917, 12), 250 => to_unsigned(211, 12), 251 => to_unsigned(4060, 12), 252 => to_unsigned(3160, 12), 253 => to_unsigned(1850, 12), 254 => to_unsigned(3285, 12), 255 => to_unsigned(1001, 12), 256 => to_unsigned(3842, 12), 257 => to_unsigned(2860, 12), 258 => to_unsigned(1415, 12), 259 => to_unsigned(3818, 12), 260 => to_unsigned(2808, 12), 261 => to_unsigned(2042, 12), 262 => to_unsigned(3397, 12), 263 => to_unsigned(761, 12), 264 => to_unsigned(1895, 12), 265 => to_unsigned(3912, 12), 266 => to_unsigned(183, 12), 267 => to_unsigned(2733, 12), 268 => to_unsigned(1378, 12), 269 => to_unsigned(3724, 12), 270 => to_unsigned(2846, 12), 271 => to_unsigned(3394, 12), 272 => to_unsigned(3314, 12), 273 => to_unsigned(3282, 12), 274 => to_unsigned(3345, 12), 275 => to_unsigned(2555, 12), 276 => to_unsigned(1976, 12), 277 => to_unsigned(2247, 12), 278 => to_unsigned(4003, 12), 279 => to_unsigned(3468, 12), 280 => to_unsigned(3626, 12), 281 => to_unsigned(4089, 12), 282 => to_unsigned(2238, 12), 283 => to_unsigned(1428, 12), 284 => to_unsigned(1665, 12), 285 => to_unsigned(519, 12), 286 => to_unsigned(766, 12), 287 => to_unsigned(438, 12), 288 => to_unsigned(3791, 12), 289 => to_unsigned(1949, 12), 290 => to_unsigned(1277, 12), 291 => to_unsigned(3524, 12), 292 => to_unsigned(140, 12), 293 => to_unsigned(839, 12), 294 => to_unsigned(1095, 12), 295 => to_unsigned(3891, 12), 296 => to_unsigned(3570, 12), 297 => to_unsigned(2666, 12), 298 => to_unsigned(2956, 12), 299 => to_unsigned(3780, 12), 300 => to_unsigned(778, 12), 301 => to_unsigned(4092, 12), 302 => to_unsigned(447, 12), 303 => to_unsigned(2174, 12), 304 => to_unsigned(2299, 12), 305 => to_unsigned(1143, 12), 306 => to_unsigned(3387, 12), 307 => to_unsigned(735, 12), 308 => to_unsigned(2573, 12), 309 => to_unsigned(88, 12), 310 => to_unsigned(471, 12), 311 => to_unsigned(3195, 12), 312 => to_unsigned(2348, 12), 313 => to_unsigned(522, 12), 314 => to_unsigned(3285, 12), 315 => to_unsigned(2794, 12), 316 => to_unsigned(2024, 12), 317 => to_unsigned(1913, 12), 318 => to_unsigned(1266, 12), 319 => to_unsigned(902, 12), 320 => to_unsigned(4052, 12), 321 => to_unsigned(3628, 12), 322 => to_unsigned(2308, 12), 323 => to_unsigned(351, 12), 324 => to_unsigned(1887, 12), 325 => to_unsigned(3943, 12), 326 => to_unsigned(988, 12), 327 => to_unsigned(2064, 12), 328 => to_unsigned(577, 12), 329 => to_unsigned(3819, 12), 330 => to_unsigned(3040, 12), 331 => to_unsigned(1218, 12), 332 => to_unsigned(1143, 12), 333 => to_unsigned(1181, 12), 334 => to_unsigned(3402, 12), 335 => to_unsigned(2200, 12), 336 => to_unsigned(2824, 12), 337 => to_unsigned(3887, 12), 338 => to_unsigned(2142, 12), 339 => to_unsigned(1817, 12), 340 => to_unsigned(1545, 12), 341 => to_unsigned(2376, 12), 342 => to_unsigned(2812, 12), 343 => to_unsigned(3831, 12), 344 => to_unsigned(3267, 12), 345 => to_unsigned(170, 12), 346 => to_unsigned(1509, 12), 347 => to_unsigned(2317, 12), 348 => to_unsigned(31, 12), 349 => to_unsigned(2094, 12), 350 => to_unsigned(661, 12), 351 => to_unsigned(3456, 12), 352 => to_unsigned(3709, 12), 353 => to_unsigned(4035, 12), 354 => to_unsigned(2811, 12), 355 => to_unsigned(1850, 12), 356 => to_unsigned(838, 12), 357 => to_unsigned(460, 12), 358 => to_unsigned(3928, 12), 359 => to_unsigned(3454, 12), 360 => to_unsigned(309, 12), 361 => to_unsigned(1039, 12), 362 => to_unsigned(1924, 12), 363 => to_unsigned(3512, 12), 364 => to_unsigned(2441, 12), 365 => to_unsigned(3613, 12), 366 => to_unsigned(1053, 12), 367 => to_unsigned(538, 12), 368 => to_unsigned(3076, 12), 369 => to_unsigned(155, 12), 370 => to_unsigned(3613, 12), 371 => to_unsigned(2448, 12), 372 => to_unsigned(3184, 12), 373 => to_unsigned(1294, 12), 374 => to_unsigned(900, 12), 375 => to_unsigned(585, 12), 376 => to_unsigned(462, 12), 377 => to_unsigned(3339, 12), 378 => to_unsigned(1047, 12), 379 => to_unsigned(1778, 12), 380 => to_unsigned(1270, 12), 381 => to_unsigned(88, 12), 382 => to_unsigned(2197, 12), 383 => to_unsigned(3689, 12), 384 => to_unsigned(2241, 12), 385 => to_unsigned(2080, 12), 386 => to_unsigned(3788, 12), 387 => to_unsigned(3584, 12), 388 => to_unsigned(2527, 12), 389 => to_unsigned(36, 12), 390 => to_unsigned(667, 12), 391 => to_unsigned(3588, 12), 392 => to_unsigned(3644, 12), 393 => to_unsigned(4022, 12), 394 => to_unsigned(2159, 12), 395 => to_unsigned(2342, 12), 396 => to_unsigned(1458, 12), 397 => to_unsigned(3490, 12), 398 => to_unsigned(323, 12), 399 => to_unsigned(595, 12), 400 => to_unsigned(2406, 12), 401 => to_unsigned(4068, 12), 402 => to_unsigned(3637, 12), 403 => to_unsigned(2493, 12), 404 => to_unsigned(2929, 12), 405 => to_unsigned(3451, 12), 406 => to_unsigned(467, 12), 407 => to_unsigned(1796, 12), 408 => to_unsigned(1881, 12), 409 => to_unsigned(1365, 12), 410 => to_unsigned(3043, 12), 411 => to_unsigned(4004, 12), 412 => to_unsigned(3549, 12), 413 => to_unsigned(274, 12), 414 => to_unsigned(2305, 12), 415 => to_unsigned(955, 12), 416 => to_unsigned(154, 12), 417 => to_unsigned(2676, 12), 418 => to_unsigned(2333, 12), 419 => to_unsigned(2712, 12), 420 => to_unsigned(3126, 12), 421 => to_unsigned(2498, 12), 422 => to_unsigned(3121, 12), 423 => to_unsigned(1243, 12), 424 => to_unsigned(2738, 12), 425 => to_unsigned(2936, 12), 426 => to_unsigned(3949, 12), 427 => to_unsigned(1117, 12), 428 => to_unsigned(1146, 12), 429 => to_unsigned(331, 12), 430 => to_unsigned(566, 12), 431 => to_unsigned(1536, 12), 432 => to_unsigned(712, 12), 433 => to_unsigned(2267, 12), 434 => to_unsigned(2312, 12), 435 => to_unsigned(2726, 12), 436 => to_unsigned(746, 12), 437 => to_unsigned(1716, 12), 438 => to_unsigned(1360, 12), 439 => to_unsigned(1677, 12), 440 => to_unsigned(1720, 12), 441 => to_unsigned(1699, 12), 442 => to_unsigned(3227, 12), 443 => to_unsigned(23, 12), 444 => to_unsigned(943, 12), 445 => to_unsigned(3957, 12), 446 => to_unsigned(911, 12), 447 => to_unsigned(178, 12), 448 => to_unsigned(2936, 12), 449 => to_unsigned(3389, 12), 450 => to_unsigned(3720, 12), 451 => to_unsigned(1745, 12), 452 => to_unsigned(464, 12), 453 => to_unsigned(3992, 12), 454 => to_unsigned(3316, 12), 455 => to_unsigned(2615, 12), 456 => to_unsigned(270, 12), 457 => to_unsigned(1360, 12), 458 => to_unsigned(2888, 12), 459 => to_unsigned(2809, 12), 460 => to_unsigned(571, 12), 461 => to_unsigned(3159, 12), 462 => to_unsigned(2965, 12), 463 => to_unsigned(3274, 12), 464 => to_unsigned(929, 12), 465 => to_unsigned(1848, 12), 466 => to_unsigned(992, 12), 467 => to_unsigned(2597, 12), 468 => to_unsigned(2790, 12), 469 => to_unsigned(110, 12), 470 => to_unsigned(1999, 12), 471 => to_unsigned(1457, 12), 472 => to_unsigned(3689, 12), 473 => to_unsigned(3276, 12), 474 => to_unsigned(1202, 12), 475 => to_unsigned(3665, 12), 476 => to_unsigned(1483, 12), 477 => to_unsigned(2852, 12), 478 => to_unsigned(824, 12), 479 => to_unsigned(1178, 12), 480 => to_unsigned(730, 12), 481 => to_unsigned(3707, 12), 482 => to_unsigned(613, 12), 483 => to_unsigned(4009, 12), 484 => to_unsigned(3606, 12), 485 => to_unsigned(454, 12), 486 => to_unsigned(1684, 12), 487 => to_unsigned(1850, 12), 488 => to_unsigned(1419, 12), 489 => to_unsigned(3880, 12), 490 => to_unsigned(2241, 12), 491 => to_unsigned(1086, 12), 492 => to_unsigned(3353, 12), 493 => to_unsigned(456, 12), 494 => to_unsigned(3049, 12), 495 => to_unsigned(2244, 12), 496 => to_unsigned(2683, 12), 497 => to_unsigned(1151, 12), 498 => to_unsigned(3691, 12), 499 => to_unsigned(1594, 12), 500 => to_unsigned(2437, 12), 501 => to_unsigned(3906, 12), 502 => to_unsigned(692, 12), 503 => to_unsigned(727, 12), 504 => to_unsigned(1228, 12), 505 => to_unsigned(2490, 12), 506 => to_unsigned(1364, 12), 507 => to_unsigned(2744, 12), 508 => to_unsigned(2173, 12), 509 => to_unsigned(1085, 12), 510 => to_unsigned(1918, 12), 511 => to_unsigned(1320, 12), 512 => to_unsigned(237, 12), 513 => to_unsigned(1214, 12), 514 => to_unsigned(4043, 12), 515 => to_unsigned(2967, 12), 516 => to_unsigned(1920, 12), 517 => to_unsigned(1897, 12), 518 => to_unsigned(2803, 12), 519 => to_unsigned(346, 12), 520 => to_unsigned(3801, 12), 521 => to_unsigned(1188, 12), 522 => to_unsigned(430, 12), 523 => to_unsigned(1337, 12), 524 => to_unsigned(2047, 12), 525 => to_unsigned(541, 12), 526 => to_unsigned(3305, 12), 527 => to_unsigned(533, 12), 528 => to_unsigned(650, 12), 529 => to_unsigned(3575, 12), 530 => to_unsigned(1908, 12), 531 => to_unsigned(2000, 12), 532 => to_unsigned(1776, 12), 533 => to_unsigned(473, 12), 534 => to_unsigned(769, 12), 535 => to_unsigned(114, 12), 536 => to_unsigned(1389, 12), 537 => to_unsigned(2355, 12), 538 => to_unsigned(2218, 12), 539 => to_unsigned(649, 12), 540 => to_unsigned(1010, 12), 541 => to_unsigned(3142, 12), 542 => to_unsigned(1205, 12), 543 => to_unsigned(1094, 12), 544 => to_unsigned(267, 12), 545 => to_unsigned(3649, 12), 546 => to_unsigned(199, 12), 547 => to_unsigned(340, 12), 548 => to_unsigned(3177, 12), 549 => to_unsigned(2787, 12), 550 => to_unsigned(807, 12), 551 => to_unsigned(1518, 12), 552 => to_unsigned(642, 12), 553 => to_unsigned(547, 12), 554 => to_unsigned(129, 12), 555 => to_unsigned(2699, 12), 556 => to_unsigned(2960, 12), 557 => to_unsigned(2297, 12), 558 => to_unsigned(3038, 12), 559 => to_unsigned(1967, 12), 560 => to_unsigned(400, 12), 561 => to_unsigned(978, 12), 562 => to_unsigned(3819, 12), 563 => to_unsigned(3065, 12), 564 => to_unsigned(3557, 12), 565 => to_unsigned(331, 12), 566 => to_unsigned(3387, 12), 567 => to_unsigned(2777, 12), 568 => to_unsigned(2584, 12), 569 => to_unsigned(446, 12), 570 => to_unsigned(2281, 12), 571 => to_unsigned(107, 12), 572 => to_unsigned(1305, 12), 573 => to_unsigned(3290, 12), 574 => to_unsigned(3060, 12), 575 => to_unsigned(145, 12), 576 => to_unsigned(3113, 12), 577 => to_unsigned(1366, 12), 578 => to_unsigned(2958, 12), 579 => to_unsigned(3396, 12), 580 => to_unsigned(2579, 12), 581 => to_unsigned(2763, 12), 582 => to_unsigned(2655, 12), 583 => to_unsigned(2419, 12), 584 => to_unsigned(2804, 12), 585 => to_unsigned(133, 12), 586 => to_unsigned(1381, 12), 587 => to_unsigned(1781, 12), 588 => to_unsigned(816, 12), 589 => to_unsigned(451, 12), 590 => to_unsigned(2657, 12), 591 => to_unsigned(2545, 12), 592 => to_unsigned(622, 12), 593 => to_unsigned(760, 12), 594 => to_unsigned(497, 12), 595 => to_unsigned(2078, 12), 596 => to_unsigned(1410, 12), 597 => to_unsigned(3942, 12), 598 => to_unsigned(2359, 12), 599 => to_unsigned(3510, 12), 600 => to_unsigned(1079, 12), 601 => to_unsigned(1048, 12), 602 => to_unsigned(1527, 12), 603 => to_unsigned(1038, 12), 604 => to_unsigned(1793, 12), 605 => to_unsigned(4022, 12), 606 => to_unsigned(1204, 12), 607 => to_unsigned(2708, 12), 608 => to_unsigned(1685, 12), 609 => to_unsigned(1351, 12), 610 => to_unsigned(406, 12), 611 => to_unsigned(1113, 12), 612 => to_unsigned(2948, 12), 613 => to_unsigned(3579, 12), 614 => to_unsigned(1360, 12), 615 => to_unsigned(2549, 12), 616 => to_unsigned(2087, 12), 617 => to_unsigned(2582, 12), 618 => to_unsigned(1324, 12), 619 => to_unsigned(616, 12), 620 => to_unsigned(3688, 12), 621 => to_unsigned(3752, 12), 622 => to_unsigned(2625, 12), 623 => to_unsigned(4040, 12), 624 => to_unsigned(3187, 12), 625 => to_unsigned(42, 12), 626 => to_unsigned(245, 12), 627 => to_unsigned(2696, 12), 628 => to_unsigned(2487, 12), 629 => to_unsigned(455, 12), 630 => to_unsigned(1343, 12), 631 => to_unsigned(3612, 12), 632 => to_unsigned(616, 12), 633 => to_unsigned(2406, 12), 634 => to_unsigned(3588, 12), 635 => to_unsigned(3412, 12), 636 => to_unsigned(1635, 12), 637 => to_unsigned(1462, 12), 638 => to_unsigned(1515, 12), 639 => to_unsigned(628, 12), 640 => to_unsigned(3322, 12), 641 => to_unsigned(3911, 12), 642 => to_unsigned(937, 12), 643 => to_unsigned(3277, 12), 644 => to_unsigned(957, 12), 645 => to_unsigned(1592, 12), 646 => to_unsigned(1683, 12), 647 => to_unsigned(2080, 12), 648 => to_unsigned(2121, 12), 649 => to_unsigned(2142, 12), 650 => to_unsigned(1655, 12), 651 => to_unsigned(933, 12), 652 => to_unsigned(2156, 12), 653 => to_unsigned(3455, 12), 654 => to_unsigned(1869, 12), 655 => to_unsigned(1262, 12), 656 => to_unsigned(2398, 12), 657 => to_unsigned(2881, 12), 658 => to_unsigned(2636, 12), 659 => to_unsigned(2038, 12), 660 => to_unsigned(1156, 12), 661 => to_unsigned(2137, 12), 662 => to_unsigned(1386, 12), 663 => to_unsigned(27, 12), 664 => to_unsigned(2057, 12), 665 => to_unsigned(1096, 12), 666 => to_unsigned(445, 12), 667 => to_unsigned(3427, 12), 668 => to_unsigned(2456, 12), 669 => to_unsigned(481, 12), 670 => to_unsigned(1545, 12), 671 => to_unsigned(1407, 12), 672 => to_unsigned(1137, 12), 673 => to_unsigned(2628, 12), 674 => to_unsigned(3857, 12), 675 => to_unsigned(3058, 12), 676 => to_unsigned(490, 12), 677 => to_unsigned(3138, 12), 678 => to_unsigned(1941, 12), 679 => to_unsigned(2166, 12), 680 => to_unsigned(2315, 12), 681 => to_unsigned(3682, 12), 682 => to_unsigned(1820, 12), 683 => to_unsigned(2173, 12), 684 => to_unsigned(989, 12), 685 => to_unsigned(2531, 12), 686 => to_unsigned(2708, 12), 687 => to_unsigned(1091, 12), 688 => to_unsigned(2239, 12), 689 => to_unsigned(1950, 12), 690 => to_unsigned(1520, 12), 691 => to_unsigned(156, 12), 692 => to_unsigned(741, 12), 693 => to_unsigned(1498, 12), 694 => to_unsigned(1748, 12), 695 => to_unsigned(2083, 12), 696 => to_unsigned(3762, 12), 697 => to_unsigned(558, 12), 698 => to_unsigned(3155, 12), 699 => to_unsigned(3485, 12), 700 => to_unsigned(3810, 12), 701 => to_unsigned(1630, 12), 702 => to_unsigned(1072, 12), 703 => to_unsigned(284, 12), 704 => to_unsigned(3023, 12), 705 => to_unsigned(3236, 12), 706 => to_unsigned(625, 12), 707 => to_unsigned(1802, 12), 708 => to_unsigned(4037, 12), 709 => to_unsigned(3731, 12), 710 => to_unsigned(2178, 12), 711 => to_unsigned(1405, 12), 712 => to_unsigned(1265, 12), 713 => to_unsigned(1734, 12), 714 => to_unsigned(3008, 12), 715 => to_unsigned(1081, 12), 716 => to_unsigned(3230, 12), 717 => to_unsigned(2948, 12), 718 => to_unsigned(3584, 12), 719 => to_unsigned(1878, 12), 720 => to_unsigned(983, 12), 721 => to_unsigned(3082, 12), 722 => to_unsigned(3974, 12), 723 => to_unsigned(1982, 12), 724 => to_unsigned(2016, 12), 725 => to_unsigned(1347, 12), 726 => to_unsigned(548, 12), 727 => to_unsigned(1761, 12), 728 => to_unsigned(638, 12), 729 => to_unsigned(2272, 12), 730 => to_unsigned(3078, 12), 731 => to_unsigned(3781, 12), 732 => to_unsigned(101, 12), 733 => to_unsigned(3903, 12), 734 => to_unsigned(1103, 12), 735 => to_unsigned(2531, 12), 736 => to_unsigned(1881, 12), 737 => to_unsigned(19, 12), 738 => to_unsigned(1409, 12), 739 => to_unsigned(3051, 12), 740 => to_unsigned(2584, 12), 741 => to_unsigned(2678, 12), 742 => to_unsigned(2261, 12), 743 => to_unsigned(226, 12), 744 => to_unsigned(3726, 12), 745 => to_unsigned(2676, 12), 746 => to_unsigned(3458, 12), 747 => to_unsigned(3655, 12), 748 => to_unsigned(3173, 12), 749 => to_unsigned(3351, 12), 750 => to_unsigned(2742, 12), 751 => to_unsigned(422, 12), 752 => to_unsigned(2335, 12), 753 => to_unsigned(705, 12), 754 => to_unsigned(3071, 12), 755 => to_unsigned(2151, 12), 756 => to_unsigned(2491, 12), 757 => to_unsigned(1786, 12), 758 => to_unsigned(3089, 12), 759 => to_unsigned(2100, 12), 760 => to_unsigned(461, 12), 761 => to_unsigned(798, 12), 762 => to_unsigned(3939, 12), 763 => to_unsigned(313, 12), 764 => to_unsigned(2902, 12), 765 => to_unsigned(211, 12), 766 => to_unsigned(2299, 12), 767 => to_unsigned(1436, 12), 768 => to_unsigned(1350, 12), 769 => to_unsigned(3265, 12), 770 => to_unsigned(505, 12), 771 => to_unsigned(1029, 12), 772 => to_unsigned(1547, 12), 773 => to_unsigned(1077, 12), 774 => to_unsigned(3992, 12), 775 => to_unsigned(1370, 12), 776 => to_unsigned(760, 12), 777 => to_unsigned(1839, 12), 778 => to_unsigned(1345, 12), 779 => to_unsigned(1893, 12), 780 => to_unsigned(2730, 12), 781 => to_unsigned(3519, 12), 782 => to_unsigned(3232, 12), 783 => to_unsigned(2571, 12), 784 => to_unsigned(3986, 12), 785 => to_unsigned(639, 12), 786 => to_unsigned(3608, 12), 787 => to_unsigned(1156, 12), 788 => to_unsigned(3975, 12), 789 => to_unsigned(1568, 12), 790 => to_unsigned(399, 12), 791 => to_unsigned(2049, 12), 792 => to_unsigned(2417, 12), 793 => to_unsigned(2136, 12), 794 => to_unsigned(4005, 12), 795 => to_unsigned(2934, 12), 796 => to_unsigned(2641, 12), 797 => to_unsigned(372, 12), 798 => to_unsigned(2079, 12), 799 => to_unsigned(2975, 12), 800 => to_unsigned(456, 12), 801 => to_unsigned(4033, 12), 802 => to_unsigned(372, 12), 803 => to_unsigned(3825, 12), 804 => to_unsigned(2100, 12), 805 => to_unsigned(256, 12), 806 => to_unsigned(669, 12), 807 => to_unsigned(3896, 12), 808 => to_unsigned(897, 12), 809 => to_unsigned(153, 12), 810 => to_unsigned(3817, 12), 811 => to_unsigned(834, 12), 812 => to_unsigned(3116, 12), 813 => to_unsigned(2834, 12), 814 => to_unsigned(2772, 12), 815 => to_unsigned(3303, 12), 816 => to_unsigned(4065, 12), 817 => to_unsigned(3581, 12), 818 => to_unsigned(1843, 12), 819 => to_unsigned(3917, 12), 820 => to_unsigned(3359, 12), 821 => to_unsigned(2933, 12), 822 => to_unsigned(1156, 12), 823 => to_unsigned(3752, 12), 824 => to_unsigned(4067, 12), 825 => to_unsigned(3448, 12), 826 => to_unsigned(3191, 12), 827 => to_unsigned(1907, 12), 828 => to_unsigned(3682, 12), 829 => to_unsigned(3454, 12), 830 => to_unsigned(1431, 12), 831 => to_unsigned(2654, 12), 832 => to_unsigned(312, 12), 833 => to_unsigned(1465, 12), 834 => to_unsigned(2877, 12), 835 => to_unsigned(1027, 12), 836 => to_unsigned(333, 12), 837 => to_unsigned(1710, 12), 838 => to_unsigned(2331, 12), 839 => to_unsigned(3566, 12), 840 => to_unsigned(2144, 12), 841 => to_unsigned(1281, 12), 842 => to_unsigned(3075, 12), 843 => to_unsigned(1122, 12), 844 => to_unsigned(1764, 12), 845 => to_unsigned(2315, 12), 846 => to_unsigned(699, 12), 847 => to_unsigned(2151, 12), 848 => to_unsigned(1494, 12), 849 => to_unsigned(401, 12), 850 => to_unsigned(2204, 12), 851 => to_unsigned(2727, 12), 852 => to_unsigned(3138, 12), 853 => to_unsigned(820, 12), 854 => to_unsigned(3929, 12), 855 => to_unsigned(2704, 12), 856 => to_unsigned(3756, 12), 857 => to_unsigned(2671, 12), 858 => to_unsigned(1776, 12), 859 => to_unsigned(1142, 12), 860 => to_unsigned(1367, 12), 861 => to_unsigned(1269, 12), 862 => to_unsigned(1770, 12), 863 => to_unsigned(3204, 12), 864 => to_unsigned(1868, 12), 865 => to_unsigned(3527, 12), 866 => to_unsigned(1002, 12), 867 => to_unsigned(2583, 12), 868 => to_unsigned(2136, 12), 869 => to_unsigned(3519, 12), 870 => to_unsigned(1233, 12), 871 => to_unsigned(3828, 12), 872 => to_unsigned(2987, 12), 873 => to_unsigned(3804, 12), 874 => to_unsigned(453, 12), 875 => to_unsigned(1386, 12), 876 => to_unsigned(342, 12), 877 => to_unsigned(912, 12), 878 => to_unsigned(1839, 12), 879 => to_unsigned(4090, 12), 880 => to_unsigned(3689, 12), 881 => to_unsigned(1666, 12), 882 => to_unsigned(2757, 12), 883 => to_unsigned(683, 12), 884 => to_unsigned(2454, 12), 885 => to_unsigned(753, 12), 886 => to_unsigned(1299, 12), 887 => to_unsigned(1748, 12), 888 => to_unsigned(3622, 12), 889 => to_unsigned(1362, 12), 890 => to_unsigned(2697, 12), 891 => to_unsigned(2135, 12), 892 => to_unsigned(3907, 12), 893 => to_unsigned(430, 12), 894 => to_unsigned(134, 12), 895 => to_unsigned(1164, 12), 896 => to_unsigned(235, 12), 897 => to_unsigned(3209, 12), 898 => to_unsigned(1050, 12), 899 => to_unsigned(2029, 12), 900 => to_unsigned(457, 12), 901 => to_unsigned(2699, 12), 902 => to_unsigned(2501, 12), 903 => to_unsigned(256, 12), 904 => to_unsigned(1991, 12), 905 => to_unsigned(2486, 12), 906 => to_unsigned(829, 12), 907 => to_unsigned(3541, 12), 908 => to_unsigned(2761, 12), 909 => to_unsigned(2460, 12), 910 => to_unsigned(3152, 12), 911 => to_unsigned(46, 12), 912 => to_unsigned(1332, 12), 913 => to_unsigned(3028, 12), 914 => to_unsigned(1659, 12), 915 => to_unsigned(3880, 12), 916 => to_unsigned(885, 12), 917 => to_unsigned(1630, 12), 918 => to_unsigned(2574, 12), 919 => to_unsigned(1576, 12), 920 => to_unsigned(4052, 12), 921 => to_unsigned(1409, 12), 922 => to_unsigned(1708, 12), 923 => to_unsigned(1564, 12), 924 => to_unsigned(505, 12), 925 => to_unsigned(1419, 12), 926 => to_unsigned(3045, 12), 927 => to_unsigned(1725, 12), 928 => to_unsigned(507, 12), 929 => to_unsigned(1730, 12), 930 => to_unsigned(1313, 12), 931 => to_unsigned(3707, 12), 932 => to_unsigned(536, 12), 933 => to_unsigned(3332, 12), 934 => to_unsigned(2980, 12), 935 => to_unsigned(2226, 12), 936 => to_unsigned(3900, 12), 937 => to_unsigned(1116, 12), 938 => to_unsigned(2693, 12), 939 => to_unsigned(4061, 12), 940 => to_unsigned(3506, 12), 941 => to_unsigned(3671, 12), 942 => to_unsigned(3365, 12), 943 => to_unsigned(2567, 12), 944 => to_unsigned(3790, 12), 945 => to_unsigned(3168, 12), 946 => to_unsigned(1890, 12), 947 => to_unsigned(2669, 12), 948 => to_unsigned(707, 12), 949 => to_unsigned(1384, 12), 950 => to_unsigned(1990, 12), 951 => to_unsigned(1124, 12), 952 => to_unsigned(3820, 12), 953 => to_unsigned(2977, 12), 954 => to_unsigned(1470, 12), 955 => to_unsigned(1596, 12), 956 => to_unsigned(1268, 12), 957 => to_unsigned(2437, 12), 958 => to_unsigned(644, 12), 959 => to_unsigned(2411, 12), 960 => to_unsigned(3244, 12), 961 => to_unsigned(1940, 12), 962 => to_unsigned(34, 12), 963 => to_unsigned(1337, 12), 964 => to_unsigned(4091, 12), 965 => to_unsigned(3198, 12), 966 => to_unsigned(1376, 12), 967 => to_unsigned(1650, 12), 968 => to_unsigned(1175, 12), 969 => to_unsigned(340, 12), 970 => to_unsigned(1804, 12), 971 => to_unsigned(3573, 12), 972 => to_unsigned(1112, 12), 973 => to_unsigned(3214, 12), 974 => to_unsigned(1486, 12), 975 => to_unsigned(1402, 12), 976 => to_unsigned(2582, 12), 977 => to_unsigned(2182, 12), 978 => to_unsigned(3065, 12), 979 => to_unsigned(3940, 12), 980 => to_unsigned(2236, 12), 981 => to_unsigned(2557, 12), 982 => to_unsigned(1265, 12), 983 => to_unsigned(2806, 12), 984 => to_unsigned(3444, 12), 985 => to_unsigned(3884, 12), 986 => to_unsigned(1876, 12), 987 => to_unsigned(1643, 12), 988 => to_unsigned(648, 12), 989 => to_unsigned(3451, 12), 990 => to_unsigned(1339, 12), 991 => to_unsigned(1599, 12), 992 => to_unsigned(468, 12), 993 => to_unsigned(2248, 12), 994 => to_unsigned(2370, 12), 995 => to_unsigned(2851, 12), 996 => to_unsigned(2489, 12), 997 => to_unsigned(2509, 12), 998 => to_unsigned(233, 12), 999 => to_unsigned(1356, 12), 1000 => to_unsigned(3053, 12), 1001 => to_unsigned(2418, 12), 1002 => to_unsigned(825, 12), 1003 => to_unsigned(562, 12), 1004 => to_unsigned(278, 12), 1005 => to_unsigned(3204, 12), 1006 => to_unsigned(2090, 12), 1007 => to_unsigned(954, 12), 1008 => to_unsigned(1066, 12), 1009 => to_unsigned(3560, 12), 1010 => to_unsigned(1517, 12), 1011 => to_unsigned(2923, 12), 1012 => to_unsigned(1568, 12), 1013 => to_unsigned(1398, 12), 1014 => to_unsigned(965, 12), 1015 => to_unsigned(619, 12), 1016 => to_unsigned(2184, 12), 1017 => to_unsigned(704, 12), 1018 => to_unsigned(303, 12), 1019 => to_unsigned(1372, 12), 1020 => to_unsigned(695, 12), 1021 => to_unsigned(3928, 12), 1022 => to_unsigned(1940, 12), 1023 => to_unsigned(267, 12), 1024 => to_unsigned(3457, 12), 1025 => to_unsigned(601, 12), 1026 => to_unsigned(3383, 12), 1027 => to_unsigned(1903, 12), 1028 => to_unsigned(1061, 12), 1029 => to_unsigned(4000, 12), 1030 => to_unsigned(1329, 12), 1031 => to_unsigned(3147, 12), 1032 => to_unsigned(2373, 12), 1033 => to_unsigned(1424, 12), 1034 => to_unsigned(3880, 12), 1035 => to_unsigned(3980, 12), 1036 => to_unsigned(1520, 12), 1037 => to_unsigned(4055, 12), 1038 => to_unsigned(3307, 12), 1039 => to_unsigned(1625, 12), 1040 => to_unsigned(680, 12), 1041 => to_unsigned(1258, 12), 1042 => to_unsigned(833, 12), 1043 => to_unsigned(1241, 12), 1044 => to_unsigned(1942, 12), 1045 => to_unsigned(3393, 12), 1046 => to_unsigned(2231, 12), 1047 => to_unsigned(3405, 12), 1048 => to_unsigned(1173, 12), 1049 => to_unsigned(358, 12), 1050 => to_unsigned(1148, 12), 1051 => to_unsigned(1187, 12), 1052 => to_unsigned(1338, 12), 1053 => to_unsigned(608, 12), 1054 => to_unsigned(2191, 12), 1055 => to_unsigned(2678, 12), 1056 => to_unsigned(1735, 12), 1057 => to_unsigned(2743, 12), 1058 => to_unsigned(393, 12), 1059 => to_unsigned(4041, 12), 1060 => to_unsigned(2841, 12), 1061 => to_unsigned(3327, 12), 1062 => to_unsigned(754, 12), 1063 => to_unsigned(1755, 12), 1064 => to_unsigned(1717, 12), 1065 => to_unsigned(2008, 12), 1066 => to_unsigned(2786, 12), 1067 => to_unsigned(2477, 12), 1068 => to_unsigned(2968, 12), 1069 => to_unsigned(3919, 12), 1070 => to_unsigned(514, 12), 1071 => to_unsigned(2348, 12), 1072 => to_unsigned(1535, 12), 1073 => to_unsigned(2430, 12), 1074 => to_unsigned(772, 12), 1075 => to_unsigned(1415, 12), 1076 => to_unsigned(25, 12), 1077 => to_unsigned(4046, 12), 1078 => to_unsigned(925, 12), 1079 => to_unsigned(2389, 12), 1080 => to_unsigned(2380, 12), 1081 => to_unsigned(2706, 12), 1082 => to_unsigned(1526, 12), 1083 => to_unsigned(1776, 12), 1084 => to_unsigned(1518, 12), 1085 => to_unsigned(2571, 12), 1086 => to_unsigned(1893, 12), 1087 => to_unsigned(3083, 12), 1088 => to_unsigned(3585, 12), 1089 => to_unsigned(2255, 12), 1090 => to_unsigned(756, 12), 1091 => to_unsigned(1936, 12), 1092 => to_unsigned(2459, 12), 1093 => to_unsigned(717, 12), 1094 => to_unsigned(2727, 12), 1095 => to_unsigned(2591, 12), 1096 => to_unsigned(356, 12), 1097 => to_unsigned(3785, 12), 1098 => to_unsigned(2727, 12), 1099 => to_unsigned(209, 12), 1100 => to_unsigned(1838, 12), 1101 => to_unsigned(584, 12), 1102 => to_unsigned(548, 12), 1103 => to_unsigned(2338, 12), 1104 => to_unsigned(171, 12), 1105 => to_unsigned(3847, 12), 1106 => to_unsigned(122, 12), 1107 => to_unsigned(675, 12), 1108 => to_unsigned(1914, 12), 1109 => to_unsigned(2457, 12), 1110 => to_unsigned(3467, 12), 1111 => to_unsigned(1058, 12), 1112 => to_unsigned(2583, 12), 1113 => to_unsigned(2151, 12), 1114 => to_unsigned(2492, 12), 1115 => to_unsigned(2449, 12), 1116 => to_unsigned(3761, 12), 1117 => to_unsigned(1716, 12), 1118 => to_unsigned(981, 12), 1119 => to_unsigned(3546, 12), 1120 => to_unsigned(3182, 12), 1121 => to_unsigned(1786, 12), 1122 => to_unsigned(3275, 12), 1123 => to_unsigned(3961, 12), 1124 => to_unsigned(34, 12), 1125 => to_unsigned(246, 12), 1126 => to_unsigned(1154, 12), 1127 => to_unsigned(73, 12), 1128 => to_unsigned(2415, 12), 1129 => to_unsigned(1444, 12), 1130 => to_unsigned(3709, 12), 1131 => to_unsigned(2433, 12), 1132 => to_unsigned(1210, 12), 1133 => to_unsigned(3391, 12), 1134 => to_unsigned(3383, 12), 1135 => to_unsigned(3645, 12), 1136 => to_unsigned(3529, 12), 1137 => to_unsigned(3883, 12), 1138 => to_unsigned(2891, 12), 1139 => to_unsigned(2836, 12), 1140 => to_unsigned(3845, 12), 1141 => to_unsigned(2084, 12), 1142 => to_unsigned(3691, 12), 1143 => to_unsigned(1080, 12), 1144 => to_unsigned(4051, 12), 1145 => to_unsigned(2998, 12), 1146 => to_unsigned(2759, 12), 1147 => to_unsigned(1970, 12), 1148 => to_unsigned(2874, 12), 1149 => to_unsigned(931, 12), 1150 => to_unsigned(1030, 12), 1151 => to_unsigned(545, 12), 1152 => to_unsigned(216, 12), 1153 => to_unsigned(259, 12), 1154 => to_unsigned(2777, 12), 1155 => to_unsigned(657, 12), 1156 => to_unsigned(2792, 12), 1157 => to_unsigned(2991, 12), 1158 => to_unsigned(1612, 12), 1159 => to_unsigned(3052, 12), 1160 => to_unsigned(1775, 12), 1161 => to_unsigned(305, 12), 1162 => to_unsigned(1589, 12), 1163 => to_unsigned(3595, 12), 1164 => to_unsigned(1672, 12), 1165 => to_unsigned(3062, 12), 1166 => to_unsigned(733, 12), 1167 => to_unsigned(2865, 12), 1168 => to_unsigned(536, 12), 1169 => to_unsigned(3740, 12), 1170 => to_unsigned(2336, 12), 1171 => to_unsigned(3411, 12), 1172 => to_unsigned(3374, 12), 1173 => to_unsigned(1864, 12), 1174 => to_unsigned(1912, 12), 1175 => to_unsigned(3417, 12), 1176 => to_unsigned(1168, 12), 1177 => to_unsigned(3532, 12), 1178 => to_unsigned(3318, 12), 1179 => to_unsigned(1390, 12), 1180 => to_unsigned(1187, 12), 1181 => to_unsigned(2942, 12), 1182 => to_unsigned(3307, 12), 1183 => to_unsigned(2174, 12), 1184 => to_unsigned(3687, 12), 1185 => to_unsigned(1336, 12), 1186 => to_unsigned(2595, 12), 1187 => to_unsigned(29, 12), 1188 => to_unsigned(2894, 12), 1189 => to_unsigned(717, 12), 1190 => to_unsigned(1133, 12), 1191 => to_unsigned(2442, 12), 1192 => to_unsigned(2960, 12), 1193 => to_unsigned(1411, 12), 1194 => to_unsigned(3839, 12), 1195 => to_unsigned(3349, 12), 1196 => to_unsigned(1566, 12), 1197 => to_unsigned(1691, 12), 1198 => to_unsigned(3687, 12), 1199 => to_unsigned(650, 12), 1200 => to_unsigned(311, 12), 1201 => to_unsigned(3936, 12), 1202 => to_unsigned(1289, 12), 1203 => to_unsigned(1498, 12), 1204 => to_unsigned(2653, 12), 1205 => to_unsigned(1007, 12), 1206 => to_unsigned(2939, 12), 1207 => to_unsigned(3507, 12), 1208 => to_unsigned(2068, 12), 1209 => to_unsigned(1948, 12), 1210 => to_unsigned(2606, 12), 1211 => to_unsigned(887, 12), 1212 => to_unsigned(1944, 12), 1213 => to_unsigned(1824, 12), 1214 => to_unsigned(2955, 12), 1215 => to_unsigned(63, 12), 1216 => to_unsigned(3268, 12), 1217 => to_unsigned(1547, 12), 1218 => to_unsigned(539, 12), 1219 => to_unsigned(3240, 12), 1220 => to_unsigned(1805, 12), 1221 => to_unsigned(3838, 12), 1222 => to_unsigned(3130, 12), 1223 => to_unsigned(2176, 12), 1224 => to_unsigned(2212, 12), 1225 => to_unsigned(1828, 12), 1226 => to_unsigned(2123, 12), 1227 => to_unsigned(661, 12), 1228 => to_unsigned(3446, 12), 1229 => to_unsigned(1484, 12), 1230 => to_unsigned(1757, 12), 1231 => to_unsigned(1206, 12), 1232 => to_unsigned(1774, 12), 1233 => to_unsigned(3062, 12), 1234 => to_unsigned(3032, 12), 1235 => to_unsigned(1674, 12), 1236 => to_unsigned(2711, 12), 1237 => to_unsigned(770, 12), 1238 => to_unsigned(2655, 12), 1239 => to_unsigned(358, 12), 1240 => to_unsigned(3548, 12), 1241 => to_unsigned(699, 12), 1242 => to_unsigned(804, 12), 1243 => to_unsigned(1399, 12), 1244 => to_unsigned(2092, 12), 1245 => to_unsigned(3884, 12), 1246 => to_unsigned(3414, 12), 1247 => to_unsigned(964, 12), 1248 => to_unsigned(3400, 12), 1249 => to_unsigned(3974, 12), 1250 => to_unsigned(3662, 12), 1251 => to_unsigned(148, 12), 1252 => to_unsigned(440, 12), 1253 => to_unsigned(3906, 12), 1254 => to_unsigned(1619, 12), 1255 => to_unsigned(371, 12), 1256 => to_unsigned(1069, 12), 1257 => to_unsigned(2628, 12), 1258 => to_unsigned(1279, 12), 1259 => to_unsigned(1862, 12), 1260 => to_unsigned(696, 12), 1261 => to_unsigned(1128, 12), 1262 => to_unsigned(3924, 12), 1263 => to_unsigned(1592, 12), 1264 => to_unsigned(673, 12), 1265 => to_unsigned(1433, 12), 1266 => to_unsigned(2688, 12), 1267 => to_unsigned(3977, 12), 1268 => to_unsigned(1114, 12), 1269 => to_unsigned(3029, 12), 1270 => to_unsigned(3789, 12), 1271 => to_unsigned(976, 12), 1272 => to_unsigned(409, 12), 1273 => to_unsigned(3978, 12), 1274 => to_unsigned(891, 12), 1275 => to_unsigned(1979, 12), 1276 => to_unsigned(2879, 12), 1277 => to_unsigned(261, 12), 1278 => to_unsigned(138, 12), 1279 => to_unsigned(3996, 12), 1280 => to_unsigned(914, 12), 1281 => to_unsigned(2155, 12), 1282 => to_unsigned(1726, 12), 1283 => to_unsigned(3733, 12), 1284 => to_unsigned(1850, 12), 1285 => to_unsigned(687, 12), 1286 => to_unsigned(2404, 12), 1287 => to_unsigned(2639, 12), 1288 => to_unsigned(2498, 12), 1289 => to_unsigned(1913, 12), 1290 => to_unsigned(1481, 12), 1291 => to_unsigned(1081, 12), 1292 => to_unsigned(3987, 12), 1293 => to_unsigned(2152, 12), 1294 => to_unsigned(1721, 12), 1295 => to_unsigned(1511, 12), 1296 => to_unsigned(2354, 12), 1297 => to_unsigned(1774, 12), 1298 => to_unsigned(669, 12), 1299 => to_unsigned(1799, 12), 1300 => to_unsigned(523, 12), 1301 => to_unsigned(1623, 12), 1302 => to_unsigned(2422, 12), 1303 => to_unsigned(2120, 12), 1304 => to_unsigned(3735, 12), 1305 => to_unsigned(3908, 12), 1306 => to_unsigned(3456, 12), 1307 => to_unsigned(3354, 12), 1308 => to_unsigned(1525, 12), 1309 => to_unsigned(3412, 12), 1310 => to_unsigned(2752, 12), 1311 => to_unsigned(3409, 12), 1312 => to_unsigned(3295, 12), 1313 => to_unsigned(4020, 12), 1314 => to_unsigned(2757, 12), 1315 => to_unsigned(3847, 12), 1316 => to_unsigned(3045, 12), 1317 => to_unsigned(2551, 12), 1318 => to_unsigned(2341, 12), 1319 => to_unsigned(1044, 12), 1320 => to_unsigned(620, 12), 1321 => to_unsigned(361, 12), 1322 => to_unsigned(84, 12), 1323 => to_unsigned(1182, 12), 1324 => to_unsigned(2447, 12), 1325 => to_unsigned(1958, 12), 1326 => to_unsigned(2204, 12), 1327 => to_unsigned(3377, 12), 1328 => to_unsigned(2645, 12), 1329 => to_unsigned(3566, 12), 1330 => to_unsigned(2009, 12), 1331 => to_unsigned(2959, 12), 1332 => to_unsigned(432, 12), 1333 => to_unsigned(3171, 12), 1334 => to_unsigned(2316, 12), 1335 => to_unsigned(3704, 12), 1336 => to_unsigned(3095, 12), 1337 => to_unsigned(1896, 12), 1338 => to_unsigned(3749, 12), 1339 => to_unsigned(3440, 12), 1340 => to_unsigned(3275, 12), 1341 => to_unsigned(2513, 12), 1342 => to_unsigned(472, 12), 1343 => to_unsigned(3468, 12), 1344 => to_unsigned(3575, 12), 1345 => to_unsigned(2474, 12), 1346 => to_unsigned(3644, 12), 1347 => to_unsigned(2459, 12), 1348 => to_unsigned(2016, 12), 1349 => to_unsigned(1926, 12), 1350 => to_unsigned(826, 12), 1351 => to_unsigned(3702, 12), 1352 => to_unsigned(813, 12), 1353 => to_unsigned(1644, 12), 1354 => to_unsigned(2792, 12), 1355 => to_unsigned(4073, 12), 1356 => to_unsigned(1430, 12), 1357 => to_unsigned(3212, 12), 1358 => to_unsigned(341, 12), 1359 => to_unsigned(3456, 12), 1360 => to_unsigned(874, 12), 1361 => to_unsigned(1180, 12), 1362 => to_unsigned(555, 12), 1363 => to_unsigned(3811, 12), 1364 => to_unsigned(4080, 12), 1365 => to_unsigned(2497, 12), 1366 => to_unsigned(3729, 12), 1367 => to_unsigned(3447, 12), 1368 => to_unsigned(3097, 12), 1369 => to_unsigned(1423, 12), 1370 => to_unsigned(717, 12), 1371 => to_unsigned(1143, 12), 1372 => to_unsigned(127, 12), 1373 => to_unsigned(3349, 12), 1374 => to_unsigned(1026, 12), 1375 => to_unsigned(3558, 12), 1376 => to_unsigned(1678, 12), 1377 => to_unsigned(2068, 12), 1378 => to_unsigned(881, 12), 1379 => to_unsigned(1559, 12), 1380 => to_unsigned(2082, 12), 1381 => to_unsigned(3686, 12), 1382 => to_unsigned(3318, 12), 1383 => to_unsigned(3400, 12), 1384 => to_unsigned(2838, 12), 1385 => to_unsigned(7, 12), 1386 => to_unsigned(1844, 12), 1387 => to_unsigned(3307, 12), 1388 => to_unsigned(2879, 12), 1389 => to_unsigned(3073, 12), 1390 => to_unsigned(968, 12), 1391 => to_unsigned(2460, 12), 1392 => to_unsigned(2011, 12), 1393 => to_unsigned(1250, 12), 1394 => to_unsigned(1181, 12), 1395 => to_unsigned(3002, 12), 1396 => to_unsigned(1246, 12), 1397 => to_unsigned(2953, 12), 1398 => to_unsigned(2108, 12), 1399 => to_unsigned(3920, 12), 1400 => to_unsigned(2038, 12), 1401 => to_unsigned(1655, 12), 1402 => to_unsigned(1256, 12), 1403 => to_unsigned(2461, 12), 1404 => to_unsigned(1200, 12), 1405 => to_unsigned(857, 12), 1406 => to_unsigned(3041, 12), 1407 => to_unsigned(2369, 12), 1408 => to_unsigned(2977, 12), 1409 => to_unsigned(2002, 12), 1410 => to_unsigned(2332, 12), 1411 => to_unsigned(1840, 12), 1412 => to_unsigned(2795, 12), 1413 => to_unsigned(3688, 12), 1414 => to_unsigned(3637, 12), 1415 => to_unsigned(850, 12), 1416 => to_unsigned(326, 12), 1417 => to_unsigned(2595, 12), 1418 => to_unsigned(3945, 12), 1419 => to_unsigned(393, 12), 1420 => to_unsigned(2328, 12), 1421 => to_unsigned(1922, 12), 1422 => to_unsigned(1051, 12), 1423 => to_unsigned(880, 12), 1424 => to_unsigned(1214, 12), 1425 => to_unsigned(3650, 12), 1426 => to_unsigned(79, 12), 1427 => to_unsigned(642, 12), 1428 => to_unsigned(1611, 12), 1429 => to_unsigned(3867, 12), 1430 => to_unsigned(995, 12), 1431 => to_unsigned(111, 12), 1432 => to_unsigned(1902, 12), 1433 => to_unsigned(271, 12), 1434 => to_unsigned(36, 12), 1435 => to_unsigned(2391, 12), 1436 => to_unsigned(1933, 12), 1437 => to_unsigned(3378, 12), 1438 => to_unsigned(1353, 12), 1439 => to_unsigned(2107, 12), 1440 => to_unsigned(3708, 12), 1441 => to_unsigned(3731, 12), 1442 => to_unsigned(1622, 12), 1443 => to_unsigned(1782, 12), 1444 => to_unsigned(2149, 12), 1445 => to_unsigned(3492, 12), 1446 => to_unsigned(1852, 12), 1447 => to_unsigned(1679, 12), 1448 => to_unsigned(937, 12), 1449 => to_unsigned(2235, 12), 1450 => to_unsigned(2142, 12), 1451 => to_unsigned(525, 12), 1452 => to_unsigned(4074, 12), 1453 => to_unsigned(3652, 12), 1454 => to_unsigned(1602, 12), 1455 => to_unsigned(278, 12), 1456 => to_unsigned(3542, 12), 1457 => to_unsigned(1995, 12), 1458 => to_unsigned(892, 12), 1459 => to_unsigned(3670, 12), 1460 => to_unsigned(2653, 12), 1461 => to_unsigned(1444, 12), 1462 => to_unsigned(3170, 12), 1463 => to_unsigned(480, 12), 1464 => to_unsigned(2656, 12), 1465 => to_unsigned(2968, 12), 1466 => to_unsigned(3896, 12), 1467 => to_unsigned(922, 12), 1468 => to_unsigned(1303, 12), 1469 => to_unsigned(1128, 12), 1470 => to_unsigned(1398, 12), 1471 => to_unsigned(3828, 12), 1472 => to_unsigned(722, 12), 1473 => to_unsigned(2883, 12), 1474 => to_unsigned(2008, 12), 1475 => to_unsigned(3410, 12), 1476 => to_unsigned(3701, 12), 1477 => to_unsigned(25, 12), 1478 => to_unsigned(1823, 12), 1479 => to_unsigned(1464, 12), 1480 => to_unsigned(553, 12), 1481 => to_unsigned(2316, 12), 1482 => to_unsigned(1586, 12), 1483 => to_unsigned(1823, 12), 1484 => to_unsigned(3232, 12), 1485 => to_unsigned(2095, 12), 1486 => to_unsigned(3336, 12), 1487 => to_unsigned(2951, 12), 1488 => to_unsigned(105, 12), 1489 => to_unsigned(3445, 12), 1490 => to_unsigned(1690, 12), 1491 => to_unsigned(2638, 12), 1492 => to_unsigned(2270, 12), 1493 => to_unsigned(40, 12), 1494 => to_unsigned(1710, 12), 1495 => to_unsigned(1674, 12), 1496 => to_unsigned(843, 12), 1497 => to_unsigned(1150, 12), 1498 => to_unsigned(1992, 12), 1499 => to_unsigned(4015, 12), 1500 => to_unsigned(1425, 12), 1501 => to_unsigned(3617, 12), 1502 => to_unsigned(3107, 12), 1503 => to_unsigned(2686, 12), 1504 => to_unsigned(928, 12), 1505 => to_unsigned(3827, 12), 1506 => to_unsigned(945, 12), 1507 => to_unsigned(1930, 12), 1508 => to_unsigned(3918, 12), 1509 => to_unsigned(3716, 12), 1510 => to_unsigned(2678, 12), 1511 => to_unsigned(1984, 12), 1512 => to_unsigned(2853, 12), 1513 => to_unsigned(2338, 12), 1514 => to_unsigned(1077, 12), 1515 => to_unsigned(2644, 12), 1516 => to_unsigned(3013, 12), 1517 => to_unsigned(3710, 12), 1518 => to_unsigned(2447, 12), 1519 => to_unsigned(3597, 12), 1520 => to_unsigned(710, 12), 1521 => to_unsigned(1644, 12), 1522 => to_unsigned(3567, 12), 1523 => to_unsigned(302, 12), 1524 => to_unsigned(2162, 12), 1525 => to_unsigned(764, 12), 1526 => to_unsigned(3267, 12), 1527 => to_unsigned(2536, 12), 1528 => to_unsigned(2293, 12), 1529 => to_unsigned(172, 12), 1530 => to_unsigned(2099, 12), 1531 => to_unsigned(2829, 12), 1532 => to_unsigned(781, 12), 1533 => to_unsigned(2439, 12), 1534 => to_unsigned(2522, 12), 1535 => to_unsigned(1714, 12), 1536 => to_unsigned(2912, 12), 1537 => to_unsigned(3942, 12), 1538 => to_unsigned(3866, 12), 1539 => to_unsigned(1356, 12), 1540 => to_unsigned(2863, 12), 1541 => to_unsigned(3183, 12), 1542 => to_unsigned(3313, 12), 1543 => to_unsigned(3773, 12), 1544 => to_unsigned(2455, 12), 1545 => to_unsigned(3074, 12), 1546 => to_unsigned(2483, 12), 1547 => to_unsigned(2003, 12), 1548 => to_unsigned(2259, 12), 1549 => to_unsigned(2779, 12), 1550 => to_unsigned(3209, 12), 1551 => to_unsigned(3492, 12), 1552 => to_unsigned(978, 12), 1553 => to_unsigned(288, 12), 1554 => to_unsigned(3985, 12), 1555 => to_unsigned(1413, 12), 1556 => to_unsigned(1694, 12), 1557 => to_unsigned(3230, 12), 1558 => to_unsigned(1017, 12), 1559 => to_unsigned(1845, 12), 1560 => to_unsigned(2817, 12), 1561 => to_unsigned(1146, 12), 1562 => to_unsigned(2492, 12), 1563 => to_unsigned(73, 12), 1564 => to_unsigned(2530, 12), 1565 => to_unsigned(3724, 12), 1566 => to_unsigned(3769, 12), 1567 => to_unsigned(694, 12), 1568 => to_unsigned(1662, 12), 1569 => to_unsigned(3272, 12), 1570 => to_unsigned(1062, 12), 1571 => to_unsigned(1079, 12), 1572 => to_unsigned(2622, 12), 1573 => to_unsigned(4058, 12), 1574 => to_unsigned(3388, 12), 1575 => to_unsigned(3467, 12), 1576 => to_unsigned(4083, 12), 1577 => to_unsigned(2865, 12), 1578 => to_unsigned(893, 12), 1579 => to_unsigned(3524, 12), 1580 => to_unsigned(2181, 12), 1581 => to_unsigned(2349, 12), 1582 => to_unsigned(289, 12), 1583 => to_unsigned(3828, 12), 1584 => to_unsigned(2904, 12), 1585 => to_unsigned(4044, 12), 1586 => to_unsigned(1885, 12), 1587 => to_unsigned(1216, 12), 1588 => to_unsigned(3291, 12), 1589 => to_unsigned(1093, 12), 1590 => to_unsigned(1000, 12), 1591 => to_unsigned(429, 12), 1592 => to_unsigned(850, 12), 1593 => to_unsigned(3762, 12), 1594 => to_unsigned(3106, 12), 1595 => to_unsigned(2554, 12), 1596 => to_unsigned(2111, 12), 1597 => to_unsigned(3601, 12), 1598 => to_unsigned(909, 12), 1599 => to_unsigned(2133, 12), 1600 => to_unsigned(3557, 12), 1601 => to_unsigned(970, 12), 1602 => to_unsigned(3651, 12), 1603 => to_unsigned(3985, 12), 1604 => to_unsigned(122, 12), 1605 => to_unsigned(1202, 12), 1606 => to_unsigned(2275, 12), 1607 => to_unsigned(588, 12), 1608 => to_unsigned(3439, 12), 1609 => to_unsigned(1200, 12), 1610 => to_unsigned(3522, 12), 1611 => to_unsigned(2705, 12), 1612 => to_unsigned(2588, 12), 1613 => to_unsigned(2320, 12), 1614 => to_unsigned(2052, 12), 1615 => to_unsigned(3104, 12), 1616 => to_unsigned(2737, 12), 1617 => to_unsigned(81, 12), 1618 => to_unsigned(1991, 12), 1619 => to_unsigned(1042, 12), 1620 => to_unsigned(312, 12), 1621 => to_unsigned(1094, 12), 1622 => to_unsigned(1986, 12), 1623 => to_unsigned(1592, 12), 1624 => to_unsigned(3538, 12), 1625 => to_unsigned(870, 12), 1626 => to_unsigned(824, 12), 1627 => to_unsigned(1680, 12), 1628 => to_unsigned(742, 12), 1629 => to_unsigned(3223, 12), 1630 => to_unsigned(1817, 12), 1631 => to_unsigned(3894, 12), 1632 => to_unsigned(556, 12), 1633 => to_unsigned(3956, 12), 1634 => to_unsigned(3159, 12), 1635 => to_unsigned(2387, 12), 1636 => to_unsigned(684, 12), 1637 => to_unsigned(1951, 12), 1638 => to_unsigned(2142, 12), 1639 => to_unsigned(1985, 12), 1640 => to_unsigned(3169, 12), 1641 => to_unsigned(2072, 12), 1642 => to_unsigned(982, 12), 1643 => to_unsigned(4001, 12), 1644 => to_unsigned(723, 12), 1645 => to_unsigned(1950, 12), 1646 => to_unsigned(4093, 12), 1647 => to_unsigned(602, 12), 1648 => to_unsigned(2594, 12), 1649 => to_unsigned(3028, 12), 1650 => to_unsigned(1008, 12), 1651 => to_unsigned(740, 12), 1652 => to_unsigned(81, 12), 1653 => to_unsigned(3600, 12), 1654 => to_unsigned(2351, 12), 1655 => to_unsigned(2874, 12), 1656 => to_unsigned(2779, 12), 1657 => to_unsigned(1881, 12), 1658 => to_unsigned(2722, 12), 1659 => to_unsigned(3299, 12), 1660 => to_unsigned(1531, 12), 1661 => to_unsigned(1894, 12), 1662 => to_unsigned(2438, 12), 1663 => to_unsigned(30, 12), 1664 => to_unsigned(824, 12), 1665 => to_unsigned(849, 12), 1666 => to_unsigned(3917, 12), 1667 => to_unsigned(3376, 12), 1668 => to_unsigned(4020, 12), 1669 => to_unsigned(493, 12), 1670 => to_unsigned(2427, 12), 1671 => to_unsigned(3701, 12), 1672 => to_unsigned(2178, 12), 1673 => to_unsigned(1050, 12), 1674 => to_unsigned(2684, 12), 1675 => to_unsigned(2999, 12), 1676 => to_unsigned(152, 12), 1677 => to_unsigned(4079, 12), 1678 => to_unsigned(3356, 12), 1679 => to_unsigned(968, 12), 1680 => to_unsigned(3575, 12), 1681 => to_unsigned(1252, 12), 1682 => to_unsigned(1228, 12), 1683 => to_unsigned(1061, 12), 1684 => to_unsigned(895, 12), 1685 => to_unsigned(1001, 12), 1686 => to_unsigned(4037, 12), 1687 => to_unsigned(1153, 12), 1688 => to_unsigned(2281, 12), 1689 => to_unsigned(808, 12), 1690 => to_unsigned(2386, 12), 1691 => to_unsigned(1272, 12), 1692 => to_unsigned(2218, 12), 1693 => to_unsigned(3413, 12), 1694 => to_unsigned(2112, 12), 1695 => to_unsigned(1360, 12), 1696 => to_unsigned(681, 12), 1697 => to_unsigned(2284, 12), 1698 => to_unsigned(39, 12), 1699 => to_unsigned(3295, 12), 1700 => to_unsigned(2661, 12), 1701 => to_unsigned(3180, 12), 1702 => to_unsigned(2520, 12), 1703 => to_unsigned(1139, 12), 1704 => to_unsigned(1563, 12), 1705 => to_unsigned(2917, 12), 1706 => to_unsigned(3661, 12), 1707 => to_unsigned(2716, 12), 1708 => to_unsigned(58, 12), 1709 => to_unsigned(3041, 12), 1710 => to_unsigned(1985, 12), 1711 => to_unsigned(1558, 12), 1712 => to_unsigned(3149, 12), 1713 => to_unsigned(2318, 12), 1714 => to_unsigned(996, 12), 1715 => to_unsigned(3161, 12), 1716 => to_unsigned(3488, 12), 1717 => to_unsigned(2246, 12), 1718 => to_unsigned(2321, 12), 1719 => to_unsigned(1063, 12), 1720 => to_unsigned(1028, 12), 1721 => to_unsigned(3700, 12), 1722 => to_unsigned(3226, 12), 1723 => to_unsigned(94, 12), 1724 => to_unsigned(3208, 12), 1725 => to_unsigned(3214, 12), 1726 => to_unsigned(3256, 12), 1727 => to_unsigned(3162, 12), 1728 => to_unsigned(2833, 12), 1729 => to_unsigned(4052, 12), 1730 => to_unsigned(2076, 12), 1731 => to_unsigned(811, 12), 1732 => to_unsigned(259, 12), 1733 => to_unsigned(3520, 12), 1734 => to_unsigned(1036, 12), 1735 => to_unsigned(1619, 12), 1736 => to_unsigned(2110, 12), 1737 => to_unsigned(1662, 12), 1738 => to_unsigned(1591, 12), 1739 => to_unsigned(1727, 12), 1740 => to_unsigned(442, 12), 1741 => to_unsigned(1364, 12), 1742 => to_unsigned(2569, 12), 1743 => to_unsigned(2984, 12), 1744 => to_unsigned(1841, 12), 1745 => to_unsigned(195, 12), 1746 => to_unsigned(1631, 12), 1747 => to_unsigned(1293, 12), 1748 => to_unsigned(3180, 12), 1749 => to_unsigned(1367, 12), 1750 => to_unsigned(3346, 12), 1751 => to_unsigned(255, 12), 1752 => to_unsigned(2620, 12), 1753 => to_unsigned(327, 12), 1754 => to_unsigned(1708, 12), 1755 => to_unsigned(3504, 12), 1756 => to_unsigned(2859, 12), 1757 => to_unsigned(4054, 12), 1758 => to_unsigned(2537, 12), 1759 => to_unsigned(1719, 12), 1760 => to_unsigned(683, 12), 1761 => to_unsigned(52, 12), 1762 => to_unsigned(181, 12), 1763 => to_unsigned(2454, 12), 1764 => to_unsigned(1346, 12), 1765 => to_unsigned(1006, 12), 1766 => to_unsigned(2614, 12), 1767 => to_unsigned(3013, 12), 1768 => to_unsigned(1615, 12), 1769 => to_unsigned(2047, 12), 1770 => to_unsigned(3975, 12), 1771 => to_unsigned(3961, 12), 1772 => to_unsigned(2273, 12), 1773 => to_unsigned(3034, 12), 1774 => to_unsigned(918, 12), 1775 => to_unsigned(1698, 12), 1776 => to_unsigned(2268, 12), 1777 => to_unsigned(2308, 12), 1778 => to_unsigned(2025, 12), 1779 => to_unsigned(3047, 12), 1780 => to_unsigned(3511, 12), 1781 => to_unsigned(3145, 12), 1782 => to_unsigned(3152, 12), 1783 => to_unsigned(3004, 12), 1784 => to_unsigned(282, 12), 1785 => to_unsigned(3877, 12), 1786 => to_unsigned(1918, 12), 1787 => to_unsigned(1069, 12), 1788 => to_unsigned(3962, 12), 1789 => to_unsigned(486, 12), 1790 => to_unsigned(2372, 12), 1791 => to_unsigned(1419, 12), 1792 => to_unsigned(1725, 12), 1793 => to_unsigned(402, 12), 1794 => to_unsigned(2016, 12), 1795 => to_unsigned(2263, 12), 1796 => to_unsigned(1424, 12), 1797 => to_unsigned(2175, 12), 1798 => to_unsigned(1165, 12), 1799 => to_unsigned(3331, 12), 1800 => to_unsigned(1264, 12), 1801 => to_unsigned(2444, 12), 1802 => to_unsigned(3195, 12), 1803 => to_unsigned(4017, 12), 1804 => to_unsigned(1863, 12), 1805 => to_unsigned(1884, 12), 1806 => to_unsigned(2330, 12), 1807 => to_unsigned(1644, 12), 1808 => to_unsigned(2139, 12), 1809 => to_unsigned(2440, 12), 1810 => to_unsigned(3941, 12), 1811 => to_unsigned(157, 12), 1812 => to_unsigned(613, 12), 1813 => to_unsigned(1253, 12), 1814 => to_unsigned(2489, 12), 1815 => to_unsigned(2747, 12), 1816 => to_unsigned(1072, 12), 1817 => to_unsigned(3215, 12), 1818 => to_unsigned(1017, 12), 1819 => to_unsigned(3809, 12), 1820 => to_unsigned(3590, 12), 1821 => to_unsigned(3271, 12), 1822 => to_unsigned(1479, 12), 1823 => to_unsigned(1188, 12), 1824 => to_unsigned(2196, 12), 1825 => to_unsigned(424, 12), 1826 => to_unsigned(1200, 12), 1827 => to_unsigned(235, 12), 1828 => to_unsigned(2132, 12), 1829 => to_unsigned(417, 12), 1830 => to_unsigned(2723, 12), 1831 => to_unsigned(214, 12), 1832 => to_unsigned(2618, 12), 1833 => to_unsigned(1933, 12), 1834 => to_unsigned(4014, 12), 1835 => to_unsigned(3523, 12), 1836 => to_unsigned(370, 12), 1837 => to_unsigned(2890, 12), 1838 => to_unsigned(32, 12), 1839 => to_unsigned(896, 12), 1840 => to_unsigned(1288, 12), 1841 => to_unsigned(2110, 12), 1842 => to_unsigned(2467, 12), 1843 => to_unsigned(2754, 12), 1844 => to_unsigned(3082, 12), 1845 => to_unsigned(176, 12), 1846 => to_unsigned(1311, 12), 1847 => to_unsigned(2989, 12), 1848 => to_unsigned(4051, 12), 1849 => to_unsigned(1470, 12), 1850 => to_unsigned(1525, 12), 1851 => to_unsigned(1363, 12), 1852 => to_unsigned(1891, 12), 1853 => to_unsigned(646, 12), 1854 => to_unsigned(3512, 12), 1855 => to_unsigned(1491, 12), 1856 => to_unsigned(1339, 12), 1857 => to_unsigned(1254, 12), 1858 => to_unsigned(1526, 12), 1859 => to_unsigned(1980, 12), 1860 => to_unsigned(849, 12), 1861 => to_unsigned(1342, 12), 1862 => to_unsigned(2330, 12), 1863 => to_unsigned(250, 12), 1864 => to_unsigned(2818, 12), 1865 => to_unsigned(1899, 12), 1866 => to_unsigned(3416, 12), 1867 => to_unsigned(2521, 12), 1868 => to_unsigned(1832, 12), 1869 => to_unsigned(499, 12), 1870 => to_unsigned(2161, 12), 1871 => to_unsigned(3412, 12), 1872 => to_unsigned(4042, 12), 1873 => to_unsigned(1715, 12), 1874 => to_unsigned(2962, 12), 1875 => to_unsigned(3261, 12), 1876 => to_unsigned(1765, 12), 1877 => to_unsigned(839, 12), 1878 => to_unsigned(2284, 12), 1879 => to_unsigned(2564, 12), 1880 => to_unsigned(2209, 12), 1881 => to_unsigned(903, 12), 1882 => to_unsigned(553, 12), 1883 => to_unsigned(2818, 12), 1884 => to_unsigned(446, 12), 1885 => to_unsigned(2986, 12), 1886 => to_unsigned(760, 12), 1887 => to_unsigned(2972, 12), 1888 => to_unsigned(537, 12), 1889 => to_unsigned(56, 12), 1890 => to_unsigned(1049, 12), 1891 => to_unsigned(982, 12), 1892 => to_unsigned(3505, 12), 1893 => to_unsigned(181, 12), 1894 => to_unsigned(221, 12), 1895 => to_unsigned(4030, 12), 1896 => to_unsigned(218, 12), 1897 => to_unsigned(3006, 12), 1898 => to_unsigned(3901, 12), 1899 => to_unsigned(371, 12), 1900 => to_unsigned(1853, 12), 1901 => to_unsigned(1662, 12), 1902 => to_unsigned(1144, 12), 1903 => to_unsigned(3672, 12), 1904 => to_unsigned(123, 12), 1905 => to_unsigned(3347, 12), 1906 => to_unsigned(3808, 12), 1907 => to_unsigned(809, 12), 1908 => to_unsigned(880, 12), 1909 => to_unsigned(3056, 12), 1910 => to_unsigned(2583, 12), 1911 => to_unsigned(53, 12), 1912 => to_unsigned(524, 12), 1913 => to_unsigned(3808, 12), 1914 => to_unsigned(78, 12), 1915 => to_unsigned(1961, 12), 1916 => to_unsigned(305, 12), 1917 => to_unsigned(2588, 12), 1918 => to_unsigned(3000, 12), 1919 => to_unsigned(3623, 12), 1920 => to_unsigned(1497, 12), 1921 => to_unsigned(2121, 12), 1922 => to_unsigned(2508, 12), 1923 => to_unsigned(1777, 12), 1924 => to_unsigned(2317, 12), 1925 => to_unsigned(1016, 12), 1926 => to_unsigned(805, 12), 1927 => to_unsigned(1499, 12), 1928 => to_unsigned(3912, 12), 1929 => to_unsigned(2601, 12), 1930 => to_unsigned(1598, 12), 1931 => to_unsigned(2856, 12), 1932 => to_unsigned(1569, 12), 1933 => to_unsigned(765, 12), 1934 => to_unsigned(1024, 12), 1935 => to_unsigned(2063, 12), 1936 => to_unsigned(3366, 12), 1937 => to_unsigned(419, 12), 1938 => to_unsigned(275, 12), 1939 => to_unsigned(1508, 12), 1940 => to_unsigned(3878, 12), 1941 => to_unsigned(3937, 12), 1942 => to_unsigned(1127, 12), 1943 => to_unsigned(1485, 12), 1944 => to_unsigned(548, 12), 1945 => to_unsigned(619, 12), 1946 => to_unsigned(3392, 12), 1947 => to_unsigned(1192, 12), 1948 => to_unsigned(2442, 12), 1949 => to_unsigned(2343, 12), 1950 => to_unsigned(1256, 12), 1951 => to_unsigned(2322, 12), 1952 => to_unsigned(3438, 12), 1953 => to_unsigned(4012, 12), 1954 => to_unsigned(3494, 12), 1955 => to_unsigned(3, 12), 1956 => to_unsigned(2787, 12), 1957 => to_unsigned(4069, 12), 1958 => to_unsigned(253, 12), 1959 => to_unsigned(2802, 12), 1960 => to_unsigned(767, 12), 1961 => to_unsigned(3406, 12), 1962 => to_unsigned(3026, 12), 1963 => to_unsigned(593, 12), 1964 => to_unsigned(2293, 12), 1965 => to_unsigned(133, 12), 1966 => to_unsigned(1097, 12), 1967 => to_unsigned(2867, 12), 1968 => to_unsigned(3663, 12), 1969 => to_unsigned(3530, 12), 1970 => to_unsigned(1958, 12), 1971 => to_unsigned(884, 12), 1972 => to_unsigned(2206, 12), 1973 => to_unsigned(3717, 12), 1974 => to_unsigned(3275, 12), 1975 => to_unsigned(2326, 12), 1976 => to_unsigned(1513, 12), 1977 => to_unsigned(1916, 12), 1978 => to_unsigned(3671, 12), 1979 => to_unsigned(1945, 12), 1980 => to_unsigned(2837, 12), 1981 => to_unsigned(2119, 12), 1982 => to_unsigned(1969, 12), 1983 => to_unsigned(2577, 12), 1984 => to_unsigned(862, 12), 1985 => to_unsigned(1738, 12), 1986 => to_unsigned(1921, 12), 1987 => to_unsigned(2377, 12), 1988 => to_unsigned(1391, 12), 1989 => to_unsigned(3720, 12), 1990 => to_unsigned(3973, 12), 1991 => to_unsigned(3018, 12), 1992 => to_unsigned(996, 12), 1993 => to_unsigned(3677, 12), 1994 => to_unsigned(1454, 12), 1995 => to_unsigned(3512, 12), 1996 => to_unsigned(699, 12), 1997 => to_unsigned(2417, 12), 1998 => to_unsigned(3360, 12), 1999 => to_unsigned(3297, 12), 2000 => to_unsigned(1535, 12), 2001 => to_unsigned(3725, 12), 2002 => to_unsigned(2325, 12), 2003 => to_unsigned(1914, 12), 2004 => to_unsigned(3610, 12), 2005 => to_unsigned(3708, 12), 2006 => to_unsigned(3976, 12), 2007 => to_unsigned(1949, 12), 2008 => to_unsigned(2796, 12), 2009 => to_unsigned(2746, 12), 2010 => to_unsigned(962, 12), 2011 => to_unsigned(2327, 12), 2012 => to_unsigned(3330, 12), 2013 => to_unsigned(725, 12), 2014 => to_unsigned(1851, 12), 2015 => to_unsigned(1755, 12), 2016 => to_unsigned(3609, 12), 2017 => to_unsigned(3264, 12), 2018 => to_unsigned(2451, 12), 2019 => to_unsigned(1155, 12), 2020 => to_unsigned(628, 12), 2021 => to_unsigned(4013, 12), 2022 => to_unsigned(483, 12), 2023 => to_unsigned(3063, 12), 2024 => to_unsigned(962, 12), 2025 => to_unsigned(1731, 12), 2026 => to_unsigned(2277, 12), 2027 => to_unsigned(1473, 12), 2028 => to_unsigned(3315, 12), 2029 => to_unsigned(1609, 12), 2030 => to_unsigned(96, 12), 2031 => to_unsigned(3302, 12), 2032 => to_unsigned(3253, 12), 2033 => to_unsigned(602, 12), 2034 => to_unsigned(2668, 12), 2035 => to_unsigned(2563, 12), 2036 => to_unsigned(1639, 12), 2037 => to_unsigned(3391, 12), 2038 => to_unsigned(2591, 12), 2039 => to_unsigned(166, 12), 2040 => to_unsigned(2172, 12), 2041 => to_unsigned(3582, 12), 2042 => to_unsigned(3172, 12), 2043 => to_unsigned(284, 12), 2044 => to_unsigned(772, 12), 2045 => to_unsigned(2226, 12), 2046 => to_unsigned(1343, 12), 2047 => to_unsigned(2441, 12)),
            1 => (0 => to_unsigned(1192, 12), 1 => to_unsigned(3856, 12), 2 => to_unsigned(4046, 12), 3 => to_unsigned(2792, 12), 4 => to_unsigned(1498, 12), 5 => to_unsigned(1759, 12), 6 => to_unsigned(1875, 12), 7 => to_unsigned(1454, 12), 8 => to_unsigned(1620, 12), 9 => to_unsigned(3019, 12), 10 => to_unsigned(3761, 12), 11 => to_unsigned(1930, 12), 12 => to_unsigned(1904, 12), 13 => to_unsigned(405, 12), 14 => to_unsigned(711, 12), 15 => to_unsigned(501, 12), 16 => to_unsigned(1964, 12), 17 => to_unsigned(886, 12), 18 => to_unsigned(3840, 12), 19 => to_unsigned(882, 12), 20 => to_unsigned(1486, 12), 21 => to_unsigned(1069, 12), 22 => to_unsigned(3275, 12), 23 => to_unsigned(560, 12), 24 => to_unsigned(3656, 12), 25 => to_unsigned(3895, 12), 26 => to_unsigned(2287, 12), 27 => to_unsigned(4087, 12), 28 => to_unsigned(3484, 12), 29 => to_unsigned(974, 12), 30 => to_unsigned(742, 12), 31 => to_unsigned(2647, 12), 32 => to_unsigned(3379, 12), 33 => to_unsigned(3778, 12), 34 => to_unsigned(3055, 12), 35 => to_unsigned(438, 12), 36 => to_unsigned(1957, 12), 37 => to_unsigned(699, 12), 38 => to_unsigned(3899, 12), 39 => to_unsigned(1767, 12), 40 => to_unsigned(614, 12), 41 => to_unsigned(2232, 12), 42 => to_unsigned(3387, 12), 43 => to_unsigned(396, 12), 44 => to_unsigned(816, 12), 45 => to_unsigned(3879, 12), 46 => to_unsigned(2822, 12), 47 => to_unsigned(1804, 12), 48 => to_unsigned(422, 12), 49 => to_unsigned(3596, 12), 50 => to_unsigned(2179, 12), 51 => to_unsigned(1360, 12), 52 => to_unsigned(728, 12), 53 => to_unsigned(3360, 12), 54 => to_unsigned(3368, 12), 55 => to_unsigned(643, 12), 56 => to_unsigned(143, 12), 57 => to_unsigned(2788, 12), 58 => to_unsigned(3983, 12), 59 => to_unsigned(1223, 12), 60 => to_unsigned(1351, 12), 61 => to_unsigned(1337, 12), 62 => to_unsigned(247, 12), 63 => to_unsigned(282, 12), 64 => to_unsigned(3334, 12), 65 => to_unsigned(3626, 12), 66 => to_unsigned(372, 12), 67 => to_unsigned(510, 12), 68 => to_unsigned(2906, 12), 69 => to_unsigned(4015, 12), 70 => to_unsigned(2098, 12), 71 => to_unsigned(3860, 12), 72 => to_unsigned(702, 12), 73 => to_unsigned(2652, 12), 74 => to_unsigned(1234, 12), 75 => to_unsigned(1407, 12), 76 => to_unsigned(2847, 12), 77 => to_unsigned(3212, 12), 78 => to_unsigned(220, 12), 79 => to_unsigned(2758, 12), 80 => to_unsigned(158, 12), 81 => to_unsigned(1256, 12), 82 => to_unsigned(373, 12), 83 => to_unsigned(820, 12), 84 => to_unsigned(585, 12), 85 => to_unsigned(1962, 12), 86 => to_unsigned(2573, 12), 87 => to_unsigned(2414, 12), 88 => to_unsigned(2145, 12), 89 => to_unsigned(241, 12), 90 => to_unsigned(642, 12), 91 => to_unsigned(1214, 12), 92 => to_unsigned(684, 12), 93 => to_unsigned(112, 12), 94 => to_unsigned(1556, 12), 95 => to_unsigned(1242, 12), 96 => to_unsigned(2973, 12), 97 => to_unsigned(2403, 12), 98 => to_unsigned(2775, 12), 99 => to_unsigned(2765, 12), 100 => to_unsigned(3517, 12), 101 => to_unsigned(3711, 12), 102 => to_unsigned(2239, 12), 103 => to_unsigned(2115, 12), 104 => to_unsigned(3034, 12), 105 => to_unsigned(870, 12), 106 => to_unsigned(3875, 12), 107 => to_unsigned(2783, 12), 108 => to_unsigned(2027, 12), 109 => to_unsigned(2909, 12), 110 => to_unsigned(1495, 12), 111 => to_unsigned(3035, 12), 112 => to_unsigned(1999, 12), 113 => to_unsigned(398, 12), 114 => to_unsigned(1275, 12), 115 => to_unsigned(1667, 12), 116 => to_unsigned(716, 12), 117 => to_unsigned(565, 12), 118 => to_unsigned(2772, 12), 119 => to_unsigned(2601, 12), 120 => to_unsigned(2347, 12), 121 => to_unsigned(1791, 12), 122 => to_unsigned(756, 12), 123 => to_unsigned(78, 12), 124 => to_unsigned(3340, 12), 125 => to_unsigned(3026, 12), 126 => to_unsigned(4083, 12), 127 => to_unsigned(1098, 12), 128 => to_unsigned(1846, 12), 129 => to_unsigned(3975, 12), 130 => to_unsigned(718, 12), 131 => to_unsigned(1863, 12), 132 => to_unsigned(1366, 12), 133 => to_unsigned(859, 12), 134 => to_unsigned(107, 12), 135 => to_unsigned(3846, 12), 136 => to_unsigned(1515, 12), 137 => to_unsigned(241, 12), 138 => to_unsigned(470, 12), 139 => to_unsigned(1134, 12), 140 => to_unsigned(3353, 12), 141 => to_unsigned(3701, 12), 142 => to_unsigned(2160, 12), 143 => to_unsigned(2938, 12), 144 => to_unsigned(566, 12), 145 => to_unsigned(1738, 12), 146 => to_unsigned(629, 12), 147 => to_unsigned(610, 12), 148 => to_unsigned(1485, 12), 149 => to_unsigned(3263, 12), 150 => to_unsigned(3054, 12), 151 => to_unsigned(1229, 12), 152 => to_unsigned(2973, 12), 153 => to_unsigned(2055, 12), 154 => to_unsigned(2730, 12), 155 => to_unsigned(2496, 12), 156 => to_unsigned(886, 12), 157 => to_unsigned(1724, 12), 158 => to_unsigned(616, 12), 159 => to_unsigned(2866, 12), 160 => to_unsigned(4095, 12), 161 => to_unsigned(3806, 12), 162 => to_unsigned(187, 12), 163 => to_unsigned(301, 12), 164 => to_unsigned(2933, 12), 165 => to_unsigned(4086, 12), 166 => to_unsigned(1906, 12), 167 => to_unsigned(2356, 12), 168 => to_unsigned(1500, 12), 169 => to_unsigned(275, 12), 170 => to_unsigned(1513, 12), 171 => to_unsigned(2642, 12), 172 => to_unsigned(807, 12), 173 => to_unsigned(1171, 12), 174 => to_unsigned(2052, 12), 175 => to_unsigned(1016, 12), 176 => to_unsigned(2335, 12), 177 => to_unsigned(3732, 12), 178 => to_unsigned(1896, 12), 179 => to_unsigned(2218, 12), 180 => to_unsigned(2120, 12), 181 => to_unsigned(1290, 12), 182 => to_unsigned(1194, 12), 183 => to_unsigned(812, 12), 184 => to_unsigned(632, 12), 185 => to_unsigned(1919, 12), 186 => to_unsigned(149, 12), 187 => to_unsigned(3319, 12), 188 => to_unsigned(392, 12), 189 => to_unsigned(567, 12), 190 => to_unsigned(1059, 12), 191 => to_unsigned(367, 12), 192 => to_unsigned(351, 12), 193 => to_unsigned(3523, 12), 194 => to_unsigned(2057, 12), 195 => to_unsigned(1581, 12), 196 => to_unsigned(46, 12), 197 => to_unsigned(3836, 12), 198 => to_unsigned(1840, 12), 199 => to_unsigned(2325, 12), 200 => to_unsigned(986, 12), 201 => to_unsigned(585, 12), 202 => to_unsigned(2599, 12), 203 => to_unsigned(1967, 12), 204 => to_unsigned(3956, 12), 205 => to_unsigned(2949, 12), 206 => to_unsigned(590, 12), 207 => to_unsigned(1296, 12), 208 => to_unsigned(147, 12), 209 => to_unsigned(49, 12), 210 => to_unsigned(1346, 12), 211 => to_unsigned(16, 12), 212 => to_unsigned(2613, 12), 213 => to_unsigned(1014, 12), 214 => to_unsigned(4074, 12), 215 => to_unsigned(3434, 12), 216 => to_unsigned(1410, 12), 217 => to_unsigned(1929, 12), 218 => to_unsigned(1831, 12), 219 => to_unsigned(3655, 12), 220 => to_unsigned(1328, 12), 221 => to_unsigned(1760, 12), 222 => to_unsigned(3415, 12), 223 => to_unsigned(2736, 12), 224 => to_unsigned(3879, 12), 225 => to_unsigned(2928, 12), 226 => to_unsigned(3579, 12), 227 => to_unsigned(1147, 12), 228 => to_unsigned(1961, 12), 229 => to_unsigned(1548, 12), 230 => to_unsigned(1612, 12), 231 => to_unsigned(3823, 12), 232 => to_unsigned(3683, 12), 233 => to_unsigned(3532, 12), 234 => to_unsigned(3688, 12), 235 => to_unsigned(383, 12), 236 => to_unsigned(2941, 12), 237 => to_unsigned(584, 12), 238 => to_unsigned(1825, 12), 239 => to_unsigned(2845, 12), 240 => to_unsigned(2096, 12), 241 => to_unsigned(1312, 12), 242 => to_unsigned(1145, 12), 243 => to_unsigned(2250, 12), 244 => to_unsigned(2800, 12), 245 => to_unsigned(3416, 12), 246 => to_unsigned(1717, 12), 247 => to_unsigned(477, 12), 248 => to_unsigned(3264, 12), 249 => to_unsigned(196, 12), 250 => to_unsigned(599, 12), 251 => to_unsigned(1040, 12), 252 => to_unsigned(3280, 12), 253 => to_unsigned(2245, 12), 254 => to_unsigned(1452, 12), 255 => to_unsigned(1218, 12), 256 => to_unsigned(3689, 12), 257 => to_unsigned(1848, 12), 258 => to_unsigned(3855, 12), 259 => to_unsigned(3763, 12), 260 => to_unsigned(1908, 12), 261 => to_unsigned(2523, 12), 262 => to_unsigned(3716, 12), 263 => to_unsigned(1913, 12), 264 => to_unsigned(3940, 12), 265 => to_unsigned(1326, 12), 266 => to_unsigned(3805, 12), 267 => to_unsigned(3410, 12), 268 => to_unsigned(1443, 12), 269 => to_unsigned(2141, 12), 270 => to_unsigned(375, 12), 271 => to_unsigned(869, 12), 272 => to_unsigned(2521, 12), 273 => to_unsigned(3088, 12), 274 => to_unsigned(1511, 12), 275 => to_unsigned(2762, 12), 276 => to_unsigned(1559, 12), 277 => to_unsigned(451, 12), 278 => to_unsigned(644, 12), 279 => to_unsigned(1581, 12), 280 => to_unsigned(3207, 12), 281 => to_unsigned(311, 12), 282 => to_unsigned(1242, 12), 283 => to_unsigned(3968, 12), 284 => to_unsigned(2771, 12), 285 => to_unsigned(1180, 12), 286 => to_unsigned(95, 12), 287 => to_unsigned(2802, 12), 288 => to_unsigned(1978, 12), 289 => to_unsigned(2118, 12), 290 => to_unsigned(871, 12), 291 => to_unsigned(3557, 12), 292 => to_unsigned(3072, 12), 293 => to_unsigned(95, 12), 294 => to_unsigned(3221, 12), 295 => to_unsigned(2736, 12), 296 => to_unsigned(3279, 12), 297 => to_unsigned(2623, 12), 298 => to_unsigned(2155, 12), 299 => to_unsigned(3342, 12), 300 => to_unsigned(2197, 12), 301 => to_unsigned(2556, 12), 302 => to_unsigned(1597, 12), 303 => to_unsigned(3182, 12), 304 => to_unsigned(3671, 12), 305 => to_unsigned(855, 12), 306 => to_unsigned(1393, 12), 307 => to_unsigned(447, 12), 308 => to_unsigned(1675, 12), 309 => to_unsigned(2087, 12), 310 => to_unsigned(3204, 12), 311 => to_unsigned(4000, 12), 312 => to_unsigned(3948, 12), 313 => to_unsigned(3259, 12), 314 => to_unsigned(114, 12), 315 => to_unsigned(3566, 12), 316 => to_unsigned(2497, 12), 317 => to_unsigned(3647, 12), 318 => to_unsigned(3993, 12), 319 => to_unsigned(2858, 12), 320 => to_unsigned(83, 12), 321 => to_unsigned(847, 12), 322 => to_unsigned(393, 12), 323 => to_unsigned(2280, 12), 324 => to_unsigned(2126, 12), 325 => to_unsigned(2506, 12), 326 => to_unsigned(1300, 12), 327 => to_unsigned(457, 12), 328 => to_unsigned(645, 12), 329 => to_unsigned(467, 12), 330 => to_unsigned(520, 12), 331 => to_unsigned(527, 12), 332 => to_unsigned(2746, 12), 333 => to_unsigned(2127, 12), 334 => to_unsigned(980, 12), 335 => to_unsigned(2186, 12), 336 => to_unsigned(294, 12), 337 => to_unsigned(106, 12), 338 => to_unsigned(4095, 12), 339 => to_unsigned(1610, 12), 340 => to_unsigned(2239, 12), 341 => to_unsigned(2407, 12), 342 => to_unsigned(2187, 12), 343 => to_unsigned(2165, 12), 344 => to_unsigned(2979, 12), 345 => to_unsigned(1826, 12), 346 => to_unsigned(753, 12), 347 => to_unsigned(2255, 12), 348 => to_unsigned(683, 12), 349 => to_unsigned(1889, 12), 350 => to_unsigned(1289, 12), 351 => to_unsigned(1874, 12), 352 => to_unsigned(1375, 12), 353 => to_unsigned(2814, 12), 354 => to_unsigned(3617, 12), 355 => to_unsigned(2097, 12), 356 => to_unsigned(3570, 12), 357 => to_unsigned(158, 12), 358 => to_unsigned(1478, 12), 359 => to_unsigned(3647, 12), 360 => to_unsigned(3341, 12), 361 => to_unsigned(1534, 12), 362 => to_unsigned(2696, 12), 363 => to_unsigned(1479, 12), 364 => to_unsigned(1826, 12), 365 => to_unsigned(1304, 12), 366 => to_unsigned(3075, 12), 367 => to_unsigned(1685, 12), 368 => to_unsigned(941, 12), 369 => to_unsigned(2179, 12), 370 => to_unsigned(2296, 12), 371 => to_unsigned(1753, 12), 372 => to_unsigned(171, 12), 373 => to_unsigned(3639, 12), 374 => to_unsigned(3299, 12), 375 => to_unsigned(423, 12), 376 => to_unsigned(3430, 12), 377 => to_unsigned(193, 12), 378 => to_unsigned(1810, 12), 379 => to_unsigned(3174, 12), 380 => to_unsigned(3287, 12), 381 => to_unsigned(3569, 12), 382 => to_unsigned(608, 12), 383 => to_unsigned(395, 12), 384 => to_unsigned(1697, 12), 385 => to_unsigned(1008, 12), 386 => to_unsigned(477, 12), 387 => to_unsigned(3931, 12), 388 => to_unsigned(3444, 12), 389 => to_unsigned(3491, 12), 390 => to_unsigned(979, 12), 391 => to_unsigned(1635, 12), 392 => to_unsigned(2893, 12), 393 => to_unsigned(2206, 12), 394 => to_unsigned(1207, 12), 395 => to_unsigned(1739, 12), 396 => to_unsigned(2317, 12), 397 => to_unsigned(3444, 12), 398 => to_unsigned(597, 12), 399 => to_unsigned(1833, 12), 400 => to_unsigned(2563, 12), 401 => to_unsigned(3870, 12), 402 => to_unsigned(2458, 12), 403 => to_unsigned(434, 12), 404 => to_unsigned(675, 12), 405 => to_unsigned(3635, 12), 406 => to_unsigned(1734, 12), 407 => to_unsigned(1345, 12), 408 => to_unsigned(892, 12), 409 => to_unsigned(3872, 12), 410 => to_unsigned(2642, 12), 411 => to_unsigned(764, 12), 412 => to_unsigned(3233, 12), 413 => to_unsigned(3409, 12), 414 => to_unsigned(897, 12), 415 => to_unsigned(3657, 12), 416 => to_unsigned(311, 12), 417 => to_unsigned(4077, 12), 418 => to_unsigned(3908, 12), 419 => to_unsigned(423, 12), 420 => to_unsigned(2145, 12), 421 => to_unsigned(3208, 12), 422 => to_unsigned(1670, 12), 423 => to_unsigned(3440, 12), 424 => to_unsigned(1928, 12), 425 => to_unsigned(1321, 12), 426 => to_unsigned(1641, 12), 427 => to_unsigned(941, 12), 428 => to_unsigned(3671, 12), 429 => to_unsigned(320, 12), 430 => to_unsigned(2055, 12), 431 => to_unsigned(2448, 12), 432 => to_unsigned(3725, 12), 433 => to_unsigned(1613, 12), 434 => to_unsigned(3500, 12), 435 => to_unsigned(2914, 12), 436 => to_unsigned(2197, 12), 437 => to_unsigned(431, 12), 438 => to_unsigned(1312, 12), 439 => to_unsigned(1253, 12), 440 => to_unsigned(475, 12), 441 => to_unsigned(1912, 12), 442 => to_unsigned(2889, 12), 443 => to_unsigned(3353, 12), 444 => to_unsigned(1915, 12), 445 => to_unsigned(206, 12), 446 => to_unsigned(1203, 12), 447 => to_unsigned(3070, 12), 448 => to_unsigned(1219, 12), 449 => to_unsigned(333, 12), 450 => to_unsigned(3700, 12), 451 => to_unsigned(1938, 12), 452 => to_unsigned(1164, 12), 453 => to_unsigned(3561, 12), 454 => to_unsigned(3105, 12), 455 => to_unsigned(551, 12), 456 => to_unsigned(1727, 12), 457 => to_unsigned(1594, 12), 458 => to_unsigned(1297, 12), 459 => to_unsigned(629, 12), 460 => to_unsigned(2973, 12), 461 => to_unsigned(3834, 12), 462 => to_unsigned(1089, 12), 463 => to_unsigned(968, 12), 464 => to_unsigned(3678, 12), 465 => to_unsigned(425, 12), 466 => to_unsigned(2133, 12), 467 => to_unsigned(1313, 12), 468 => to_unsigned(2905, 12), 469 => to_unsigned(358, 12), 470 => to_unsigned(822, 12), 471 => to_unsigned(3698, 12), 472 => to_unsigned(3993, 12), 473 => to_unsigned(3712, 12), 474 => to_unsigned(1540, 12), 475 => to_unsigned(3633, 12), 476 => to_unsigned(51, 12), 477 => to_unsigned(3815, 12), 478 => to_unsigned(3018, 12), 479 => to_unsigned(1689, 12), 480 => to_unsigned(4001, 12), 481 => to_unsigned(2308, 12), 482 => to_unsigned(2714, 12), 483 => to_unsigned(2354, 12), 484 => to_unsigned(3503, 12), 485 => to_unsigned(2397, 12), 486 => to_unsigned(2730, 12), 487 => to_unsigned(3532, 12), 488 => to_unsigned(1464, 12), 489 => to_unsigned(3587, 12), 490 => to_unsigned(1191, 12), 491 => to_unsigned(3998, 12), 492 => to_unsigned(3158, 12), 493 => to_unsigned(266, 12), 494 => to_unsigned(929, 12), 495 => to_unsigned(2320, 12), 496 => to_unsigned(1345, 12), 497 => to_unsigned(3366, 12), 498 => to_unsigned(365, 12), 499 => to_unsigned(2831, 12), 500 => to_unsigned(125, 12), 501 => to_unsigned(1570, 12), 502 => to_unsigned(3288, 12), 503 => to_unsigned(4048, 12), 504 => to_unsigned(1736, 12), 505 => to_unsigned(3010, 12), 506 => to_unsigned(2602, 12), 507 => to_unsigned(2382, 12), 508 => to_unsigned(3818, 12), 509 => to_unsigned(519, 12), 510 => to_unsigned(1208, 12), 511 => to_unsigned(938, 12), 512 => to_unsigned(1277, 12), 513 => to_unsigned(1877, 12), 514 => to_unsigned(2757, 12), 515 => to_unsigned(2561, 12), 516 => to_unsigned(741, 12), 517 => to_unsigned(3146, 12), 518 => to_unsigned(544, 12), 519 => to_unsigned(584, 12), 520 => to_unsigned(3334, 12), 521 => to_unsigned(873, 12), 522 => to_unsigned(9, 12), 523 => to_unsigned(1074, 12), 524 => to_unsigned(1327, 12), 525 => to_unsigned(2205, 12), 526 => to_unsigned(2252, 12), 527 => to_unsigned(2834, 12), 528 => to_unsigned(2203, 12), 529 => to_unsigned(4078, 12), 530 => to_unsigned(3988, 12), 531 => to_unsigned(580, 12), 532 => to_unsigned(2796, 12), 533 => to_unsigned(3326, 12), 534 => to_unsigned(1419, 12), 535 => to_unsigned(80, 12), 536 => to_unsigned(2409, 12), 537 => to_unsigned(3111, 12), 538 => to_unsigned(3716, 12), 539 => to_unsigned(3121, 12), 540 => to_unsigned(2735, 12), 541 => to_unsigned(2918, 12), 542 => to_unsigned(463, 12), 543 => to_unsigned(3164, 12), 544 => to_unsigned(4053, 12), 545 => to_unsigned(3798, 12), 546 => to_unsigned(2951, 12), 547 => to_unsigned(2275, 12), 548 => to_unsigned(1489, 12), 549 => to_unsigned(3461, 12), 550 => to_unsigned(4092, 12), 551 => to_unsigned(3259, 12), 552 => to_unsigned(3001, 12), 553 => to_unsigned(528, 12), 554 => to_unsigned(536, 12), 555 => to_unsigned(2977, 12), 556 => to_unsigned(1746, 12), 557 => to_unsigned(1164, 12), 558 => to_unsigned(3664, 12), 559 => to_unsigned(1983, 12), 560 => to_unsigned(1801, 12), 561 => to_unsigned(2594, 12), 562 => to_unsigned(823, 12), 563 => to_unsigned(1888, 12), 564 => to_unsigned(217, 12), 565 => to_unsigned(153, 12), 566 => to_unsigned(2618, 12), 567 => to_unsigned(1183, 12), 568 => to_unsigned(1700, 12), 569 => to_unsigned(1119, 12), 570 => to_unsigned(972, 12), 571 => to_unsigned(2060, 12), 572 => to_unsigned(1362, 12), 573 => to_unsigned(1266, 12), 574 => to_unsigned(2983, 12), 575 => to_unsigned(1866, 12), 576 => to_unsigned(2630, 12), 577 => to_unsigned(2236, 12), 578 => to_unsigned(3481, 12), 579 => to_unsigned(3194, 12), 580 => to_unsigned(3847, 12), 581 => to_unsigned(1800, 12), 582 => to_unsigned(3583, 12), 583 => to_unsigned(3248, 12), 584 => to_unsigned(805, 12), 585 => to_unsigned(173, 12), 586 => to_unsigned(1409, 12), 587 => to_unsigned(506, 12), 588 => to_unsigned(122, 12), 589 => to_unsigned(1859, 12), 590 => to_unsigned(1735, 12), 591 => to_unsigned(535, 12), 592 => to_unsigned(2659, 12), 593 => to_unsigned(2647, 12), 594 => to_unsigned(2178, 12), 595 => to_unsigned(3793, 12), 596 => to_unsigned(15, 12), 597 => to_unsigned(638, 12), 598 => to_unsigned(3433, 12), 599 => to_unsigned(2190, 12), 600 => to_unsigned(2379, 12), 601 => to_unsigned(3307, 12), 602 => to_unsigned(1508, 12), 603 => to_unsigned(2833, 12), 604 => to_unsigned(1461, 12), 605 => to_unsigned(742, 12), 606 => to_unsigned(3872, 12), 607 => to_unsigned(3383, 12), 608 => to_unsigned(3645, 12), 609 => to_unsigned(1829, 12), 610 => to_unsigned(2308, 12), 611 => to_unsigned(2319, 12), 612 => to_unsigned(1862, 12), 613 => to_unsigned(326, 12), 614 => to_unsigned(1652, 12), 615 => to_unsigned(1593, 12), 616 => to_unsigned(2390, 12), 617 => to_unsigned(1809, 12), 618 => to_unsigned(3664, 12), 619 => to_unsigned(3139, 12), 620 => to_unsigned(576, 12), 621 => to_unsigned(3550, 12), 622 => to_unsigned(2463, 12), 623 => to_unsigned(1899, 12), 624 => to_unsigned(799, 12), 625 => to_unsigned(787, 12), 626 => to_unsigned(3917, 12), 627 => to_unsigned(500, 12), 628 => to_unsigned(1150, 12), 629 => to_unsigned(2221, 12), 630 => to_unsigned(350, 12), 631 => to_unsigned(3523, 12), 632 => to_unsigned(3382, 12), 633 => to_unsigned(986, 12), 634 => to_unsigned(3909, 12), 635 => to_unsigned(2102, 12), 636 => to_unsigned(3894, 12), 637 => to_unsigned(1856, 12), 638 => to_unsigned(1147, 12), 639 => to_unsigned(3148, 12), 640 => to_unsigned(2093, 12), 641 => to_unsigned(688, 12), 642 => to_unsigned(261, 12), 643 => to_unsigned(2025, 12), 644 => to_unsigned(2701, 12), 645 => to_unsigned(237, 12), 646 => to_unsigned(1375, 12), 647 => to_unsigned(2635, 12), 648 => to_unsigned(3116, 12), 649 => to_unsigned(2144, 12), 650 => to_unsigned(3023, 12), 651 => to_unsigned(1696, 12), 652 => to_unsigned(2343, 12), 653 => to_unsigned(2739, 12), 654 => to_unsigned(2355, 12), 655 => to_unsigned(3771, 12), 656 => to_unsigned(2036, 12), 657 => to_unsigned(1500, 12), 658 => to_unsigned(1650, 12), 659 => to_unsigned(1903, 12), 660 => to_unsigned(1824, 12), 661 => to_unsigned(1606, 12), 662 => to_unsigned(3594, 12), 663 => to_unsigned(1755, 12), 664 => to_unsigned(1492, 12), 665 => to_unsigned(988, 12), 666 => to_unsigned(1128, 12), 667 => to_unsigned(1130, 12), 668 => to_unsigned(204, 12), 669 => to_unsigned(3501, 12), 670 => to_unsigned(2120, 12), 671 => to_unsigned(386, 12), 672 => to_unsigned(2780, 12), 673 => to_unsigned(3117, 12), 674 => to_unsigned(3624, 12), 675 => to_unsigned(3372, 12), 676 => to_unsigned(493, 12), 677 => to_unsigned(3564, 12), 678 => to_unsigned(3217, 12), 679 => to_unsigned(2250, 12), 680 => to_unsigned(1542, 12), 681 => to_unsigned(386, 12), 682 => to_unsigned(2392, 12), 683 => to_unsigned(2334, 12), 684 => to_unsigned(3484, 12), 685 => to_unsigned(2494, 12), 686 => to_unsigned(3944, 12), 687 => to_unsigned(1243, 12), 688 => to_unsigned(470, 12), 689 => to_unsigned(1676, 12), 690 => to_unsigned(452, 12), 691 => to_unsigned(2835, 12), 692 => to_unsigned(3673, 12), 693 => to_unsigned(1458, 12), 694 => to_unsigned(1559, 12), 695 => to_unsigned(2145, 12), 696 => to_unsigned(2090, 12), 697 => to_unsigned(1643, 12), 698 => to_unsigned(3501, 12), 699 => to_unsigned(2062, 12), 700 => to_unsigned(1627, 12), 701 => to_unsigned(2900, 12), 702 => to_unsigned(1424, 12), 703 => to_unsigned(4005, 12), 704 => to_unsigned(2459, 12), 705 => to_unsigned(3799, 12), 706 => to_unsigned(3953, 12), 707 => to_unsigned(152, 12), 708 => to_unsigned(2677, 12), 709 => to_unsigned(2567, 12), 710 => to_unsigned(403, 12), 711 => to_unsigned(113, 12), 712 => to_unsigned(2655, 12), 713 => to_unsigned(3378, 12), 714 => to_unsigned(2883, 12), 715 => to_unsigned(302, 12), 716 => to_unsigned(3058, 12), 717 => to_unsigned(678, 12), 718 => to_unsigned(2234, 12), 719 => to_unsigned(1516, 12), 720 => to_unsigned(817, 12), 721 => to_unsigned(3576, 12), 722 => to_unsigned(3140, 12), 723 => to_unsigned(576, 12), 724 => to_unsigned(1378, 12), 725 => to_unsigned(1135, 12), 726 => to_unsigned(675, 12), 727 => to_unsigned(3692, 12), 728 => to_unsigned(1330, 12), 729 => to_unsigned(1871, 12), 730 => to_unsigned(458, 12), 731 => to_unsigned(600, 12), 732 => to_unsigned(576, 12), 733 => to_unsigned(3932, 12), 734 => to_unsigned(3879, 12), 735 => to_unsigned(942, 12), 736 => to_unsigned(891, 12), 737 => to_unsigned(159, 12), 738 => to_unsigned(168, 12), 739 => to_unsigned(3855, 12), 740 => to_unsigned(710, 12), 741 => to_unsigned(2099, 12), 742 => to_unsigned(448, 12), 743 => to_unsigned(3443, 12), 744 => to_unsigned(1714, 12), 745 => to_unsigned(1875, 12), 746 => to_unsigned(3495, 12), 747 => to_unsigned(235, 12), 748 => to_unsigned(1483, 12), 749 => to_unsigned(2004, 12), 750 => to_unsigned(2619, 12), 751 => to_unsigned(3410, 12), 752 => to_unsigned(1172, 12), 753 => to_unsigned(1332, 12), 754 => to_unsigned(116, 12), 755 => to_unsigned(344, 12), 756 => to_unsigned(498, 12), 757 => to_unsigned(3875, 12), 758 => to_unsigned(3849, 12), 759 => to_unsigned(2072, 12), 760 => to_unsigned(1478, 12), 761 => to_unsigned(3348, 12), 762 => to_unsigned(3870, 12), 763 => to_unsigned(671, 12), 764 => to_unsigned(3464, 12), 765 => to_unsigned(3279, 12), 766 => to_unsigned(2227, 12), 767 => to_unsigned(3898, 12), 768 => to_unsigned(2361, 12), 769 => to_unsigned(2778, 12), 770 => to_unsigned(405, 12), 771 => to_unsigned(2690, 12), 772 => to_unsigned(847, 12), 773 => to_unsigned(1408, 12), 774 => to_unsigned(2077, 12), 775 => to_unsigned(3477, 12), 776 => to_unsigned(812, 12), 777 => to_unsigned(1325, 12), 778 => to_unsigned(1988, 12), 779 => to_unsigned(1672, 12), 780 => to_unsigned(2271, 12), 781 => to_unsigned(674, 12), 782 => to_unsigned(2221, 12), 783 => to_unsigned(2100, 12), 784 => to_unsigned(595, 12), 785 => to_unsigned(1361, 12), 786 => to_unsigned(2742, 12), 787 => to_unsigned(2833, 12), 788 => to_unsigned(957, 12), 789 => to_unsigned(291, 12), 790 => to_unsigned(3864, 12), 791 => to_unsigned(929, 12), 792 => to_unsigned(1535, 12), 793 => to_unsigned(1155, 12), 794 => to_unsigned(1996, 12), 795 => to_unsigned(1240, 12), 796 => to_unsigned(804, 12), 797 => to_unsigned(3369, 12), 798 => to_unsigned(3219, 12), 799 => to_unsigned(1284, 12), 800 => to_unsigned(1512, 12), 801 => to_unsigned(695, 12), 802 => to_unsigned(2682, 12), 803 => to_unsigned(2026, 12), 804 => to_unsigned(3714, 12), 805 => to_unsigned(2502, 12), 806 => to_unsigned(1620, 12), 807 => to_unsigned(490, 12), 808 => to_unsigned(3718, 12), 809 => to_unsigned(1151, 12), 810 => to_unsigned(2712, 12), 811 => to_unsigned(2671, 12), 812 => to_unsigned(2636, 12), 813 => to_unsigned(4043, 12), 814 => to_unsigned(1489, 12), 815 => to_unsigned(1055, 12), 816 => to_unsigned(3172, 12), 817 => to_unsigned(1236, 12), 818 => to_unsigned(1672, 12), 819 => to_unsigned(646, 12), 820 => to_unsigned(3653, 12), 821 => to_unsigned(386, 12), 822 => to_unsigned(2540, 12), 823 => to_unsigned(144, 12), 824 => to_unsigned(3185, 12), 825 => to_unsigned(1036, 12), 826 => to_unsigned(1575, 12), 827 => to_unsigned(390, 12), 828 => to_unsigned(4053, 12), 829 => to_unsigned(1194, 12), 830 => to_unsigned(3159, 12), 831 => to_unsigned(1055, 12), 832 => to_unsigned(1655, 12), 833 => to_unsigned(146, 12), 834 => to_unsigned(3768, 12), 835 => to_unsigned(97, 12), 836 => to_unsigned(122, 12), 837 => to_unsigned(3232, 12), 838 => to_unsigned(3749, 12), 839 => to_unsigned(1852, 12), 840 => to_unsigned(3581, 12), 841 => to_unsigned(3943, 12), 842 => to_unsigned(1913, 12), 843 => to_unsigned(2457, 12), 844 => to_unsigned(2911, 12), 845 => to_unsigned(2277, 12), 846 => to_unsigned(601, 12), 847 => to_unsigned(3039, 12), 848 => to_unsigned(2220, 12), 849 => to_unsigned(2827, 12), 850 => to_unsigned(2294, 12), 851 => to_unsigned(3700, 12), 852 => to_unsigned(640, 12), 853 => to_unsigned(1378, 12), 854 => to_unsigned(3546, 12), 855 => to_unsigned(982, 12), 856 => to_unsigned(1293, 12), 857 => to_unsigned(1532, 12), 858 => to_unsigned(2776, 12), 859 => to_unsigned(2562, 12), 860 => to_unsigned(2946, 12), 861 => to_unsigned(1139, 12), 862 => to_unsigned(1660, 12), 863 => to_unsigned(1180, 12), 864 => to_unsigned(3629, 12), 865 => to_unsigned(2382, 12), 866 => to_unsigned(3391, 12), 867 => to_unsigned(1743, 12), 868 => to_unsigned(3227, 12), 869 => to_unsigned(66, 12), 870 => to_unsigned(2488, 12), 871 => to_unsigned(1105, 12), 872 => to_unsigned(2608, 12), 873 => to_unsigned(3208, 12), 874 => to_unsigned(2523, 12), 875 => to_unsigned(2367, 12), 876 => to_unsigned(1656, 12), 877 => to_unsigned(990, 12), 878 => to_unsigned(3845, 12), 879 => to_unsigned(1597, 12), 880 => to_unsigned(1691, 12), 881 => to_unsigned(1528, 12), 882 => to_unsigned(4094, 12), 883 => to_unsigned(2089, 12), 884 => to_unsigned(146, 12), 885 => to_unsigned(145, 12), 886 => to_unsigned(704, 12), 887 => to_unsigned(3012, 12), 888 => to_unsigned(2145, 12), 889 => to_unsigned(1126, 12), 890 => to_unsigned(361, 12), 891 => to_unsigned(1932, 12), 892 => to_unsigned(2018, 12), 893 => to_unsigned(890, 12), 894 => to_unsigned(3798, 12), 895 => to_unsigned(2202, 12), 896 => to_unsigned(3340, 12), 897 => to_unsigned(1229, 12), 898 => to_unsigned(2297, 12), 899 => to_unsigned(2400, 12), 900 => to_unsigned(3955, 12), 901 => to_unsigned(320, 12), 902 => to_unsigned(791, 12), 903 => to_unsigned(3291, 12), 904 => to_unsigned(268, 12), 905 => to_unsigned(3022, 12), 906 => to_unsigned(284, 12), 907 => to_unsigned(3124, 12), 908 => to_unsigned(2243, 12), 909 => to_unsigned(153, 12), 910 => to_unsigned(2938, 12), 911 => to_unsigned(2887, 12), 912 => to_unsigned(3392, 12), 913 => to_unsigned(2389, 12), 914 => to_unsigned(1776, 12), 915 => to_unsigned(2058, 12), 916 => to_unsigned(968, 12), 917 => to_unsigned(116, 12), 918 => to_unsigned(107, 12), 919 => to_unsigned(1939, 12), 920 => to_unsigned(138, 12), 921 => to_unsigned(3233, 12), 922 => to_unsigned(2813, 12), 923 => to_unsigned(524, 12), 924 => to_unsigned(2428, 12), 925 => to_unsigned(2588, 12), 926 => to_unsigned(2973, 12), 927 => to_unsigned(1344, 12), 928 => to_unsigned(3295, 12), 929 => to_unsigned(3508, 12), 930 => to_unsigned(2982, 12), 931 => to_unsigned(2358, 12), 932 => to_unsigned(1800, 12), 933 => to_unsigned(3819, 12), 934 => to_unsigned(2709, 12), 935 => to_unsigned(1517, 12), 936 => to_unsigned(864, 12), 937 => to_unsigned(1943, 12), 938 => to_unsigned(600, 12), 939 => to_unsigned(1405, 12), 940 => to_unsigned(2170, 12), 941 => to_unsigned(1670, 12), 942 => to_unsigned(910, 12), 943 => to_unsigned(3365, 12), 944 => to_unsigned(2511, 12), 945 => to_unsigned(1499, 12), 946 => to_unsigned(2304, 12), 947 => to_unsigned(837, 12), 948 => to_unsigned(3740, 12), 949 => to_unsigned(2895, 12), 950 => to_unsigned(421, 12), 951 => to_unsigned(2881, 12), 952 => to_unsigned(3533, 12), 953 => to_unsigned(2222, 12), 954 => to_unsigned(2129, 12), 955 => to_unsigned(2170, 12), 956 => to_unsigned(2594, 12), 957 => to_unsigned(2071, 12), 958 => to_unsigned(3899, 12), 959 => to_unsigned(3173, 12), 960 => to_unsigned(1206, 12), 961 => to_unsigned(1588, 12), 962 => to_unsigned(2963, 12), 963 => to_unsigned(1903, 12), 964 => to_unsigned(2255, 12), 965 => to_unsigned(344, 12), 966 => to_unsigned(650, 12), 967 => to_unsigned(120, 12), 968 => to_unsigned(2769, 12), 969 => to_unsigned(1870, 12), 970 => to_unsigned(1295, 12), 971 => to_unsigned(2279, 12), 972 => to_unsigned(2800, 12), 973 => to_unsigned(2992, 12), 974 => to_unsigned(1465, 12), 975 => to_unsigned(3039, 12), 976 => to_unsigned(1233, 12), 977 => to_unsigned(3510, 12), 978 => to_unsigned(1732, 12), 979 => to_unsigned(3242, 12), 980 => to_unsigned(1450, 12), 981 => to_unsigned(655, 12), 982 => to_unsigned(4012, 12), 983 => to_unsigned(1865, 12), 984 => to_unsigned(2467, 12), 985 => to_unsigned(498, 12), 986 => to_unsigned(3476, 12), 987 => to_unsigned(2423, 12), 988 => to_unsigned(2164, 12), 989 => to_unsigned(796, 12), 990 => to_unsigned(2821, 12), 991 => to_unsigned(2824, 12), 992 => to_unsigned(2312, 12), 993 => to_unsigned(214, 12), 994 => to_unsigned(1338, 12), 995 => to_unsigned(1915, 12), 996 => to_unsigned(1239, 12), 997 => to_unsigned(2725, 12), 998 => to_unsigned(956, 12), 999 => to_unsigned(1656, 12), 1000 => to_unsigned(3889, 12), 1001 => to_unsigned(3968, 12), 1002 => to_unsigned(3289, 12), 1003 => to_unsigned(1547, 12), 1004 => to_unsigned(3238, 12), 1005 => to_unsigned(2291, 12), 1006 => to_unsigned(1726, 12), 1007 => to_unsigned(1860, 12), 1008 => to_unsigned(3749, 12), 1009 => to_unsigned(1516, 12), 1010 => to_unsigned(2151, 12), 1011 => to_unsigned(531, 12), 1012 => to_unsigned(1266, 12), 1013 => to_unsigned(389, 12), 1014 => to_unsigned(2229, 12), 1015 => to_unsigned(1032, 12), 1016 => to_unsigned(1565, 12), 1017 => to_unsigned(1338, 12), 1018 => to_unsigned(3573, 12), 1019 => to_unsigned(2033, 12), 1020 => to_unsigned(985, 12), 1021 => to_unsigned(191, 12), 1022 => to_unsigned(928, 12), 1023 => to_unsigned(1310, 12), 1024 => to_unsigned(2376, 12), 1025 => to_unsigned(2816, 12), 1026 => to_unsigned(1206, 12), 1027 => to_unsigned(1940, 12), 1028 => to_unsigned(2542, 12), 1029 => to_unsigned(4082, 12), 1030 => to_unsigned(2586, 12), 1031 => to_unsigned(2436, 12), 1032 => to_unsigned(2888, 12), 1033 => to_unsigned(3124, 12), 1034 => to_unsigned(3339, 12), 1035 => to_unsigned(1395, 12), 1036 => to_unsigned(228, 12), 1037 => to_unsigned(2910, 12), 1038 => to_unsigned(2408, 12), 1039 => to_unsigned(3497, 12), 1040 => to_unsigned(2525, 12), 1041 => to_unsigned(487, 12), 1042 => to_unsigned(1754, 12), 1043 => to_unsigned(848, 12), 1044 => to_unsigned(629, 12), 1045 => to_unsigned(404, 12), 1046 => to_unsigned(2639, 12), 1047 => to_unsigned(2379, 12), 1048 => to_unsigned(1756, 12), 1049 => to_unsigned(2995, 12), 1050 => to_unsigned(1995, 12), 1051 => to_unsigned(2700, 12), 1052 => to_unsigned(55, 12), 1053 => to_unsigned(2148, 12), 1054 => to_unsigned(830, 12), 1055 => to_unsigned(1376, 12), 1056 => to_unsigned(3851, 12), 1057 => to_unsigned(883, 12), 1058 => to_unsigned(3906, 12), 1059 => to_unsigned(1895, 12), 1060 => to_unsigned(201, 12), 1061 => to_unsigned(2033, 12), 1062 => to_unsigned(300, 12), 1063 => to_unsigned(2058, 12), 1064 => to_unsigned(1749, 12), 1065 => to_unsigned(885, 12), 1066 => to_unsigned(1443, 12), 1067 => to_unsigned(3444, 12), 1068 => to_unsigned(3340, 12), 1069 => to_unsigned(1677, 12), 1070 => to_unsigned(1655, 12), 1071 => to_unsigned(3199, 12), 1072 => to_unsigned(1911, 12), 1073 => to_unsigned(3835, 12), 1074 => to_unsigned(366, 12), 1075 => to_unsigned(2351, 12), 1076 => to_unsigned(2473, 12), 1077 => to_unsigned(115, 12), 1078 => to_unsigned(3857, 12), 1079 => to_unsigned(3747, 12), 1080 => to_unsigned(806, 12), 1081 => to_unsigned(1211, 12), 1082 => to_unsigned(3747, 12), 1083 => to_unsigned(1006, 12), 1084 => to_unsigned(610, 12), 1085 => to_unsigned(3293, 12), 1086 => to_unsigned(3111, 12), 1087 => to_unsigned(2993, 12), 1088 => to_unsigned(1464, 12), 1089 => to_unsigned(3165, 12), 1090 => to_unsigned(1109, 12), 1091 => to_unsigned(3722, 12), 1092 => to_unsigned(2123, 12), 1093 => to_unsigned(1637, 12), 1094 => to_unsigned(3188, 12), 1095 => to_unsigned(620, 12), 1096 => to_unsigned(1607, 12), 1097 => to_unsigned(2429, 12), 1098 => to_unsigned(2837, 12), 1099 => to_unsigned(520, 12), 1100 => to_unsigned(1619, 12), 1101 => to_unsigned(526, 12), 1102 => to_unsigned(2986, 12), 1103 => to_unsigned(1303, 12), 1104 => to_unsigned(501, 12), 1105 => to_unsigned(284, 12), 1106 => to_unsigned(1562, 12), 1107 => to_unsigned(3290, 12), 1108 => to_unsigned(715, 12), 1109 => to_unsigned(1526, 12), 1110 => to_unsigned(2020, 12), 1111 => to_unsigned(3088, 12), 1112 => to_unsigned(2619, 12), 1113 => to_unsigned(3248, 12), 1114 => to_unsigned(174, 12), 1115 => to_unsigned(3738, 12), 1116 => to_unsigned(1152, 12), 1117 => to_unsigned(2299, 12), 1118 => to_unsigned(688, 12), 1119 => to_unsigned(3771, 12), 1120 => to_unsigned(1196, 12), 1121 => to_unsigned(3620, 12), 1122 => to_unsigned(3362, 12), 1123 => to_unsigned(3230, 12), 1124 => to_unsigned(3959, 12), 1125 => to_unsigned(1498, 12), 1126 => to_unsigned(3238, 12), 1127 => to_unsigned(693, 12), 1128 => to_unsigned(1303, 12), 1129 => to_unsigned(839, 12), 1130 => to_unsigned(1864, 12), 1131 => to_unsigned(2325, 12), 1132 => to_unsigned(821, 12), 1133 => to_unsigned(3125, 12), 1134 => to_unsigned(3659, 12), 1135 => to_unsigned(1855, 12), 1136 => to_unsigned(1104, 12), 1137 => to_unsigned(1118, 12), 1138 => to_unsigned(3742, 12), 1139 => to_unsigned(2782, 12), 1140 => to_unsigned(3002, 12), 1141 => to_unsigned(3394, 12), 1142 => to_unsigned(3976, 12), 1143 => to_unsigned(4015, 12), 1144 => to_unsigned(2395, 12), 1145 => to_unsigned(3101, 12), 1146 => to_unsigned(1742, 12), 1147 => to_unsigned(1842, 12), 1148 => to_unsigned(693, 12), 1149 => to_unsigned(3372, 12), 1150 => to_unsigned(2778, 12), 1151 => to_unsigned(379, 12), 1152 => to_unsigned(248, 12), 1153 => to_unsigned(562, 12), 1154 => to_unsigned(1765, 12), 1155 => to_unsigned(495, 12), 1156 => to_unsigned(2748, 12), 1157 => to_unsigned(552, 12), 1158 => to_unsigned(636, 12), 1159 => to_unsigned(585, 12), 1160 => to_unsigned(3879, 12), 1161 => to_unsigned(3023, 12), 1162 => to_unsigned(508, 12), 1163 => to_unsigned(821, 12), 1164 => to_unsigned(25, 12), 1165 => to_unsigned(2683, 12), 1166 => to_unsigned(182, 12), 1167 => to_unsigned(3953, 12), 1168 => to_unsigned(3818, 12), 1169 => to_unsigned(1883, 12), 1170 => to_unsigned(959, 12), 1171 => to_unsigned(2127, 12), 1172 => to_unsigned(2333, 12), 1173 => to_unsigned(2788, 12), 1174 => to_unsigned(3937, 12), 1175 => to_unsigned(1352, 12), 1176 => to_unsigned(2523, 12), 1177 => to_unsigned(2673, 12), 1178 => to_unsigned(358, 12), 1179 => to_unsigned(3394, 12), 1180 => to_unsigned(2832, 12), 1181 => to_unsigned(3461, 12), 1182 => to_unsigned(272, 12), 1183 => to_unsigned(2678, 12), 1184 => to_unsigned(3829, 12), 1185 => to_unsigned(443, 12), 1186 => to_unsigned(2509, 12), 1187 => to_unsigned(1086, 12), 1188 => to_unsigned(2166, 12), 1189 => to_unsigned(3792, 12), 1190 => to_unsigned(319, 12), 1191 => to_unsigned(442, 12), 1192 => to_unsigned(2520, 12), 1193 => to_unsigned(198, 12), 1194 => to_unsigned(903, 12), 1195 => to_unsigned(44, 12), 1196 => to_unsigned(310, 12), 1197 => to_unsigned(2516, 12), 1198 => to_unsigned(2713, 12), 1199 => to_unsigned(1726, 12), 1200 => to_unsigned(599, 12), 1201 => to_unsigned(2743, 12), 1202 => to_unsigned(2896, 12), 1203 => to_unsigned(1946, 12), 1204 => to_unsigned(3750, 12), 1205 => to_unsigned(2169, 12), 1206 => to_unsigned(980, 12), 1207 => to_unsigned(3513, 12), 1208 => to_unsigned(3682, 12), 1209 => to_unsigned(3212, 12), 1210 => to_unsigned(1912, 12), 1211 => to_unsigned(436, 12), 1212 => to_unsigned(562, 12), 1213 => to_unsigned(3193, 12), 1214 => to_unsigned(3871, 12), 1215 => to_unsigned(1217, 12), 1216 => to_unsigned(3525, 12), 1217 => to_unsigned(2933, 12), 1218 => to_unsigned(4085, 12), 1219 => to_unsigned(1507, 12), 1220 => to_unsigned(941, 12), 1221 => to_unsigned(393, 12), 1222 => to_unsigned(2226, 12), 1223 => to_unsigned(1579, 12), 1224 => to_unsigned(3184, 12), 1225 => to_unsigned(2649, 12), 1226 => to_unsigned(148, 12), 1227 => to_unsigned(2347, 12), 1228 => to_unsigned(1882, 12), 1229 => to_unsigned(2489, 12), 1230 => to_unsigned(1236, 12), 1231 => to_unsigned(125, 12), 1232 => to_unsigned(2915, 12), 1233 => to_unsigned(1853, 12), 1234 => to_unsigned(1516, 12), 1235 => to_unsigned(1982, 12), 1236 => to_unsigned(2996, 12), 1237 => to_unsigned(3906, 12), 1238 => to_unsigned(588, 12), 1239 => to_unsigned(1681, 12), 1240 => to_unsigned(1301, 12), 1241 => to_unsigned(3366, 12), 1242 => to_unsigned(3555, 12), 1243 => to_unsigned(3197, 12), 1244 => to_unsigned(1536, 12), 1245 => to_unsigned(2379, 12), 1246 => to_unsigned(1231, 12), 1247 => to_unsigned(690, 12), 1248 => to_unsigned(413, 12), 1249 => to_unsigned(2651, 12), 1250 => to_unsigned(2917, 12), 1251 => to_unsigned(2353, 12), 1252 => to_unsigned(1668, 12), 1253 => to_unsigned(3002, 12), 1254 => to_unsigned(3692, 12), 1255 => to_unsigned(3713, 12), 1256 => to_unsigned(3449, 12), 1257 => to_unsigned(978, 12), 1258 => to_unsigned(2446, 12), 1259 => to_unsigned(2374, 12), 1260 => to_unsigned(1186, 12), 1261 => to_unsigned(194, 12), 1262 => to_unsigned(1695, 12), 1263 => to_unsigned(3183, 12), 1264 => to_unsigned(1153, 12), 1265 => to_unsigned(2361, 12), 1266 => to_unsigned(3256, 12), 1267 => to_unsigned(3212, 12), 1268 => to_unsigned(172, 12), 1269 => to_unsigned(109, 12), 1270 => to_unsigned(2274, 12), 1271 => to_unsigned(1307, 12), 1272 => to_unsigned(2513, 12), 1273 => to_unsigned(244, 12), 1274 => to_unsigned(739, 12), 1275 => to_unsigned(3964, 12), 1276 => to_unsigned(1231, 12), 1277 => to_unsigned(3035, 12), 1278 => to_unsigned(3236, 12), 1279 => to_unsigned(3597, 12), 1280 => to_unsigned(3051, 12), 1281 => to_unsigned(397, 12), 1282 => to_unsigned(2216, 12), 1283 => to_unsigned(1368, 12), 1284 => to_unsigned(1483, 12), 1285 => to_unsigned(3487, 12), 1286 => to_unsigned(3560, 12), 1287 => to_unsigned(1642, 12), 1288 => to_unsigned(1304, 12), 1289 => to_unsigned(790, 12), 1290 => to_unsigned(4020, 12), 1291 => to_unsigned(309, 12), 1292 => to_unsigned(4002, 12), 1293 => to_unsigned(925, 12), 1294 => to_unsigned(2770, 12), 1295 => to_unsigned(1487, 12), 1296 => to_unsigned(1226, 12), 1297 => to_unsigned(3622, 12), 1298 => to_unsigned(1482, 12), 1299 => to_unsigned(3662, 12), 1300 => to_unsigned(1496, 12), 1301 => to_unsigned(1775, 12), 1302 => to_unsigned(1986, 12), 1303 => to_unsigned(2941, 12), 1304 => to_unsigned(3956, 12), 1305 => to_unsigned(590, 12), 1306 => to_unsigned(1391, 12), 1307 => to_unsigned(3195, 12), 1308 => to_unsigned(996, 12), 1309 => to_unsigned(1887, 12), 1310 => to_unsigned(2297, 12), 1311 => to_unsigned(1242, 12), 1312 => to_unsigned(3834, 12), 1313 => to_unsigned(1899, 12), 1314 => to_unsigned(3612, 12), 1315 => to_unsigned(625, 12), 1316 => to_unsigned(2334, 12), 1317 => to_unsigned(2709, 12), 1318 => to_unsigned(3935, 12), 1319 => to_unsigned(1233, 12), 1320 => to_unsigned(2431, 12), 1321 => to_unsigned(1942, 12), 1322 => to_unsigned(1157, 12), 1323 => to_unsigned(2460, 12), 1324 => to_unsigned(3597, 12), 1325 => to_unsigned(979, 12), 1326 => to_unsigned(4018, 12), 1327 => to_unsigned(1345, 12), 1328 => to_unsigned(3072, 12), 1329 => to_unsigned(23, 12), 1330 => to_unsigned(874, 12), 1331 => to_unsigned(3917, 12), 1332 => to_unsigned(929, 12), 1333 => to_unsigned(2763, 12), 1334 => to_unsigned(1227, 12), 1335 => to_unsigned(2489, 12), 1336 => to_unsigned(909, 12), 1337 => to_unsigned(2243, 12), 1338 => to_unsigned(3179, 12), 1339 => to_unsigned(2950, 12), 1340 => to_unsigned(446, 12), 1341 => to_unsigned(3480, 12), 1342 => to_unsigned(2011, 12), 1343 => to_unsigned(3571, 12), 1344 => to_unsigned(3253, 12), 1345 => to_unsigned(477, 12), 1346 => to_unsigned(1361, 12), 1347 => to_unsigned(2574, 12), 1348 => to_unsigned(2543, 12), 1349 => to_unsigned(2525, 12), 1350 => to_unsigned(2080, 12), 1351 => to_unsigned(1205, 12), 1352 => to_unsigned(5, 12), 1353 => to_unsigned(3084, 12), 1354 => to_unsigned(3149, 12), 1355 => to_unsigned(2063, 12), 1356 => to_unsigned(2338, 12), 1357 => to_unsigned(3787, 12), 1358 => to_unsigned(239, 12), 1359 => to_unsigned(1200, 12), 1360 => to_unsigned(3755, 12), 1361 => to_unsigned(1391, 12), 1362 => to_unsigned(3176, 12), 1363 => to_unsigned(2176, 12), 1364 => to_unsigned(2114, 12), 1365 => to_unsigned(3025, 12), 1366 => to_unsigned(530, 12), 1367 => to_unsigned(1883, 12), 1368 => to_unsigned(3357, 12), 1369 => to_unsigned(3693, 12), 1370 => to_unsigned(3716, 12), 1371 => to_unsigned(2267, 12), 1372 => to_unsigned(849, 12), 1373 => to_unsigned(79, 12), 1374 => to_unsigned(3957, 12), 1375 => to_unsigned(2446, 12), 1376 => to_unsigned(2037, 12), 1377 => to_unsigned(3749, 12), 1378 => to_unsigned(3572, 12), 1379 => to_unsigned(2176, 12), 1380 => to_unsigned(1733, 12), 1381 => to_unsigned(3763, 12), 1382 => to_unsigned(2076, 12), 1383 => to_unsigned(2174, 12), 1384 => to_unsigned(4004, 12), 1385 => to_unsigned(801, 12), 1386 => to_unsigned(3005, 12), 1387 => to_unsigned(378, 12), 1388 => to_unsigned(180, 12), 1389 => to_unsigned(989, 12), 1390 => to_unsigned(1793, 12), 1391 => to_unsigned(3950, 12), 1392 => to_unsigned(2009, 12), 1393 => to_unsigned(301, 12), 1394 => to_unsigned(443, 12), 1395 => to_unsigned(2731, 12), 1396 => to_unsigned(3602, 12), 1397 => to_unsigned(600, 12), 1398 => to_unsigned(1669, 12), 1399 => to_unsigned(963, 12), 1400 => to_unsigned(1545, 12), 1401 => to_unsigned(3002, 12), 1402 => to_unsigned(3401, 12), 1403 => to_unsigned(1402, 12), 1404 => to_unsigned(3182, 12), 1405 => to_unsigned(1733, 12), 1406 => to_unsigned(1542, 12), 1407 => to_unsigned(1026, 12), 1408 => to_unsigned(1096, 12), 1409 => to_unsigned(2606, 12), 1410 => to_unsigned(1056, 12), 1411 => to_unsigned(764, 12), 1412 => to_unsigned(29, 12), 1413 => to_unsigned(614, 12), 1414 => to_unsigned(1046, 12), 1415 => to_unsigned(208, 12), 1416 => to_unsigned(2358, 12), 1417 => to_unsigned(246, 12), 1418 => to_unsigned(157, 12), 1419 => to_unsigned(3926, 12), 1420 => to_unsigned(401, 12), 1421 => to_unsigned(443, 12), 1422 => to_unsigned(1853, 12), 1423 => to_unsigned(3945, 12), 1424 => to_unsigned(508, 12), 1425 => to_unsigned(3106, 12), 1426 => to_unsigned(1066, 12), 1427 => to_unsigned(2143, 12), 1428 => to_unsigned(2740, 12), 1429 => to_unsigned(844, 12), 1430 => to_unsigned(1186, 12), 1431 => to_unsigned(214, 12), 1432 => to_unsigned(1491, 12), 1433 => to_unsigned(2882, 12), 1434 => to_unsigned(4055, 12), 1435 => to_unsigned(2177, 12), 1436 => to_unsigned(2490, 12), 1437 => to_unsigned(2010, 12), 1438 => to_unsigned(3895, 12), 1439 => to_unsigned(3325, 12), 1440 => to_unsigned(1186, 12), 1441 => to_unsigned(2133, 12), 1442 => to_unsigned(1293, 12), 1443 => to_unsigned(183, 12), 1444 => to_unsigned(2259, 12), 1445 => to_unsigned(1559, 12), 1446 => to_unsigned(3621, 12), 1447 => to_unsigned(285, 12), 1448 => to_unsigned(626, 12), 1449 => to_unsigned(4033, 12), 1450 => to_unsigned(1926, 12), 1451 => to_unsigned(761, 12), 1452 => to_unsigned(66, 12), 1453 => to_unsigned(2140, 12), 1454 => to_unsigned(2818, 12), 1455 => to_unsigned(562, 12), 1456 => to_unsigned(1846, 12), 1457 => to_unsigned(521, 12), 1458 => to_unsigned(3013, 12), 1459 => to_unsigned(361, 12), 1460 => to_unsigned(2151, 12), 1461 => to_unsigned(601, 12), 1462 => to_unsigned(1812, 12), 1463 => to_unsigned(2524, 12), 1464 => to_unsigned(992, 12), 1465 => to_unsigned(3894, 12), 1466 => to_unsigned(3820, 12), 1467 => to_unsigned(3754, 12), 1468 => to_unsigned(346, 12), 1469 => to_unsigned(110, 12), 1470 => to_unsigned(2961, 12), 1471 => to_unsigned(2755, 12), 1472 => to_unsigned(1599, 12), 1473 => to_unsigned(3610, 12), 1474 => to_unsigned(2126, 12), 1475 => to_unsigned(1404, 12), 1476 => to_unsigned(728, 12), 1477 => to_unsigned(3168, 12), 1478 => to_unsigned(1244, 12), 1479 => to_unsigned(3645, 12), 1480 => to_unsigned(692, 12), 1481 => to_unsigned(1171, 12), 1482 => to_unsigned(2980, 12), 1483 => to_unsigned(875, 12), 1484 => to_unsigned(3421, 12), 1485 => to_unsigned(3590, 12), 1486 => to_unsigned(2408, 12), 1487 => to_unsigned(1634, 12), 1488 => to_unsigned(1006, 12), 1489 => to_unsigned(3616, 12), 1490 => to_unsigned(2046, 12), 1491 => to_unsigned(2787, 12), 1492 => to_unsigned(959, 12), 1493 => to_unsigned(894, 12), 1494 => to_unsigned(1628, 12), 1495 => to_unsigned(212, 12), 1496 => to_unsigned(3477, 12), 1497 => to_unsigned(1899, 12), 1498 => to_unsigned(399, 12), 1499 => to_unsigned(3740, 12), 1500 => to_unsigned(154, 12), 1501 => to_unsigned(2315, 12), 1502 => to_unsigned(2827, 12), 1503 => to_unsigned(3205, 12), 1504 => to_unsigned(1144, 12), 1505 => to_unsigned(1295, 12), 1506 => to_unsigned(3618, 12), 1507 => to_unsigned(3661, 12), 1508 => to_unsigned(1867, 12), 1509 => to_unsigned(1655, 12), 1510 => to_unsigned(328, 12), 1511 => to_unsigned(1898, 12), 1512 => to_unsigned(2409, 12), 1513 => to_unsigned(537, 12), 1514 => to_unsigned(19, 12), 1515 => to_unsigned(2757, 12), 1516 => to_unsigned(627, 12), 1517 => to_unsigned(2112, 12), 1518 => to_unsigned(3532, 12), 1519 => to_unsigned(2697, 12), 1520 => to_unsigned(2176, 12), 1521 => to_unsigned(1591, 12), 1522 => to_unsigned(802, 12), 1523 => to_unsigned(3844, 12), 1524 => to_unsigned(2288, 12), 1525 => to_unsigned(3593, 12), 1526 => to_unsigned(3819, 12), 1527 => to_unsigned(1865, 12), 1528 => to_unsigned(3889, 12), 1529 => to_unsigned(2926, 12), 1530 => to_unsigned(3978, 12), 1531 => to_unsigned(491, 12), 1532 => to_unsigned(2279, 12), 1533 => to_unsigned(767, 12), 1534 => to_unsigned(4087, 12), 1535 => to_unsigned(1493, 12), 1536 => to_unsigned(3771, 12), 1537 => to_unsigned(1705, 12), 1538 => to_unsigned(296, 12), 1539 => to_unsigned(880, 12), 1540 => to_unsigned(1693, 12), 1541 => to_unsigned(700, 12), 1542 => to_unsigned(1502, 12), 1543 => to_unsigned(3949, 12), 1544 => to_unsigned(1541, 12), 1545 => to_unsigned(2900, 12), 1546 => to_unsigned(1682, 12), 1547 => to_unsigned(149, 12), 1548 => to_unsigned(3191, 12), 1549 => to_unsigned(2754, 12), 1550 => to_unsigned(2579, 12), 1551 => to_unsigned(1793, 12), 1552 => to_unsigned(918, 12), 1553 => to_unsigned(1648, 12), 1554 => to_unsigned(1833, 12), 1555 => to_unsigned(1802, 12), 1556 => to_unsigned(916, 12), 1557 => to_unsigned(2750, 12), 1558 => to_unsigned(1607, 12), 1559 => to_unsigned(112, 12), 1560 => to_unsigned(3383, 12), 1561 => to_unsigned(2650, 12), 1562 => to_unsigned(2711, 12), 1563 => to_unsigned(2088, 12), 1564 => to_unsigned(3690, 12), 1565 => to_unsigned(1635, 12), 1566 => to_unsigned(3311, 12), 1567 => to_unsigned(3449, 12), 1568 => to_unsigned(584, 12), 1569 => to_unsigned(2466, 12), 1570 => to_unsigned(2715, 12), 1571 => to_unsigned(4, 12), 1572 => to_unsigned(2500, 12), 1573 => to_unsigned(3602, 12), 1574 => to_unsigned(2697, 12), 1575 => to_unsigned(3304, 12), 1576 => to_unsigned(2951, 12), 1577 => to_unsigned(2994, 12), 1578 => to_unsigned(3102, 12), 1579 => to_unsigned(1486, 12), 1580 => to_unsigned(1364, 12), 1581 => to_unsigned(189, 12), 1582 => to_unsigned(253, 12), 1583 => to_unsigned(315, 12), 1584 => to_unsigned(1014, 12), 1585 => to_unsigned(1237, 12), 1586 => to_unsigned(1818, 12), 1587 => to_unsigned(3829, 12), 1588 => to_unsigned(99, 12), 1589 => to_unsigned(2247, 12), 1590 => to_unsigned(238, 12), 1591 => to_unsigned(198, 12), 1592 => to_unsigned(2443, 12), 1593 => to_unsigned(2268, 12), 1594 => to_unsigned(1786, 12), 1595 => to_unsigned(2671, 12), 1596 => to_unsigned(423, 12), 1597 => to_unsigned(3911, 12), 1598 => to_unsigned(671, 12), 1599 => to_unsigned(497, 12), 1600 => to_unsigned(1659, 12), 1601 => to_unsigned(443, 12), 1602 => to_unsigned(79, 12), 1603 => to_unsigned(1930, 12), 1604 => to_unsigned(2460, 12), 1605 => to_unsigned(2164, 12), 1606 => to_unsigned(3462, 12), 1607 => to_unsigned(2905, 12), 1608 => to_unsigned(2842, 12), 1609 => to_unsigned(54, 12), 1610 => to_unsigned(273, 12), 1611 => to_unsigned(1511, 12), 1612 => to_unsigned(2060, 12), 1613 => to_unsigned(3674, 12), 1614 => to_unsigned(3427, 12), 1615 => to_unsigned(578, 12), 1616 => to_unsigned(3837, 12), 1617 => to_unsigned(67, 12), 1618 => to_unsigned(668, 12), 1619 => to_unsigned(3523, 12), 1620 => to_unsigned(354, 12), 1621 => to_unsigned(2939, 12), 1622 => to_unsigned(2998, 12), 1623 => to_unsigned(2068, 12), 1624 => to_unsigned(1264, 12), 1625 => to_unsigned(257, 12), 1626 => to_unsigned(3687, 12), 1627 => to_unsigned(2260, 12), 1628 => to_unsigned(222, 12), 1629 => to_unsigned(3488, 12), 1630 => to_unsigned(1693, 12), 1631 => to_unsigned(1039, 12), 1632 => to_unsigned(2054, 12), 1633 => to_unsigned(809, 12), 1634 => to_unsigned(1290, 12), 1635 => to_unsigned(1498, 12), 1636 => to_unsigned(3845, 12), 1637 => to_unsigned(2831, 12), 1638 => to_unsigned(220, 12), 1639 => to_unsigned(1859, 12), 1640 => to_unsigned(2173, 12), 1641 => to_unsigned(2875, 12), 1642 => to_unsigned(2613, 12), 1643 => to_unsigned(2007, 12), 1644 => to_unsigned(3834, 12), 1645 => to_unsigned(1224, 12), 1646 => to_unsigned(2986, 12), 1647 => to_unsigned(2139, 12), 1648 => to_unsigned(1656, 12), 1649 => to_unsigned(37, 12), 1650 => to_unsigned(3609, 12), 1651 => to_unsigned(114, 12), 1652 => to_unsigned(1681, 12), 1653 => to_unsigned(2400, 12), 1654 => to_unsigned(3031, 12), 1655 => to_unsigned(1102, 12), 1656 => to_unsigned(2767, 12), 1657 => to_unsigned(1095, 12), 1658 => to_unsigned(3285, 12), 1659 => to_unsigned(3229, 12), 1660 => to_unsigned(636, 12), 1661 => to_unsigned(2593, 12), 1662 => to_unsigned(455, 12), 1663 => to_unsigned(4055, 12), 1664 => to_unsigned(387, 12), 1665 => to_unsigned(3843, 12), 1666 => to_unsigned(258, 12), 1667 => to_unsigned(1891, 12), 1668 => to_unsigned(2948, 12), 1669 => to_unsigned(2238, 12), 1670 => to_unsigned(794, 12), 1671 => to_unsigned(3465, 12), 1672 => to_unsigned(591, 12), 1673 => to_unsigned(2048, 12), 1674 => to_unsigned(3920, 12), 1675 => to_unsigned(1496, 12), 1676 => to_unsigned(1468, 12), 1677 => to_unsigned(2804, 12), 1678 => to_unsigned(840, 12), 1679 => to_unsigned(1937, 12), 1680 => to_unsigned(1026, 12), 1681 => to_unsigned(3108, 12), 1682 => to_unsigned(1035, 12), 1683 => to_unsigned(1352, 12), 1684 => to_unsigned(2487, 12), 1685 => to_unsigned(786, 12), 1686 => to_unsigned(2714, 12), 1687 => to_unsigned(2967, 12), 1688 => to_unsigned(3980, 12), 1689 => to_unsigned(1939, 12), 1690 => to_unsigned(2983, 12), 1691 => to_unsigned(1247, 12), 1692 => to_unsigned(2813, 12), 1693 => to_unsigned(774, 12), 1694 => to_unsigned(1586, 12), 1695 => to_unsigned(985, 12), 1696 => to_unsigned(1785, 12), 1697 => to_unsigned(1292, 12), 1698 => to_unsigned(832, 12), 1699 => to_unsigned(1594, 12), 1700 => to_unsigned(418, 12), 1701 => to_unsigned(1955, 12), 1702 => to_unsigned(1270, 12), 1703 => to_unsigned(680, 12), 1704 => to_unsigned(1022, 12), 1705 => to_unsigned(3458, 12), 1706 => to_unsigned(2278, 12), 1707 => to_unsigned(192, 12), 1708 => to_unsigned(1604, 12), 1709 => to_unsigned(1093, 12), 1710 => to_unsigned(3939, 12), 1711 => to_unsigned(484, 12), 1712 => to_unsigned(3145, 12), 1713 => to_unsigned(1197, 12), 1714 => to_unsigned(1873, 12), 1715 => to_unsigned(2781, 12), 1716 => to_unsigned(1344, 12), 1717 => to_unsigned(2572, 12), 1718 => to_unsigned(180, 12), 1719 => to_unsigned(95, 12), 1720 => to_unsigned(3823, 12), 1721 => to_unsigned(3090, 12), 1722 => to_unsigned(835, 12), 1723 => to_unsigned(1549, 12), 1724 => to_unsigned(1538, 12), 1725 => to_unsigned(1232, 12), 1726 => to_unsigned(277, 12), 1727 => to_unsigned(3241, 12), 1728 => to_unsigned(3160, 12), 1729 => to_unsigned(302, 12), 1730 => to_unsigned(3464, 12), 1731 => to_unsigned(434, 12), 1732 => to_unsigned(304, 12), 1733 => to_unsigned(1519, 12), 1734 => to_unsigned(3946, 12), 1735 => to_unsigned(2980, 12), 1736 => to_unsigned(2107, 12), 1737 => to_unsigned(2404, 12), 1738 => to_unsigned(4059, 12), 1739 => to_unsigned(2650, 12), 1740 => to_unsigned(3982, 12), 1741 => to_unsigned(2472, 12), 1742 => to_unsigned(2692, 12), 1743 => to_unsigned(547, 12), 1744 => to_unsigned(1090, 12), 1745 => to_unsigned(2451, 12), 1746 => to_unsigned(2076, 12), 1747 => to_unsigned(1042, 12), 1748 => to_unsigned(3660, 12), 1749 => to_unsigned(2839, 12), 1750 => to_unsigned(1871, 12), 1751 => to_unsigned(110, 12), 1752 => to_unsigned(1707, 12), 1753 => to_unsigned(2191, 12), 1754 => to_unsigned(3454, 12), 1755 => to_unsigned(3554, 12), 1756 => to_unsigned(1126, 12), 1757 => to_unsigned(1837, 12), 1758 => to_unsigned(97, 12), 1759 => to_unsigned(1780, 12), 1760 => to_unsigned(443, 12), 1761 => to_unsigned(2714, 12), 1762 => to_unsigned(3097, 12), 1763 => to_unsigned(1191, 12), 1764 => to_unsigned(3265, 12), 1765 => to_unsigned(3775, 12), 1766 => to_unsigned(1194, 12), 1767 => to_unsigned(1874, 12), 1768 => to_unsigned(621, 12), 1769 => to_unsigned(971, 12), 1770 => to_unsigned(1317, 12), 1771 => to_unsigned(3132, 12), 1772 => to_unsigned(720, 12), 1773 => to_unsigned(3938, 12), 1774 => to_unsigned(2283, 12), 1775 => to_unsigned(1308, 12), 1776 => to_unsigned(2956, 12), 1777 => to_unsigned(770, 12), 1778 => to_unsigned(2350, 12), 1779 => to_unsigned(1130, 12), 1780 => to_unsigned(3501, 12), 1781 => to_unsigned(3338, 12), 1782 => to_unsigned(2468, 12), 1783 => to_unsigned(3144, 12), 1784 => to_unsigned(3507, 12), 1785 => to_unsigned(1978, 12), 1786 => to_unsigned(2547, 12), 1787 => to_unsigned(3071, 12), 1788 => to_unsigned(3959, 12), 1789 => to_unsigned(1808, 12), 1790 => to_unsigned(1406, 12), 1791 => to_unsigned(1840, 12), 1792 => to_unsigned(2840, 12), 1793 => to_unsigned(3801, 12), 1794 => to_unsigned(3300, 12), 1795 => to_unsigned(1151, 12), 1796 => to_unsigned(2781, 12), 1797 => to_unsigned(768, 12), 1798 => to_unsigned(957, 12), 1799 => to_unsigned(2016, 12), 1800 => to_unsigned(1194, 12), 1801 => to_unsigned(899, 12), 1802 => to_unsigned(944, 12), 1803 => to_unsigned(4008, 12), 1804 => to_unsigned(3048, 12), 1805 => to_unsigned(2801, 12), 1806 => to_unsigned(1438, 12), 1807 => to_unsigned(425, 12), 1808 => to_unsigned(2809, 12), 1809 => to_unsigned(1691, 12), 1810 => to_unsigned(458, 12), 1811 => to_unsigned(2617, 12), 1812 => to_unsigned(3775, 12), 1813 => to_unsigned(1225, 12), 1814 => to_unsigned(930, 12), 1815 => to_unsigned(2601, 12), 1816 => to_unsigned(2200, 12), 1817 => to_unsigned(1018, 12), 1818 => to_unsigned(1424, 12), 1819 => to_unsigned(2311, 12), 1820 => to_unsigned(3376, 12), 1821 => to_unsigned(1778, 12), 1822 => to_unsigned(1314, 12), 1823 => to_unsigned(1359, 12), 1824 => to_unsigned(68, 12), 1825 => to_unsigned(1914, 12), 1826 => to_unsigned(1894, 12), 1827 => to_unsigned(3752, 12), 1828 => to_unsigned(2183, 12), 1829 => to_unsigned(3498, 12), 1830 => to_unsigned(291, 12), 1831 => to_unsigned(3828, 12), 1832 => to_unsigned(971, 12), 1833 => to_unsigned(3788, 12), 1834 => to_unsigned(2272, 12), 1835 => to_unsigned(3955, 12), 1836 => to_unsigned(1771, 12), 1837 => to_unsigned(2503, 12), 1838 => to_unsigned(680, 12), 1839 => to_unsigned(3304, 12), 1840 => to_unsigned(1069, 12), 1841 => to_unsigned(207, 12), 1842 => to_unsigned(593, 12), 1843 => to_unsigned(3530, 12), 1844 => to_unsigned(2426, 12), 1845 => to_unsigned(1755, 12), 1846 => to_unsigned(2160, 12), 1847 => to_unsigned(2194, 12), 1848 => to_unsigned(3830, 12), 1849 => to_unsigned(3185, 12), 1850 => to_unsigned(1398, 12), 1851 => to_unsigned(423, 12), 1852 => to_unsigned(3777, 12), 1853 => to_unsigned(911, 12), 1854 => to_unsigned(749, 12), 1855 => to_unsigned(252, 12), 1856 => to_unsigned(3573, 12), 1857 => to_unsigned(4026, 12), 1858 => to_unsigned(1495, 12), 1859 => to_unsigned(3654, 12), 1860 => to_unsigned(4022, 12), 1861 => to_unsigned(1693, 12), 1862 => to_unsigned(3277, 12), 1863 => to_unsigned(863, 12), 1864 => to_unsigned(1349, 12), 1865 => to_unsigned(3150, 12), 1866 => to_unsigned(1755, 12), 1867 => to_unsigned(1697, 12), 1868 => to_unsigned(797, 12), 1869 => to_unsigned(3451, 12), 1870 => to_unsigned(3610, 12), 1871 => to_unsigned(1571, 12), 1872 => to_unsigned(1144, 12), 1873 => to_unsigned(4084, 12), 1874 => to_unsigned(1304, 12), 1875 => to_unsigned(3771, 12), 1876 => to_unsigned(3941, 12), 1877 => to_unsigned(902, 12), 1878 => to_unsigned(766, 12), 1879 => to_unsigned(1346, 12), 1880 => to_unsigned(36, 12), 1881 => to_unsigned(3569, 12), 1882 => to_unsigned(3771, 12), 1883 => to_unsigned(956, 12), 1884 => to_unsigned(3822, 12), 1885 => to_unsigned(2871, 12), 1886 => to_unsigned(1188, 12), 1887 => to_unsigned(1295, 12), 1888 => to_unsigned(3869, 12), 1889 => to_unsigned(2780, 12), 1890 => to_unsigned(2470, 12), 1891 => to_unsigned(2180, 12), 1892 => to_unsigned(3544, 12), 1893 => to_unsigned(1917, 12), 1894 => to_unsigned(429, 12), 1895 => to_unsigned(996, 12), 1896 => to_unsigned(3329, 12), 1897 => to_unsigned(1883, 12), 1898 => to_unsigned(2502, 12), 1899 => to_unsigned(3744, 12), 1900 => to_unsigned(659, 12), 1901 => to_unsigned(3942, 12), 1902 => to_unsigned(3617, 12), 1903 => to_unsigned(375, 12), 1904 => to_unsigned(3885, 12), 1905 => to_unsigned(2928, 12), 1906 => to_unsigned(1924, 12), 1907 => to_unsigned(1010, 12), 1908 => to_unsigned(1219, 12), 1909 => to_unsigned(770, 12), 1910 => to_unsigned(2862, 12), 1911 => to_unsigned(3953, 12), 1912 => to_unsigned(1529, 12), 1913 => to_unsigned(3370, 12), 1914 => to_unsigned(2754, 12), 1915 => to_unsigned(892, 12), 1916 => to_unsigned(1569, 12), 1917 => to_unsigned(3785, 12), 1918 => to_unsigned(654, 12), 1919 => to_unsigned(2897, 12), 1920 => to_unsigned(1069, 12), 1921 => to_unsigned(973, 12), 1922 => to_unsigned(146, 12), 1923 => to_unsigned(804, 12), 1924 => to_unsigned(1402, 12), 1925 => to_unsigned(2450, 12), 1926 => to_unsigned(3957, 12), 1927 => to_unsigned(2518, 12), 1928 => to_unsigned(1935, 12), 1929 => to_unsigned(823, 12), 1930 => to_unsigned(3702, 12), 1931 => to_unsigned(462, 12), 1932 => to_unsigned(3037, 12), 1933 => to_unsigned(636, 12), 1934 => to_unsigned(3687, 12), 1935 => to_unsigned(3467, 12), 1936 => to_unsigned(2131, 12), 1937 => to_unsigned(989, 12), 1938 => to_unsigned(2353, 12), 1939 => to_unsigned(3900, 12), 1940 => to_unsigned(1128, 12), 1941 => to_unsigned(2692, 12), 1942 => to_unsigned(1947, 12), 1943 => to_unsigned(2936, 12), 1944 => to_unsigned(609, 12), 1945 => to_unsigned(1370, 12), 1946 => to_unsigned(2480, 12), 1947 => to_unsigned(500, 12), 1948 => to_unsigned(2766, 12), 1949 => to_unsigned(2822, 12), 1950 => to_unsigned(1393, 12), 1951 => to_unsigned(3394, 12), 1952 => to_unsigned(1288, 12), 1953 => to_unsigned(1152, 12), 1954 => to_unsigned(3116, 12), 1955 => to_unsigned(1008, 12), 1956 => to_unsigned(3391, 12), 1957 => to_unsigned(2316, 12), 1958 => to_unsigned(915, 12), 1959 => to_unsigned(2999, 12), 1960 => to_unsigned(1783, 12), 1961 => to_unsigned(2155, 12), 1962 => to_unsigned(1024, 12), 1963 => to_unsigned(1363, 12), 1964 => to_unsigned(1413, 12), 1965 => to_unsigned(3808, 12), 1966 => to_unsigned(2368, 12), 1967 => to_unsigned(3258, 12), 1968 => to_unsigned(2334, 12), 1969 => to_unsigned(1983, 12), 1970 => to_unsigned(2771, 12), 1971 => to_unsigned(3171, 12), 1972 => to_unsigned(635, 12), 1973 => to_unsigned(2935, 12), 1974 => to_unsigned(376, 12), 1975 => to_unsigned(155, 12), 1976 => to_unsigned(2253, 12), 1977 => to_unsigned(2449, 12), 1978 => to_unsigned(1957, 12), 1979 => to_unsigned(1201, 12), 1980 => to_unsigned(708, 12), 1981 => to_unsigned(221, 12), 1982 => to_unsigned(1553, 12), 1983 => to_unsigned(224, 12), 1984 => to_unsigned(2731, 12), 1985 => to_unsigned(3923, 12), 1986 => to_unsigned(2792, 12), 1987 => to_unsigned(2276, 12), 1988 => to_unsigned(2539, 12), 1989 => to_unsigned(1490, 12), 1990 => to_unsigned(71, 12), 1991 => to_unsigned(2534, 12), 1992 => to_unsigned(2642, 12), 1993 => to_unsigned(3713, 12), 1994 => to_unsigned(830, 12), 1995 => to_unsigned(50, 12), 1996 => to_unsigned(908, 12), 1997 => to_unsigned(2946, 12), 1998 => to_unsigned(3442, 12), 1999 => to_unsigned(3807, 12), 2000 => to_unsigned(1110, 12), 2001 => to_unsigned(817, 12), 2002 => to_unsigned(2953, 12), 2003 => to_unsigned(2990, 12), 2004 => to_unsigned(1012, 12), 2005 => to_unsigned(3958, 12), 2006 => to_unsigned(1007, 12), 2007 => to_unsigned(3107, 12), 2008 => to_unsigned(2266, 12), 2009 => to_unsigned(880, 12), 2010 => to_unsigned(1190, 12), 2011 => to_unsigned(1254, 12), 2012 => to_unsigned(1214, 12), 2013 => to_unsigned(755, 12), 2014 => to_unsigned(298, 12), 2015 => to_unsigned(1073, 12), 2016 => to_unsigned(3718, 12), 2017 => to_unsigned(2936, 12), 2018 => to_unsigned(1744, 12), 2019 => to_unsigned(3205, 12), 2020 => to_unsigned(2105, 12), 2021 => to_unsigned(2000, 12), 2022 => to_unsigned(2204, 12), 2023 => to_unsigned(2376, 12), 2024 => to_unsigned(2086, 12), 2025 => to_unsigned(1407, 12), 2026 => to_unsigned(2639, 12), 2027 => to_unsigned(937, 12), 2028 => to_unsigned(1081, 12), 2029 => to_unsigned(2295, 12), 2030 => to_unsigned(1451, 12), 2031 => to_unsigned(1495, 12), 2032 => to_unsigned(2972, 12), 2033 => to_unsigned(1709, 12), 2034 => to_unsigned(1028, 12), 2035 => to_unsigned(1744, 12), 2036 => to_unsigned(582, 12), 2037 => to_unsigned(3030, 12), 2038 => to_unsigned(1499, 12), 2039 => to_unsigned(3761, 12), 2040 => to_unsigned(2551, 12), 2041 => to_unsigned(815, 12), 2042 => to_unsigned(3949, 12), 2043 => to_unsigned(1523, 12), 2044 => to_unsigned(2796, 12), 2045 => to_unsigned(3382, 12), 2046 => to_unsigned(33, 12), 2047 => to_unsigned(1151, 12)),
            2 => (0 => to_unsigned(3226, 12), 1 => to_unsigned(3394, 12), 2 => to_unsigned(3577, 12), 3 => to_unsigned(1519, 12), 4 => to_unsigned(781, 12), 5 => to_unsigned(703, 12), 6 => to_unsigned(331, 12), 7 => to_unsigned(1934, 12), 8 => to_unsigned(2812, 12), 9 => to_unsigned(3082, 12), 10 => to_unsigned(2377, 12), 11 => to_unsigned(409, 12), 12 => to_unsigned(3722, 12), 13 => to_unsigned(3994, 12), 14 => to_unsigned(764, 12), 15 => to_unsigned(890, 12), 16 => to_unsigned(2321, 12), 17 => to_unsigned(2389, 12), 18 => to_unsigned(2211, 12), 19 => to_unsigned(930, 12), 20 => to_unsigned(2976, 12), 21 => to_unsigned(189, 12), 22 => to_unsigned(3002, 12), 23 => to_unsigned(2496, 12), 24 => to_unsigned(580, 12), 25 => to_unsigned(2831, 12), 26 => to_unsigned(2665, 12), 27 => to_unsigned(1817, 12), 28 => to_unsigned(3580, 12), 29 => to_unsigned(1340, 12), 30 => to_unsigned(1548, 12), 31 => to_unsigned(1074, 12), 32 => to_unsigned(1859, 12), 33 => to_unsigned(3992, 12), 34 => to_unsigned(2809, 12), 35 => to_unsigned(1603, 12), 36 => to_unsigned(2253, 12), 37 => to_unsigned(1077, 12), 38 => to_unsigned(1926, 12), 39 => to_unsigned(2597, 12), 40 => to_unsigned(967, 12), 41 => to_unsigned(2247, 12), 42 => to_unsigned(183, 12), 43 => to_unsigned(63, 12), 44 => to_unsigned(1841, 12), 45 => to_unsigned(3545, 12), 46 => to_unsigned(1033, 12), 47 => to_unsigned(2489, 12), 48 => to_unsigned(1479, 12), 49 => to_unsigned(3786, 12), 50 => to_unsigned(3238, 12), 51 => to_unsigned(975, 12), 52 => to_unsigned(1490, 12), 53 => to_unsigned(597, 12), 54 => to_unsigned(2594, 12), 55 => to_unsigned(931, 12), 56 => to_unsigned(1105, 12), 57 => to_unsigned(1343, 12), 58 => to_unsigned(3227, 12), 59 => to_unsigned(3671, 12), 60 => to_unsigned(2211, 12), 61 => to_unsigned(2517, 12), 62 => to_unsigned(745, 12), 63 => to_unsigned(1313, 12), 64 => to_unsigned(160, 12), 65 => to_unsigned(848, 12), 66 => to_unsigned(1383, 12), 67 => to_unsigned(1110, 12), 68 => to_unsigned(2123, 12), 69 => to_unsigned(3607, 12), 70 => to_unsigned(2651, 12), 71 => to_unsigned(3910, 12), 72 => to_unsigned(2437, 12), 73 => to_unsigned(232, 12), 74 => to_unsigned(1910, 12), 75 => to_unsigned(3278, 12), 76 => to_unsigned(1549, 12), 77 => to_unsigned(3377, 12), 78 => to_unsigned(2877, 12), 79 => to_unsigned(4079, 12), 80 => to_unsigned(2400, 12), 81 => to_unsigned(3713, 12), 82 => to_unsigned(2404, 12), 83 => to_unsigned(3106, 12), 84 => to_unsigned(1723, 12), 85 => to_unsigned(122, 12), 86 => to_unsigned(3584, 12), 87 => to_unsigned(1569, 12), 88 => to_unsigned(2314, 12), 89 => to_unsigned(3329, 12), 90 => to_unsigned(3659, 12), 91 => to_unsigned(2479, 12), 92 => to_unsigned(3313, 12), 93 => to_unsigned(3582, 12), 94 => to_unsigned(699, 12), 95 => to_unsigned(2658, 12), 96 => to_unsigned(2754, 12), 97 => to_unsigned(1708, 12), 98 => to_unsigned(3914, 12), 99 => to_unsigned(3748, 12), 100 => to_unsigned(1086, 12), 101 => to_unsigned(273, 12), 102 => to_unsigned(761, 12), 103 => to_unsigned(3305, 12), 104 => to_unsigned(3642, 12), 105 => to_unsigned(136, 12), 106 => to_unsigned(896, 12), 107 => to_unsigned(3196, 12), 108 => to_unsigned(290, 12), 109 => to_unsigned(3796, 12), 110 => to_unsigned(2471, 12), 111 => to_unsigned(1545, 12), 112 => to_unsigned(2722, 12), 113 => to_unsigned(1627, 12), 114 => to_unsigned(1266, 12), 115 => to_unsigned(4, 12), 116 => to_unsigned(4034, 12), 117 => to_unsigned(3851, 12), 118 => to_unsigned(1789, 12), 119 => to_unsigned(3958, 12), 120 => to_unsigned(3088, 12), 121 => to_unsigned(3790, 12), 122 => to_unsigned(2478, 12), 123 => to_unsigned(889, 12), 124 => to_unsigned(2338, 12), 125 => to_unsigned(3310, 12), 126 => to_unsigned(3285, 12), 127 => to_unsigned(2825, 12), 128 => to_unsigned(1943, 12), 129 => to_unsigned(174, 12), 130 => to_unsigned(30, 12), 131 => to_unsigned(3800, 12), 132 => to_unsigned(3007, 12), 133 => to_unsigned(1153, 12), 134 => to_unsigned(3552, 12), 135 => to_unsigned(3017, 12), 136 => to_unsigned(3265, 12), 137 => to_unsigned(67, 12), 138 => to_unsigned(198, 12), 139 => to_unsigned(502, 12), 140 => to_unsigned(2008, 12), 141 => to_unsigned(3516, 12), 142 => to_unsigned(1795, 12), 143 => to_unsigned(1205, 12), 144 => to_unsigned(1217, 12), 145 => to_unsigned(470, 12), 146 => to_unsigned(2931, 12), 147 => to_unsigned(1793, 12), 148 => to_unsigned(3328, 12), 149 => to_unsigned(694, 12), 150 => to_unsigned(2278, 12), 151 => to_unsigned(2124, 12), 152 => to_unsigned(2371, 12), 153 => to_unsigned(140, 12), 154 => to_unsigned(2487, 12), 155 => to_unsigned(102, 12), 156 => to_unsigned(2213, 12), 157 => to_unsigned(2830, 12), 158 => to_unsigned(2221, 12), 159 => to_unsigned(421, 12), 160 => to_unsigned(1975, 12), 161 => to_unsigned(2385, 12), 162 => to_unsigned(1330, 12), 163 => to_unsigned(870, 12), 164 => to_unsigned(551, 12), 165 => to_unsigned(72, 12), 166 => to_unsigned(173, 12), 167 => to_unsigned(3680, 12), 168 => to_unsigned(280, 12), 169 => to_unsigned(3233, 12), 170 => to_unsigned(245, 12), 171 => to_unsigned(309, 12), 172 => to_unsigned(3515, 12), 173 => to_unsigned(927, 12), 174 => to_unsigned(3457, 12), 175 => to_unsigned(2909, 12), 176 => to_unsigned(2468, 12), 177 => to_unsigned(305, 12), 178 => to_unsigned(2494, 12), 179 => to_unsigned(3827, 12), 180 => to_unsigned(2914, 12), 181 => to_unsigned(1770, 12), 182 => to_unsigned(3199, 12), 183 => to_unsigned(2085, 12), 184 => to_unsigned(3258, 12), 185 => to_unsigned(1649, 12), 186 => to_unsigned(3693, 12), 187 => to_unsigned(2692, 12), 188 => to_unsigned(480, 12), 189 => to_unsigned(3971, 12), 190 => to_unsigned(2430, 12), 191 => to_unsigned(1763, 12), 192 => to_unsigned(1934, 12), 193 => to_unsigned(2028, 12), 194 => to_unsigned(1725, 12), 195 => to_unsigned(3185, 12), 196 => to_unsigned(1156, 12), 197 => to_unsigned(2310, 12), 198 => to_unsigned(3315, 12), 199 => to_unsigned(748, 12), 200 => to_unsigned(766, 12), 201 => to_unsigned(2595, 12), 202 => to_unsigned(1143, 12), 203 => to_unsigned(3637, 12), 204 => to_unsigned(2684, 12), 205 => to_unsigned(1947, 12), 206 => to_unsigned(3133, 12), 207 => to_unsigned(3373, 12), 208 => to_unsigned(2312, 12), 209 => to_unsigned(4033, 12), 210 => to_unsigned(2603, 12), 211 => to_unsigned(3947, 12), 212 => to_unsigned(959, 12), 213 => to_unsigned(32, 12), 214 => to_unsigned(1047, 12), 215 => to_unsigned(4072, 12), 216 => to_unsigned(2713, 12), 217 => to_unsigned(2557, 12), 218 => to_unsigned(2417, 12), 219 => to_unsigned(1006, 12), 220 => to_unsigned(3650, 12), 221 => to_unsigned(501, 12), 222 => to_unsigned(3064, 12), 223 => to_unsigned(3107, 12), 224 => to_unsigned(2908, 12), 225 => to_unsigned(3787, 12), 226 => to_unsigned(562, 12), 227 => to_unsigned(3249, 12), 228 => to_unsigned(577, 12), 229 => to_unsigned(1573, 12), 230 => to_unsigned(1564, 12), 231 => to_unsigned(3973, 12), 232 => to_unsigned(3134, 12), 233 => to_unsigned(2913, 12), 234 => to_unsigned(1585, 12), 235 => to_unsigned(2906, 12), 236 => to_unsigned(520, 12), 237 => to_unsigned(3366, 12), 238 => to_unsigned(40, 12), 239 => to_unsigned(3852, 12), 240 => to_unsigned(3070, 12), 241 => to_unsigned(2511, 12), 242 => to_unsigned(3247, 12), 243 => to_unsigned(470, 12), 244 => to_unsigned(3082, 12), 245 => to_unsigned(2167, 12), 246 => to_unsigned(1571, 12), 247 => to_unsigned(275, 12), 248 => to_unsigned(2722, 12), 249 => to_unsigned(952, 12), 250 => to_unsigned(3337, 12), 251 => to_unsigned(1113, 12), 252 => to_unsigned(2686, 12), 253 => to_unsigned(1716, 12), 254 => to_unsigned(1478, 12), 255 => to_unsigned(935, 12), 256 => to_unsigned(1099, 12), 257 => to_unsigned(3212, 12), 258 => to_unsigned(4066, 12), 259 => to_unsigned(2464, 12), 260 => to_unsigned(1589, 12), 261 => to_unsigned(2170, 12), 262 => to_unsigned(2640, 12), 263 => to_unsigned(3011, 12), 264 => to_unsigned(2126, 12), 265 => to_unsigned(2276, 12), 266 => to_unsigned(3127, 12), 267 => to_unsigned(3281, 12), 268 => to_unsigned(2761, 12), 269 => to_unsigned(61, 12), 270 => to_unsigned(930, 12), 271 => to_unsigned(155, 12), 272 => to_unsigned(2204, 12), 273 => to_unsigned(3757, 12), 274 => to_unsigned(3594, 12), 275 => to_unsigned(3589, 12), 276 => to_unsigned(3807, 12), 277 => to_unsigned(719, 12), 278 => to_unsigned(3628, 12), 279 => to_unsigned(2637, 12), 280 => to_unsigned(3255, 12), 281 => to_unsigned(3270, 12), 282 => to_unsigned(1935, 12), 283 => to_unsigned(7, 12), 284 => to_unsigned(2156, 12), 285 => to_unsigned(850, 12), 286 => to_unsigned(293, 12), 287 => to_unsigned(2841, 12), 288 => to_unsigned(2619, 12), 289 => to_unsigned(3356, 12), 290 => to_unsigned(2866, 12), 291 => to_unsigned(2394, 12), 292 => to_unsigned(200, 12), 293 => to_unsigned(1327, 12), 294 => to_unsigned(2235, 12), 295 => to_unsigned(1437, 12), 296 => to_unsigned(147, 12), 297 => to_unsigned(1571, 12), 298 => to_unsigned(3442, 12), 299 => to_unsigned(57, 12), 300 => to_unsigned(419, 12), 301 => to_unsigned(925, 12), 302 => to_unsigned(2384, 12), 303 => to_unsigned(3524, 12), 304 => to_unsigned(739, 12), 305 => to_unsigned(2098, 12), 306 => to_unsigned(2736, 12), 307 => to_unsigned(3775, 12), 308 => to_unsigned(164, 12), 309 => to_unsigned(1621, 12), 310 => to_unsigned(1795, 12), 311 => to_unsigned(265, 12), 312 => to_unsigned(3490, 12), 313 => to_unsigned(50, 12), 314 => to_unsigned(1999, 12), 315 => to_unsigned(933, 12), 316 => to_unsigned(2956, 12), 317 => to_unsigned(1482, 12), 318 => to_unsigned(1556, 12), 319 => to_unsigned(3793, 12), 320 => to_unsigned(3028, 12), 321 => to_unsigned(2454, 12), 322 => to_unsigned(527, 12), 323 => to_unsigned(3043, 12), 324 => to_unsigned(1882, 12), 325 => to_unsigned(2818, 12), 326 => to_unsigned(2835, 12), 327 => to_unsigned(3408, 12), 328 => to_unsigned(2942, 12), 329 => to_unsigned(1587, 12), 330 => to_unsigned(1764, 12), 331 => to_unsigned(3406, 12), 332 => to_unsigned(3174, 12), 333 => to_unsigned(562, 12), 334 => to_unsigned(1751, 12), 335 => to_unsigned(1211, 12), 336 => to_unsigned(939, 12), 337 => to_unsigned(900, 12), 338 => to_unsigned(2866, 12), 339 => to_unsigned(906, 12), 340 => to_unsigned(1132, 12), 341 => to_unsigned(2078, 12), 342 => to_unsigned(800, 12), 343 => to_unsigned(2212, 12), 344 => to_unsigned(1426, 12), 345 => to_unsigned(3607, 12), 346 => to_unsigned(2138, 12), 347 => to_unsigned(3301, 12), 348 => to_unsigned(2735, 12), 349 => to_unsigned(1827, 12), 350 => to_unsigned(1584, 12), 351 => to_unsigned(1663, 12), 352 => to_unsigned(3884, 12), 353 => to_unsigned(61, 12), 354 => to_unsigned(3167, 12), 355 => to_unsigned(2330, 12), 356 => to_unsigned(2021, 12), 357 => to_unsigned(3956, 12), 358 => to_unsigned(2478, 12), 359 => to_unsigned(3617, 12), 360 => to_unsigned(382, 12), 361 => to_unsigned(3640, 12), 362 => to_unsigned(1912, 12), 363 => to_unsigned(2021, 12), 364 => to_unsigned(3271, 12), 365 => to_unsigned(4008, 12), 366 => to_unsigned(1810, 12), 367 => to_unsigned(1257, 12), 368 => to_unsigned(671, 12), 369 => to_unsigned(126, 12), 370 => to_unsigned(3708, 12), 371 => to_unsigned(3903, 12), 372 => to_unsigned(2334, 12), 373 => to_unsigned(3146, 12), 374 => to_unsigned(1949, 12), 375 => to_unsigned(1747, 12), 376 => to_unsigned(2469, 12), 377 => to_unsigned(3985, 12), 378 => to_unsigned(9, 12), 379 => to_unsigned(2446, 12), 380 => to_unsigned(3719, 12), 381 => to_unsigned(2683, 12), 382 => to_unsigned(3726, 12), 383 => to_unsigned(2481, 12), 384 => to_unsigned(3995, 12), 385 => to_unsigned(155, 12), 386 => to_unsigned(2592, 12), 387 => to_unsigned(3506, 12), 388 => to_unsigned(3809, 12), 389 => to_unsigned(480, 12), 390 => to_unsigned(3958, 12), 391 => to_unsigned(487, 12), 392 => to_unsigned(503, 12), 393 => to_unsigned(608, 12), 394 => to_unsigned(855, 12), 395 => to_unsigned(2501, 12), 396 => to_unsigned(81, 12), 397 => to_unsigned(633, 12), 398 => to_unsigned(995, 12), 399 => to_unsigned(996, 12), 400 => to_unsigned(3968, 12), 401 => to_unsigned(2844, 12), 402 => to_unsigned(2476, 12), 403 => to_unsigned(1089, 12), 404 => to_unsigned(2288, 12), 405 => to_unsigned(3760, 12), 406 => to_unsigned(702, 12), 407 => to_unsigned(580, 12), 408 => to_unsigned(125, 12), 409 => to_unsigned(1572, 12), 410 => to_unsigned(3966, 12), 411 => to_unsigned(222, 12), 412 => to_unsigned(2688, 12), 413 => to_unsigned(2613, 12), 414 => to_unsigned(754, 12), 415 => to_unsigned(2346, 12), 416 => to_unsigned(1813, 12), 417 => to_unsigned(2962, 12), 418 => to_unsigned(2859, 12), 419 => to_unsigned(502, 12), 420 => to_unsigned(3681, 12), 421 => to_unsigned(128, 12), 422 => to_unsigned(2174, 12), 423 => to_unsigned(3758, 12), 424 => to_unsigned(2503, 12), 425 => to_unsigned(3628, 12), 426 => to_unsigned(4087, 12), 427 => to_unsigned(590, 12), 428 => to_unsigned(2978, 12), 429 => to_unsigned(2136, 12), 430 => to_unsigned(499, 12), 431 => to_unsigned(318, 12), 432 => to_unsigned(3139, 12), 433 => to_unsigned(2239, 12), 434 => to_unsigned(963, 12), 435 => to_unsigned(1514, 12), 436 => to_unsigned(267, 12), 437 => to_unsigned(2922, 12), 438 => to_unsigned(2088, 12), 439 => to_unsigned(1641, 12), 440 => to_unsigned(291, 12), 441 => to_unsigned(66, 12), 442 => to_unsigned(2788, 12), 443 => to_unsigned(1485, 12), 444 => to_unsigned(1933, 12), 445 => to_unsigned(737, 12), 446 => to_unsigned(2222, 12), 447 => to_unsigned(3906, 12), 448 => to_unsigned(1500, 12), 449 => to_unsigned(3500, 12), 450 => to_unsigned(2064, 12), 451 => to_unsigned(505, 12), 452 => to_unsigned(3873, 12), 453 => to_unsigned(48, 12), 454 => to_unsigned(2744, 12), 455 => to_unsigned(83, 12), 456 => to_unsigned(1078, 12), 457 => to_unsigned(1219, 12), 458 => to_unsigned(2646, 12), 459 => to_unsigned(2900, 12), 460 => to_unsigned(2886, 12), 461 => to_unsigned(3340, 12), 462 => to_unsigned(1331, 12), 463 => to_unsigned(164, 12), 464 => to_unsigned(2009, 12), 465 => to_unsigned(2600, 12), 466 => to_unsigned(70, 12), 467 => to_unsigned(3953, 12), 468 => to_unsigned(3608, 12), 469 => to_unsigned(1463, 12), 470 => to_unsigned(3881, 12), 471 => to_unsigned(3003, 12), 472 => to_unsigned(1013, 12), 473 => to_unsigned(3974, 12), 474 => to_unsigned(2350, 12), 475 => to_unsigned(2424, 12), 476 => to_unsigned(614, 12), 477 => to_unsigned(2625, 12), 478 => to_unsigned(1501, 12), 479 => to_unsigned(4036, 12), 480 => to_unsigned(1305, 12), 481 => to_unsigned(4008, 12), 482 => to_unsigned(795, 12), 483 => to_unsigned(1360, 12), 484 => to_unsigned(3787, 12), 485 => to_unsigned(2513, 12), 486 => to_unsigned(882, 12), 487 => to_unsigned(880, 12), 488 => to_unsigned(3128, 12), 489 => to_unsigned(1486, 12), 490 => to_unsigned(2232, 12), 491 => to_unsigned(2278, 12), 492 => to_unsigned(1553, 12), 493 => to_unsigned(2409, 12), 494 => to_unsigned(751, 12), 495 => to_unsigned(170, 12), 496 => to_unsigned(3616, 12), 497 => to_unsigned(2893, 12), 498 => to_unsigned(3191, 12), 499 => to_unsigned(1032, 12), 500 => to_unsigned(2974, 12), 501 => to_unsigned(2041, 12), 502 => to_unsigned(3152, 12), 503 => to_unsigned(577, 12), 504 => to_unsigned(1715, 12), 505 => to_unsigned(3166, 12), 506 => to_unsigned(2432, 12), 507 => to_unsigned(2630, 12), 508 => to_unsigned(2996, 12), 509 => to_unsigned(3156, 12), 510 => to_unsigned(1963, 12), 511 => to_unsigned(3928, 12), 512 => to_unsigned(1125, 12), 513 => to_unsigned(363, 12), 514 => to_unsigned(3939, 12), 515 => to_unsigned(694, 12), 516 => to_unsigned(402, 12), 517 => to_unsigned(1950, 12), 518 => to_unsigned(390, 12), 519 => to_unsigned(1761, 12), 520 => to_unsigned(1110, 12), 521 => to_unsigned(3903, 12), 522 => to_unsigned(2803, 12), 523 => to_unsigned(3036, 12), 524 => to_unsigned(2264, 12), 525 => to_unsigned(2836, 12), 526 => to_unsigned(669, 12), 527 => to_unsigned(1282, 12), 528 => to_unsigned(1529, 12), 529 => to_unsigned(3670, 12), 530 => to_unsigned(1345, 12), 531 => to_unsigned(2803, 12), 532 => to_unsigned(1860, 12), 533 => to_unsigned(247, 12), 534 => to_unsigned(1911, 12), 535 => to_unsigned(2362, 12), 536 => to_unsigned(2940, 12), 537 => to_unsigned(3245, 12), 538 => to_unsigned(308, 12), 539 => to_unsigned(2487, 12), 540 => to_unsigned(2436, 12), 541 => to_unsigned(3669, 12), 542 => to_unsigned(2682, 12), 543 => to_unsigned(1766, 12), 544 => to_unsigned(1324, 12), 545 => to_unsigned(433, 12), 546 => to_unsigned(817, 12), 547 => to_unsigned(3767, 12), 548 => to_unsigned(1999, 12), 549 => to_unsigned(2175, 12), 550 => to_unsigned(904, 12), 551 => to_unsigned(2204, 12), 552 => to_unsigned(3652, 12), 553 => to_unsigned(673, 12), 554 => to_unsigned(3700, 12), 555 => to_unsigned(1060, 12), 556 => to_unsigned(3698, 12), 557 => to_unsigned(3138, 12), 558 => to_unsigned(750, 12), 559 => to_unsigned(1756, 12), 560 => to_unsigned(3121, 12), 561 => to_unsigned(559, 12), 562 => to_unsigned(1215, 12), 563 => to_unsigned(832, 12), 564 => to_unsigned(2462, 12), 565 => to_unsigned(2931, 12), 566 => to_unsigned(1925, 12), 567 => to_unsigned(2321, 12), 568 => to_unsigned(3221, 12), 569 => to_unsigned(1120, 12), 570 => to_unsigned(229, 12), 571 => to_unsigned(2627, 12), 572 => to_unsigned(2864, 12), 573 => to_unsigned(635, 12), 574 => to_unsigned(1990, 12), 575 => to_unsigned(1561, 12), 576 => to_unsigned(3886, 12), 577 => to_unsigned(1147, 12), 578 => to_unsigned(1012, 12), 579 => to_unsigned(1582, 12), 580 => to_unsigned(2949, 12), 581 => to_unsigned(1636, 12), 582 => to_unsigned(1063, 12), 583 => to_unsigned(1269, 12), 584 => to_unsigned(320, 12), 585 => to_unsigned(3101, 12), 586 => to_unsigned(1080, 12), 587 => to_unsigned(2257, 12), 588 => to_unsigned(1482, 12), 589 => to_unsigned(3967, 12), 590 => to_unsigned(893, 12), 591 => to_unsigned(3217, 12), 592 => to_unsigned(1666, 12), 593 => to_unsigned(1050, 12), 594 => to_unsigned(2355, 12), 595 => to_unsigned(428, 12), 596 => to_unsigned(3945, 12), 597 => to_unsigned(3268, 12), 598 => to_unsigned(344, 12), 599 => to_unsigned(3789, 12), 600 => to_unsigned(1386, 12), 601 => to_unsigned(1795, 12), 602 => to_unsigned(738, 12), 603 => to_unsigned(1668, 12), 604 => to_unsigned(1454, 12), 605 => to_unsigned(3787, 12), 606 => to_unsigned(2106, 12), 607 => to_unsigned(726, 12), 608 => to_unsigned(2696, 12), 609 => to_unsigned(3542, 12), 610 => to_unsigned(398, 12), 611 => to_unsigned(1772, 12), 612 => to_unsigned(3213, 12), 613 => to_unsigned(3721, 12), 614 => to_unsigned(849, 12), 615 => to_unsigned(3378, 12), 616 => to_unsigned(8, 12), 617 => to_unsigned(2672, 12), 618 => to_unsigned(3161, 12), 619 => to_unsigned(329, 12), 620 => to_unsigned(3566, 12), 621 => to_unsigned(2464, 12), 622 => to_unsigned(2209, 12), 623 => to_unsigned(3931, 12), 624 => to_unsigned(421, 12), 625 => to_unsigned(807, 12), 626 => to_unsigned(658, 12), 627 => to_unsigned(2948, 12), 628 => to_unsigned(3765, 12), 629 => to_unsigned(3718, 12), 630 => to_unsigned(1039, 12), 631 => to_unsigned(944, 12), 632 => to_unsigned(1162, 12), 633 => to_unsigned(3700, 12), 634 => to_unsigned(2106, 12), 635 => to_unsigned(3204, 12), 636 => to_unsigned(1607, 12), 637 => to_unsigned(51, 12), 638 => to_unsigned(3297, 12), 639 => to_unsigned(3481, 12), 640 => to_unsigned(1725, 12), 641 => to_unsigned(1703, 12), 642 => to_unsigned(3374, 12), 643 => to_unsigned(1142, 12), 644 => to_unsigned(1014, 12), 645 => to_unsigned(133, 12), 646 => to_unsigned(2022, 12), 647 => to_unsigned(1608, 12), 648 => to_unsigned(3732, 12), 649 => to_unsigned(67, 12), 650 => to_unsigned(116, 12), 651 => to_unsigned(3169, 12), 652 => to_unsigned(4016, 12), 653 => to_unsigned(409, 12), 654 => to_unsigned(3419, 12), 655 => to_unsigned(2446, 12), 656 => to_unsigned(3226, 12), 657 => to_unsigned(612, 12), 658 => to_unsigned(3324, 12), 659 => to_unsigned(824, 12), 660 => to_unsigned(2664, 12), 661 => to_unsigned(3203, 12), 662 => to_unsigned(3054, 12), 663 => to_unsigned(3887, 12), 664 => to_unsigned(297, 12), 665 => to_unsigned(3748, 12), 666 => to_unsigned(2575, 12), 667 => to_unsigned(3336, 12), 668 => to_unsigned(1631, 12), 669 => to_unsigned(2218, 12), 670 => to_unsigned(2230, 12), 671 => to_unsigned(27, 12), 672 => to_unsigned(3024, 12), 673 => to_unsigned(559, 12), 674 => to_unsigned(3247, 12), 675 => to_unsigned(2555, 12), 676 => to_unsigned(1872, 12), 677 => to_unsigned(1946, 12), 678 => to_unsigned(3154, 12), 679 => to_unsigned(1494, 12), 680 => to_unsigned(0, 12), 681 => to_unsigned(3513, 12), 682 => to_unsigned(3038, 12), 683 => to_unsigned(2500, 12), 684 => to_unsigned(84, 12), 685 => to_unsigned(3039, 12), 686 => to_unsigned(2603, 12), 687 => to_unsigned(3644, 12), 688 => to_unsigned(2859, 12), 689 => to_unsigned(202, 12), 690 => to_unsigned(1825, 12), 691 => to_unsigned(1198, 12), 692 => to_unsigned(1171, 12), 693 => to_unsigned(684, 12), 694 => to_unsigned(1537, 12), 695 => to_unsigned(3595, 12), 696 => to_unsigned(2357, 12), 697 => to_unsigned(337, 12), 698 => to_unsigned(3847, 12), 699 => to_unsigned(3193, 12), 700 => to_unsigned(1908, 12), 701 => to_unsigned(5, 12), 702 => to_unsigned(1634, 12), 703 => to_unsigned(3213, 12), 704 => to_unsigned(117, 12), 705 => to_unsigned(1752, 12), 706 => to_unsigned(2233, 12), 707 => to_unsigned(1376, 12), 708 => to_unsigned(3198, 12), 709 => to_unsigned(3209, 12), 710 => to_unsigned(3276, 12), 711 => to_unsigned(3252, 12), 712 => to_unsigned(843, 12), 713 => to_unsigned(3197, 12), 714 => to_unsigned(2057, 12), 715 => to_unsigned(2808, 12), 716 => to_unsigned(3991, 12), 717 => to_unsigned(2902, 12), 718 => to_unsigned(3346, 12), 719 => to_unsigned(3970, 12), 720 => to_unsigned(133, 12), 721 => to_unsigned(2801, 12), 722 => to_unsigned(144, 12), 723 => to_unsigned(3345, 12), 724 => to_unsigned(3983, 12), 725 => to_unsigned(146, 12), 726 => to_unsigned(3123, 12), 727 => to_unsigned(1383, 12), 728 => to_unsigned(1386, 12), 729 => to_unsigned(3154, 12), 730 => to_unsigned(118, 12), 731 => to_unsigned(3338, 12), 732 => to_unsigned(1132, 12), 733 => to_unsigned(3933, 12), 734 => to_unsigned(2663, 12), 735 => to_unsigned(859, 12), 736 => to_unsigned(1171, 12), 737 => to_unsigned(721, 12), 738 => to_unsigned(3720, 12), 739 => to_unsigned(1327, 12), 740 => to_unsigned(1921, 12), 741 => to_unsigned(89, 12), 742 => to_unsigned(1569, 12), 743 => to_unsigned(26, 12), 744 => to_unsigned(2373, 12), 745 => to_unsigned(1789, 12), 746 => to_unsigned(2824, 12), 747 => to_unsigned(3735, 12), 748 => to_unsigned(873, 12), 749 => to_unsigned(3159, 12), 750 => to_unsigned(631, 12), 751 => to_unsigned(2533, 12), 752 => to_unsigned(2320, 12), 753 => to_unsigned(2647, 12), 754 => to_unsigned(3266, 12), 755 => to_unsigned(2755, 12), 756 => to_unsigned(2687, 12), 757 => to_unsigned(3167, 12), 758 => to_unsigned(2058, 12), 759 => to_unsigned(681, 12), 760 => to_unsigned(831, 12), 761 => to_unsigned(1141, 12), 762 => to_unsigned(790, 12), 763 => to_unsigned(1122, 12), 764 => to_unsigned(2871, 12), 765 => to_unsigned(2559, 12), 766 => to_unsigned(3653, 12), 767 => to_unsigned(1586, 12), 768 => to_unsigned(101, 12), 769 => to_unsigned(210, 12), 770 => to_unsigned(3444, 12), 771 => to_unsigned(1618, 12), 772 => to_unsigned(2070, 12), 773 => to_unsigned(2368, 12), 774 => to_unsigned(3795, 12), 775 => to_unsigned(1751, 12), 776 => to_unsigned(2642, 12), 777 => to_unsigned(3994, 12), 778 => to_unsigned(1294, 12), 779 => to_unsigned(888, 12), 780 => to_unsigned(2568, 12), 781 => to_unsigned(3170, 12), 782 => to_unsigned(941, 12), 783 => to_unsigned(929, 12), 784 => to_unsigned(1323, 12), 785 => to_unsigned(2128, 12), 786 => to_unsigned(4025, 12), 787 => to_unsigned(2057, 12), 788 => to_unsigned(257, 12), 789 => to_unsigned(3695, 12), 790 => to_unsigned(2144, 12), 791 => to_unsigned(3372, 12), 792 => to_unsigned(2792, 12), 793 => to_unsigned(981, 12), 794 => to_unsigned(1737, 12), 795 => to_unsigned(2038, 12), 796 => to_unsigned(1600, 12), 797 => to_unsigned(705, 12), 798 => to_unsigned(1152, 12), 799 => to_unsigned(272, 12), 800 => to_unsigned(1066, 12), 801 => to_unsigned(3445, 12), 802 => to_unsigned(222, 12), 803 => to_unsigned(862, 12), 804 => to_unsigned(304, 12), 805 => to_unsigned(3374, 12), 806 => to_unsigned(2024, 12), 807 => to_unsigned(1084, 12), 808 => to_unsigned(2994, 12), 809 => to_unsigned(1160, 12), 810 => to_unsigned(2728, 12), 811 => to_unsigned(2502, 12), 812 => to_unsigned(2363, 12), 813 => to_unsigned(1237, 12), 814 => to_unsigned(2314, 12), 815 => to_unsigned(2359, 12), 816 => to_unsigned(388, 12), 817 => to_unsigned(2963, 12), 818 => to_unsigned(3206, 12), 819 => to_unsigned(113, 12), 820 => to_unsigned(3948, 12), 821 => to_unsigned(3397, 12), 822 => to_unsigned(1377, 12), 823 => to_unsigned(3818, 12), 824 => to_unsigned(1069, 12), 825 => to_unsigned(2052, 12), 826 => to_unsigned(745, 12), 827 => to_unsigned(1539, 12), 828 => to_unsigned(3145, 12), 829 => to_unsigned(2946, 12), 830 => to_unsigned(361, 12), 831 => to_unsigned(651, 12), 832 => to_unsigned(4044, 12), 833 => to_unsigned(3526, 12), 834 => to_unsigned(2802, 12), 835 => to_unsigned(2162, 12), 836 => to_unsigned(3972, 12), 837 => to_unsigned(3368, 12), 838 => to_unsigned(1549, 12), 839 => to_unsigned(2873, 12), 840 => to_unsigned(3146, 12), 841 => to_unsigned(458, 12), 842 => to_unsigned(3530, 12), 843 => to_unsigned(1548, 12), 844 => to_unsigned(2373, 12), 845 => to_unsigned(2512, 12), 846 => to_unsigned(2603, 12), 847 => to_unsigned(1619, 12), 848 => to_unsigned(3602, 12), 849 => to_unsigned(3398, 12), 850 => to_unsigned(1403, 12), 851 => to_unsigned(2138, 12), 852 => to_unsigned(4078, 12), 853 => to_unsigned(1542, 12), 854 => to_unsigned(2, 12), 855 => to_unsigned(541, 12), 856 => to_unsigned(3522, 12), 857 => to_unsigned(1205, 12), 858 => to_unsigned(3458, 12), 859 => to_unsigned(3346, 12), 860 => to_unsigned(1943, 12), 861 => to_unsigned(1287, 12), 862 => to_unsigned(2707, 12), 863 => to_unsigned(3429, 12), 864 => to_unsigned(988, 12), 865 => to_unsigned(1009, 12), 866 => to_unsigned(2757, 12), 867 => to_unsigned(2292, 12), 868 => to_unsigned(635, 12), 869 => to_unsigned(2245, 12), 870 => to_unsigned(50, 12), 871 => to_unsigned(1337, 12), 872 => to_unsigned(3555, 12), 873 => to_unsigned(3436, 12), 874 => to_unsigned(287, 12), 875 => to_unsigned(2691, 12), 876 => to_unsigned(785, 12), 877 => to_unsigned(3758, 12), 878 => to_unsigned(1737, 12), 879 => to_unsigned(905, 12), 880 => to_unsigned(837, 12), 881 => to_unsigned(3234, 12), 882 => to_unsigned(3069, 12), 883 => to_unsigned(615, 12), 884 => to_unsigned(1824, 12), 885 => to_unsigned(3935, 12), 886 => to_unsigned(873, 12), 887 => to_unsigned(736, 12), 888 => to_unsigned(153, 12), 889 => to_unsigned(3539, 12), 890 => to_unsigned(3231, 12), 891 => to_unsigned(1715, 12), 892 => to_unsigned(3719, 12), 893 => to_unsigned(3380, 12), 894 => to_unsigned(2006, 12), 895 => to_unsigned(1679, 12), 896 => to_unsigned(3250, 12), 897 => to_unsigned(2992, 12), 898 => to_unsigned(548, 12), 899 => to_unsigned(2906, 12), 900 => to_unsigned(294, 12), 901 => to_unsigned(1254, 12), 902 => to_unsigned(738, 12), 903 => to_unsigned(1176, 12), 904 => to_unsigned(2665, 12), 905 => to_unsigned(2654, 12), 906 => to_unsigned(1793, 12), 907 => to_unsigned(3113, 12), 908 => to_unsigned(3831, 12), 909 => to_unsigned(1528, 12), 910 => to_unsigned(3288, 12), 911 => to_unsigned(1371, 12), 912 => to_unsigned(2219, 12), 913 => to_unsigned(3728, 12), 914 => to_unsigned(972, 12), 915 => to_unsigned(1097, 12), 916 => to_unsigned(193, 12), 917 => to_unsigned(843, 12), 918 => to_unsigned(1710, 12), 919 => to_unsigned(122, 12), 920 => to_unsigned(904, 12), 921 => to_unsigned(530, 12), 922 => to_unsigned(3856, 12), 923 => to_unsigned(3624, 12), 924 => to_unsigned(874, 12), 925 => to_unsigned(242, 12), 926 => to_unsigned(2905, 12), 927 => to_unsigned(3208, 12), 928 => to_unsigned(1646, 12), 929 => to_unsigned(2806, 12), 930 => to_unsigned(1242, 12), 931 => to_unsigned(1922, 12), 932 => to_unsigned(3352, 12), 933 => to_unsigned(318, 12), 934 => to_unsigned(587, 12), 935 => to_unsigned(1256, 12), 936 => to_unsigned(2758, 12), 937 => to_unsigned(3389, 12), 938 => to_unsigned(1773, 12), 939 => to_unsigned(514, 12), 940 => to_unsigned(2257, 12), 941 => to_unsigned(512, 12), 942 => to_unsigned(661, 12), 943 => to_unsigned(2464, 12), 944 => to_unsigned(954, 12), 945 => to_unsigned(3308, 12), 946 => to_unsigned(3612, 12), 947 => to_unsigned(332, 12), 948 => to_unsigned(1211, 12), 949 => to_unsigned(637, 12), 950 => to_unsigned(3228, 12), 951 => to_unsigned(1253, 12), 952 => to_unsigned(3195, 12), 953 => to_unsigned(1534, 12), 954 => to_unsigned(4055, 12), 955 => to_unsigned(2866, 12), 956 => to_unsigned(3161, 12), 957 => to_unsigned(3510, 12), 958 => to_unsigned(747, 12), 959 => to_unsigned(1679, 12), 960 => to_unsigned(1228, 12), 961 => to_unsigned(3949, 12), 962 => to_unsigned(2664, 12), 963 => to_unsigned(3791, 12), 964 => to_unsigned(1626, 12), 965 => to_unsigned(2471, 12), 966 => to_unsigned(132, 12), 967 => to_unsigned(3250, 12), 968 => to_unsigned(3969, 12), 969 => to_unsigned(3567, 12), 970 => to_unsigned(3999, 12), 971 => to_unsigned(2557, 12), 972 => to_unsigned(2160, 12), 973 => to_unsigned(753, 12), 974 => to_unsigned(3513, 12), 975 => to_unsigned(2687, 12), 976 => to_unsigned(1924, 12), 977 => to_unsigned(3694, 12), 978 => to_unsigned(1237, 12), 979 => to_unsigned(2125, 12), 980 => to_unsigned(1563, 12), 981 => to_unsigned(1348, 12), 982 => to_unsigned(324, 12), 983 => to_unsigned(4012, 12), 984 => to_unsigned(1149, 12), 985 => to_unsigned(2822, 12), 986 => to_unsigned(2463, 12), 987 => to_unsigned(634, 12), 988 => to_unsigned(250, 12), 989 => to_unsigned(2552, 12), 990 => to_unsigned(3332, 12), 991 => to_unsigned(3631, 12), 992 => to_unsigned(1480, 12), 993 => to_unsigned(3616, 12), 994 => to_unsigned(233, 12), 995 => to_unsigned(2797, 12), 996 => to_unsigned(2568, 12), 997 => to_unsigned(884, 12), 998 => to_unsigned(3610, 12), 999 => to_unsigned(4030, 12), 1000 => to_unsigned(2444, 12), 1001 => to_unsigned(3532, 12), 1002 => to_unsigned(3511, 12), 1003 => to_unsigned(1829, 12), 1004 => to_unsigned(970, 12), 1005 => to_unsigned(2311, 12), 1006 => to_unsigned(1875, 12), 1007 => to_unsigned(2071, 12), 1008 => to_unsigned(1280, 12), 1009 => to_unsigned(2028, 12), 1010 => to_unsigned(2289, 12), 1011 => to_unsigned(466, 12), 1012 => to_unsigned(1636, 12), 1013 => to_unsigned(3938, 12), 1014 => to_unsigned(3573, 12), 1015 => to_unsigned(385, 12), 1016 => to_unsigned(3455, 12), 1017 => to_unsigned(3288, 12), 1018 => to_unsigned(4084, 12), 1019 => to_unsigned(2728, 12), 1020 => to_unsigned(620, 12), 1021 => to_unsigned(1895, 12), 1022 => to_unsigned(2455, 12), 1023 => to_unsigned(419, 12), 1024 => to_unsigned(800, 12), 1025 => to_unsigned(2750, 12), 1026 => to_unsigned(3796, 12), 1027 => to_unsigned(1064, 12), 1028 => to_unsigned(3933, 12), 1029 => to_unsigned(2392, 12), 1030 => to_unsigned(2605, 12), 1031 => to_unsigned(197, 12), 1032 => to_unsigned(2327, 12), 1033 => to_unsigned(2896, 12), 1034 => to_unsigned(2410, 12), 1035 => to_unsigned(963, 12), 1036 => to_unsigned(2040, 12), 1037 => to_unsigned(758, 12), 1038 => to_unsigned(653, 12), 1039 => to_unsigned(3840, 12), 1040 => to_unsigned(4079, 12), 1041 => to_unsigned(801, 12), 1042 => to_unsigned(1723, 12), 1043 => to_unsigned(1330, 12), 1044 => to_unsigned(2061, 12), 1045 => to_unsigned(1736, 12), 1046 => to_unsigned(146, 12), 1047 => to_unsigned(1453, 12), 1048 => to_unsigned(2756, 12), 1049 => to_unsigned(1010, 12), 1050 => to_unsigned(1312, 12), 1051 => to_unsigned(2680, 12), 1052 => to_unsigned(733, 12), 1053 => to_unsigned(973, 12), 1054 => to_unsigned(3896, 12), 1055 => to_unsigned(1741, 12), 1056 => to_unsigned(1016, 12), 1057 => to_unsigned(2437, 12), 1058 => to_unsigned(1219, 12), 1059 => to_unsigned(3928, 12), 1060 => to_unsigned(953, 12), 1061 => to_unsigned(1630, 12), 1062 => to_unsigned(2501, 12), 1063 => to_unsigned(4047, 12), 1064 => to_unsigned(2197, 12), 1065 => to_unsigned(2552, 12), 1066 => to_unsigned(1563, 12), 1067 => to_unsigned(1741, 12), 1068 => to_unsigned(27, 12), 1069 => to_unsigned(877, 12), 1070 => to_unsigned(1655, 12), 1071 => to_unsigned(2652, 12), 1072 => to_unsigned(3916, 12), 1073 => to_unsigned(2095, 12), 1074 => to_unsigned(2725, 12), 1075 => to_unsigned(772, 12), 1076 => to_unsigned(3267, 12), 1077 => to_unsigned(3051, 12), 1078 => to_unsigned(1882, 12), 1079 => to_unsigned(399, 12), 1080 => to_unsigned(926, 12), 1081 => to_unsigned(2997, 12), 1082 => to_unsigned(45, 12), 1083 => to_unsigned(1079, 12), 1084 => to_unsigned(642, 12), 1085 => to_unsigned(2286, 12), 1086 => to_unsigned(2166, 12), 1087 => to_unsigned(2712, 12), 1088 => to_unsigned(1874, 12), 1089 => to_unsigned(152, 12), 1090 => to_unsigned(2452, 12), 1091 => to_unsigned(218, 12), 1092 => to_unsigned(3807, 12), 1093 => to_unsigned(1099, 12), 1094 => to_unsigned(2793, 12), 1095 => to_unsigned(3974, 12), 1096 => to_unsigned(3060, 12), 1097 => to_unsigned(3274, 12), 1098 => to_unsigned(2104, 12), 1099 => to_unsigned(2940, 12), 1100 => to_unsigned(688, 12), 1101 => to_unsigned(47, 12), 1102 => to_unsigned(70, 12), 1103 => to_unsigned(3509, 12), 1104 => to_unsigned(3239, 12), 1105 => to_unsigned(3678, 12), 1106 => to_unsigned(2534, 12), 1107 => to_unsigned(1620, 12), 1108 => to_unsigned(3632, 12), 1109 => to_unsigned(3717, 12), 1110 => to_unsigned(33, 12), 1111 => to_unsigned(3866, 12), 1112 => to_unsigned(2780, 12), 1113 => to_unsigned(691, 12), 1114 => to_unsigned(3705, 12), 1115 => to_unsigned(3278, 12), 1116 => to_unsigned(121, 12), 1117 => to_unsigned(912, 12), 1118 => to_unsigned(3693, 12), 1119 => to_unsigned(3283, 12), 1120 => to_unsigned(2379, 12), 1121 => to_unsigned(2573, 12), 1122 => to_unsigned(57, 12), 1123 => to_unsigned(3509, 12), 1124 => to_unsigned(1829, 12), 1125 => to_unsigned(285, 12), 1126 => to_unsigned(1771, 12), 1127 => to_unsigned(3240, 12), 1128 => to_unsigned(2719, 12), 1129 => to_unsigned(475, 12), 1130 => to_unsigned(347, 12), 1131 => to_unsigned(3842, 12), 1132 => to_unsigned(2261, 12), 1133 => to_unsigned(3838, 12), 1134 => to_unsigned(447, 12), 1135 => to_unsigned(4054, 12), 1136 => to_unsigned(510, 12), 1137 => to_unsigned(733, 12), 1138 => to_unsigned(364, 12), 1139 => to_unsigned(38, 12), 1140 => to_unsigned(2478, 12), 1141 => to_unsigned(3992, 12), 1142 => to_unsigned(3404, 12), 1143 => to_unsigned(3677, 12), 1144 => to_unsigned(401, 12), 1145 => to_unsigned(460, 12), 1146 => to_unsigned(1220, 12), 1147 => to_unsigned(1801, 12), 1148 => to_unsigned(1938, 12), 1149 => to_unsigned(1830, 12), 1150 => to_unsigned(4057, 12), 1151 => to_unsigned(1615, 12), 1152 => to_unsigned(3672, 12), 1153 => to_unsigned(3063, 12), 1154 => to_unsigned(2771, 12), 1155 => to_unsigned(3735, 12), 1156 => to_unsigned(3945, 12), 1157 => to_unsigned(2876, 12), 1158 => to_unsigned(3124, 12), 1159 => to_unsigned(274, 12), 1160 => to_unsigned(2886, 12), 1161 => to_unsigned(3400, 12), 1162 => to_unsigned(3722, 12), 1163 => to_unsigned(3864, 12), 1164 => to_unsigned(1773, 12), 1165 => to_unsigned(1708, 12), 1166 => to_unsigned(3563, 12), 1167 => to_unsigned(1793, 12), 1168 => to_unsigned(723, 12), 1169 => to_unsigned(114, 12), 1170 => to_unsigned(3250, 12), 1171 => to_unsigned(2342, 12), 1172 => to_unsigned(1179, 12), 1173 => to_unsigned(3731, 12), 1174 => to_unsigned(323, 12), 1175 => to_unsigned(3450, 12), 1176 => to_unsigned(3144, 12), 1177 => to_unsigned(598, 12), 1178 => to_unsigned(3258, 12), 1179 => to_unsigned(574, 12), 1180 => to_unsigned(2572, 12), 1181 => to_unsigned(704, 12), 1182 => to_unsigned(1808, 12), 1183 => to_unsigned(3864, 12), 1184 => to_unsigned(3442, 12), 1185 => to_unsigned(3423, 12), 1186 => to_unsigned(2528, 12), 1187 => to_unsigned(1123, 12), 1188 => to_unsigned(1605, 12), 1189 => to_unsigned(885, 12), 1190 => to_unsigned(3126, 12), 1191 => to_unsigned(3194, 12), 1192 => to_unsigned(3269, 12), 1193 => to_unsigned(317, 12), 1194 => to_unsigned(2689, 12), 1195 => to_unsigned(2584, 12), 1196 => to_unsigned(1804, 12), 1197 => to_unsigned(1969, 12), 1198 => to_unsigned(4009, 12), 1199 => to_unsigned(1718, 12), 1200 => to_unsigned(3411, 12), 1201 => to_unsigned(1206, 12), 1202 => to_unsigned(3487, 12), 1203 => to_unsigned(490, 12), 1204 => to_unsigned(967, 12), 1205 => to_unsigned(2836, 12), 1206 => to_unsigned(538, 12), 1207 => to_unsigned(541, 12), 1208 => to_unsigned(307, 12), 1209 => to_unsigned(3533, 12), 1210 => to_unsigned(2131, 12), 1211 => to_unsigned(2002, 12), 1212 => to_unsigned(2112, 12), 1213 => to_unsigned(1001, 12), 1214 => to_unsigned(609, 12), 1215 => to_unsigned(2980, 12), 1216 => to_unsigned(2266, 12), 1217 => to_unsigned(1277, 12), 1218 => to_unsigned(3610, 12), 1219 => to_unsigned(2302, 12), 1220 => to_unsigned(1509, 12), 1221 => to_unsigned(1163, 12), 1222 => to_unsigned(2171, 12), 1223 => to_unsigned(3208, 12), 1224 => to_unsigned(3194, 12), 1225 => to_unsigned(602, 12), 1226 => to_unsigned(1053, 12), 1227 => to_unsigned(1261, 12), 1228 => to_unsigned(191, 12), 1229 => to_unsigned(1724, 12), 1230 => to_unsigned(791, 12), 1231 => to_unsigned(4050, 12), 1232 => to_unsigned(3952, 12), 1233 => to_unsigned(150, 12), 1234 => to_unsigned(867, 12), 1235 => to_unsigned(1127, 12), 1236 => to_unsigned(3243, 12), 1237 => to_unsigned(1425, 12), 1238 => to_unsigned(3134, 12), 1239 => to_unsigned(1368, 12), 1240 => to_unsigned(3732, 12), 1241 => to_unsigned(3990, 12), 1242 => to_unsigned(3657, 12), 1243 => to_unsigned(2858, 12), 1244 => to_unsigned(1877, 12), 1245 => to_unsigned(3197, 12), 1246 => to_unsigned(1597, 12), 1247 => to_unsigned(1101, 12), 1248 => to_unsigned(1967, 12), 1249 => to_unsigned(2029, 12), 1250 => to_unsigned(625, 12), 1251 => to_unsigned(2174, 12), 1252 => to_unsigned(901, 12), 1253 => to_unsigned(3741, 12), 1254 => to_unsigned(683, 12), 1255 => to_unsigned(2113, 12), 1256 => to_unsigned(3547, 12), 1257 => to_unsigned(3395, 12), 1258 => to_unsigned(2841, 12), 1259 => to_unsigned(144, 12), 1260 => to_unsigned(2640, 12), 1261 => to_unsigned(2284, 12), 1262 => to_unsigned(1711, 12), 1263 => to_unsigned(2494, 12), 1264 => to_unsigned(11, 12), 1265 => to_unsigned(2632, 12), 1266 => to_unsigned(2078, 12), 1267 => to_unsigned(495, 12), 1268 => to_unsigned(1198, 12), 1269 => to_unsigned(2836, 12), 1270 => to_unsigned(3659, 12), 1271 => to_unsigned(3868, 12), 1272 => to_unsigned(3346, 12), 1273 => to_unsigned(2756, 12), 1274 => to_unsigned(2118, 12), 1275 => to_unsigned(1301, 12), 1276 => to_unsigned(363, 12), 1277 => to_unsigned(3960, 12), 1278 => to_unsigned(3205, 12), 1279 => to_unsigned(1, 12), 1280 => to_unsigned(3934, 12), 1281 => to_unsigned(3915, 12), 1282 => to_unsigned(1117, 12), 1283 => to_unsigned(1899, 12), 1284 => to_unsigned(1280, 12), 1285 => to_unsigned(1772, 12), 1286 => to_unsigned(1426, 12), 1287 => to_unsigned(2497, 12), 1288 => to_unsigned(212, 12), 1289 => to_unsigned(1209, 12), 1290 => to_unsigned(499, 12), 1291 => to_unsigned(2143, 12), 1292 => to_unsigned(2163, 12), 1293 => to_unsigned(550, 12), 1294 => to_unsigned(3163, 12), 1295 => to_unsigned(2285, 12), 1296 => to_unsigned(2318, 12), 1297 => to_unsigned(1949, 12), 1298 => to_unsigned(3196, 12), 1299 => to_unsigned(734, 12), 1300 => to_unsigned(257, 12), 1301 => to_unsigned(2619, 12), 1302 => to_unsigned(134, 12), 1303 => to_unsigned(2381, 12), 1304 => to_unsigned(1061, 12), 1305 => to_unsigned(1570, 12), 1306 => to_unsigned(3866, 12), 1307 => to_unsigned(2228, 12), 1308 => to_unsigned(1283, 12), 1309 => to_unsigned(417, 12), 1310 => to_unsigned(2773, 12), 1311 => to_unsigned(3816, 12), 1312 => to_unsigned(4030, 12), 1313 => to_unsigned(1910, 12), 1314 => to_unsigned(1688, 12), 1315 => to_unsigned(3112, 12), 1316 => to_unsigned(1918, 12), 1317 => to_unsigned(1607, 12), 1318 => to_unsigned(2215, 12), 1319 => to_unsigned(2665, 12), 1320 => to_unsigned(249, 12), 1321 => to_unsigned(66, 12), 1322 => to_unsigned(682, 12), 1323 => to_unsigned(775, 12), 1324 => to_unsigned(3040, 12), 1325 => to_unsigned(191, 12), 1326 => to_unsigned(1993, 12), 1327 => to_unsigned(3483, 12), 1328 => to_unsigned(908, 12), 1329 => to_unsigned(2045, 12), 1330 => to_unsigned(2945, 12), 1331 => to_unsigned(145, 12), 1332 => to_unsigned(3741, 12), 1333 => to_unsigned(1746, 12), 1334 => to_unsigned(641, 12), 1335 => to_unsigned(1850, 12), 1336 => to_unsigned(3172, 12), 1337 => to_unsigned(1095, 12), 1338 => to_unsigned(3830, 12), 1339 => to_unsigned(447, 12), 1340 => to_unsigned(1494, 12), 1341 => to_unsigned(2935, 12), 1342 => to_unsigned(955, 12), 1343 => to_unsigned(3070, 12), 1344 => to_unsigned(235, 12), 1345 => to_unsigned(2581, 12), 1346 => to_unsigned(3884, 12), 1347 => to_unsigned(2643, 12), 1348 => to_unsigned(3044, 12), 1349 => to_unsigned(2340, 12), 1350 => to_unsigned(1206, 12), 1351 => to_unsigned(1182, 12), 1352 => to_unsigned(2146, 12), 1353 => to_unsigned(895, 12), 1354 => to_unsigned(4081, 12), 1355 => to_unsigned(3644, 12), 1356 => to_unsigned(3195, 12), 1357 => to_unsigned(1066, 12), 1358 => to_unsigned(3678, 12), 1359 => to_unsigned(3122, 12), 1360 => to_unsigned(1213, 12), 1361 => to_unsigned(328, 12), 1362 => to_unsigned(3675, 12), 1363 => to_unsigned(3819, 12), 1364 => to_unsigned(1988, 12), 1365 => to_unsigned(1191, 12), 1366 => to_unsigned(3891, 12), 1367 => to_unsigned(3370, 12), 1368 => to_unsigned(1650, 12), 1369 => to_unsigned(3917, 12), 1370 => to_unsigned(2084, 12), 1371 => to_unsigned(2538, 12), 1372 => to_unsigned(301, 12), 1373 => to_unsigned(747, 12), 1374 => to_unsigned(712, 12), 1375 => to_unsigned(1803, 12), 1376 => to_unsigned(785, 12), 1377 => to_unsigned(1999, 12), 1378 => to_unsigned(3346, 12), 1379 => to_unsigned(1472, 12), 1380 => to_unsigned(4087, 12), 1381 => to_unsigned(182, 12), 1382 => to_unsigned(1204, 12), 1383 => to_unsigned(2257, 12), 1384 => to_unsigned(105, 12), 1385 => to_unsigned(2986, 12), 1386 => to_unsigned(3927, 12), 1387 => to_unsigned(2974, 12), 1388 => to_unsigned(2585, 12), 1389 => to_unsigned(3901, 12), 1390 => to_unsigned(1541, 12), 1391 => to_unsigned(2447, 12), 1392 => to_unsigned(873, 12), 1393 => to_unsigned(1429, 12), 1394 => to_unsigned(912, 12), 1395 => to_unsigned(786, 12), 1396 => to_unsigned(3849, 12), 1397 => to_unsigned(1571, 12), 1398 => to_unsigned(1065, 12), 1399 => to_unsigned(1874, 12), 1400 => to_unsigned(579, 12), 1401 => to_unsigned(2626, 12), 1402 => to_unsigned(2191, 12), 1403 => to_unsigned(3728, 12), 1404 => to_unsigned(1162, 12), 1405 => to_unsigned(2025, 12), 1406 => to_unsigned(1828, 12), 1407 => to_unsigned(2160, 12), 1408 => to_unsigned(3267, 12), 1409 => to_unsigned(2771, 12), 1410 => to_unsigned(2021, 12), 1411 => to_unsigned(1817, 12), 1412 => to_unsigned(3632, 12), 1413 => to_unsigned(1690, 12), 1414 => to_unsigned(3977, 12), 1415 => to_unsigned(1494, 12), 1416 => to_unsigned(1818, 12), 1417 => to_unsigned(2169, 12), 1418 => to_unsigned(3072, 12), 1419 => to_unsigned(961, 12), 1420 => to_unsigned(3537, 12), 1421 => to_unsigned(2420, 12), 1422 => to_unsigned(3153, 12), 1423 => to_unsigned(1135, 12), 1424 => to_unsigned(495, 12), 1425 => to_unsigned(2998, 12), 1426 => to_unsigned(624, 12), 1427 => to_unsigned(447, 12), 1428 => to_unsigned(446, 12), 1429 => to_unsigned(2102, 12), 1430 => to_unsigned(7, 12), 1431 => to_unsigned(1179, 12), 1432 => to_unsigned(1274, 12), 1433 => to_unsigned(2536, 12), 1434 => to_unsigned(286, 12), 1435 => to_unsigned(2147, 12), 1436 => to_unsigned(2466, 12), 1437 => to_unsigned(3630, 12), 1438 => to_unsigned(803, 12), 1439 => to_unsigned(2129, 12), 1440 => to_unsigned(2519, 12), 1441 => to_unsigned(1006, 12), 1442 => to_unsigned(820, 12), 1443 => to_unsigned(2270, 12), 1444 => to_unsigned(2836, 12), 1445 => to_unsigned(4094, 12), 1446 => to_unsigned(82, 12), 1447 => to_unsigned(964, 12), 1448 => to_unsigned(1652, 12), 1449 => to_unsigned(292, 12), 1450 => to_unsigned(1925, 12), 1451 => to_unsigned(2628, 12), 1452 => to_unsigned(2368, 12), 1453 => to_unsigned(1905, 12), 1454 => to_unsigned(315, 12), 1455 => to_unsigned(799, 12), 1456 => to_unsigned(3128, 12), 1457 => to_unsigned(3667, 12), 1458 => to_unsigned(1872, 12), 1459 => to_unsigned(2664, 12), 1460 => to_unsigned(784, 12), 1461 => to_unsigned(3981, 12), 1462 => to_unsigned(1447, 12), 1463 => to_unsigned(1396, 12), 1464 => to_unsigned(495, 12), 1465 => to_unsigned(1275, 12), 1466 => to_unsigned(1795, 12), 1467 => to_unsigned(2532, 12), 1468 => to_unsigned(2073, 12), 1469 => to_unsigned(1238, 12), 1470 => to_unsigned(797, 12), 1471 => to_unsigned(3011, 12), 1472 => to_unsigned(2497, 12), 1473 => to_unsigned(2846, 12), 1474 => to_unsigned(3670, 12), 1475 => to_unsigned(3106, 12), 1476 => to_unsigned(2792, 12), 1477 => to_unsigned(875, 12), 1478 => to_unsigned(916, 12), 1479 => to_unsigned(3565, 12), 1480 => to_unsigned(3852, 12), 1481 => to_unsigned(3672, 12), 1482 => to_unsigned(2050, 12), 1483 => to_unsigned(2731, 12), 1484 => to_unsigned(3546, 12), 1485 => to_unsigned(540, 12), 1486 => to_unsigned(702, 12), 1487 => to_unsigned(943, 12), 1488 => to_unsigned(1252, 12), 1489 => to_unsigned(3500, 12), 1490 => to_unsigned(138, 12), 1491 => to_unsigned(3779, 12), 1492 => to_unsigned(2203, 12), 1493 => to_unsigned(3278, 12), 1494 => to_unsigned(1102, 12), 1495 => to_unsigned(2851, 12), 1496 => to_unsigned(927, 12), 1497 => to_unsigned(1195, 12), 1498 => to_unsigned(2080, 12), 1499 => to_unsigned(3157, 12), 1500 => to_unsigned(1959, 12), 1501 => to_unsigned(1300, 12), 1502 => to_unsigned(2273, 12), 1503 => to_unsigned(751, 12), 1504 => to_unsigned(536, 12), 1505 => to_unsigned(805, 12), 1506 => to_unsigned(2822, 12), 1507 => to_unsigned(2085, 12), 1508 => to_unsigned(1075, 12), 1509 => to_unsigned(62, 12), 1510 => to_unsigned(3892, 12), 1511 => to_unsigned(3996, 12), 1512 => to_unsigned(554, 12), 1513 => to_unsigned(2021, 12), 1514 => to_unsigned(1892, 12), 1515 => to_unsigned(1217, 12), 1516 => to_unsigned(1962, 12), 1517 => to_unsigned(668, 12), 1518 => to_unsigned(2233, 12), 1519 => to_unsigned(428, 12), 1520 => to_unsigned(1289, 12), 1521 => to_unsigned(3158, 12), 1522 => to_unsigned(609, 12), 1523 => to_unsigned(2312, 12), 1524 => to_unsigned(207, 12), 1525 => to_unsigned(4001, 12), 1526 => to_unsigned(888, 12), 1527 => to_unsigned(3193, 12), 1528 => to_unsigned(26, 12), 1529 => to_unsigned(497, 12), 1530 => to_unsigned(3196, 12), 1531 => to_unsigned(2728, 12), 1532 => to_unsigned(2174, 12), 1533 => to_unsigned(3355, 12), 1534 => to_unsigned(84, 12), 1535 => to_unsigned(3556, 12), 1536 => to_unsigned(1879, 12), 1537 => to_unsigned(2895, 12), 1538 => to_unsigned(1747, 12), 1539 => to_unsigned(899, 12), 1540 => to_unsigned(130, 12), 1541 => to_unsigned(1077, 12), 1542 => to_unsigned(4072, 12), 1543 => to_unsigned(2322, 12), 1544 => to_unsigned(3497, 12), 1545 => to_unsigned(3764, 12), 1546 => to_unsigned(1863, 12), 1547 => to_unsigned(3578, 12), 1548 => to_unsigned(163, 12), 1549 => to_unsigned(634, 12), 1550 => to_unsigned(717, 12), 1551 => to_unsigned(2650, 12), 1552 => to_unsigned(2602, 12), 1553 => to_unsigned(1359, 12), 1554 => to_unsigned(2898, 12), 1555 => to_unsigned(3293, 12), 1556 => to_unsigned(109, 12), 1557 => to_unsigned(2882, 12), 1558 => to_unsigned(3427, 12), 1559 => to_unsigned(3967, 12), 1560 => to_unsigned(3101, 12), 1561 => to_unsigned(910, 12), 1562 => to_unsigned(49, 12), 1563 => to_unsigned(2022, 12), 1564 => to_unsigned(2724, 12), 1565 => to_unsigned(43, 12), 1566 => to_unsigned(3405, 12), 1567 => to_unsigned(3596, 12), 1568 => to_unsigned(2334, 12), 1569 => to_unsigned(1328, 12), 1570 => to_unsigned(990, 12), 1571 => to_unsigned(3282, 12), 1572 => to_unsigned(220, 12), 1573 => to_unsigned(396, 12), 1574 => to_unsigned(2428, 12), 1575 => to_unsigned(972, 12), 1576 => to_unsigned(684, 12), 1577 => to_unsigned(2821, 12), 1578 => to_unsigned(1017, 12), 1579 => to_unsigned(1867, 12), 1580 => to_unsigned(889, 12), 1581 => to_unsigned(136, 12), 1582 => to_unsigned(1839, 12), 1583 => to_unsigned(168, 12), 1584 => to_unsigned(1739, 12), 1585 => to_unsigned(1391, 12), 1586 => to_unsigned(438, 12), 1587 => to_unsigned(3921, 12), 1588 => to_unsigned(539, 12), 1589 => to_unsigned(2437, 12), 1590 => to_unsigned(3768, 12), 1591 => to_unsigned(1938, 12), 1592 => to_unsigned(315, 12), 1593 => to_unsigned(3660, 12), 1594 => to_unsigned(767, 12), 1595 => to_unsigned(4016, 12), 1596 => to_unsigned(1712, 12), 1597 => to_unsigned(2226, 12), 1598 => to_unsigned(2479, 12), 1599 => to_unsigned(706, 12), 1600 => to_unsigned(1807, 12), 1601 => to_unsigned(456, 12), 1602 => to_unsigned(1609, 12), 1603 => to_unsigned(3300, 12), 1604 => to_unsigned(1257, 12), 1605 => to_unsigned(3311, 12), 1606 => to_unsigned(60, 12), 1607 => to_unsigned(255, 12), 1608 => to_unsigned(2061, 12), 1609 => to_unsigned(556, 12), 1610 => to_unsigned(2224, 12), 1611 => to_unsigned(3166, 12), 1612 => to_unsigned(2576, 12), 1613 => to_unsigned(2456, 12), 1614 => to_unsigned(2336, 12), 1615 => to_unsigned(2330, 12), 1616 => to_unsigned(1540, 12), 1617 => to_unsigned(885, 12), 1618 => to_unsigned(2543, 12), 1619 => to_unsigned(968, 12), 1620 => to_unsigned(1740, 12), 1621 => to_unsigned(1270, 12), 1622 => to_unsigned(940, 12), 1623 => to_unsigned(268, 12), 1624 => to_unsigned(2297, 12), 1625 => to_unsigned(2588, 12), 1626 => to_unsigned(5, 12), 1627 => to_unsigned(1403, 12), 1628 => to_unsigned(1292, 12), 1629 => to_unsigned(593, 12), 1630 => to_unsigned(936, 12), 1631 => to_unsigned(497, 12), 1632 => to_unsigned(3389, 12), 1633 => to_unsigned(4064, 12), 1634 => to_unsigned(1858, 12), 1635 => to_unsigned(2960, 12), 1636 => to_unsigned(1685, 12), 1637 => to_unsigned(3928, 12), 1638 => to_unsigned(2797, 12), 1639 => to_unsigned(1536, 12), 1640 => to_unsigned(590, 12), 1641 => to_unsigned(571, 12), 1642 => to_unsigned(1472, 12), 1643 => to_unsigned(3684, 12), 1644 => to_unsigned(2794, 12), 1645 => to_unsigned(1653, 12), 1646 => to_unsigned(1735, 12), 1647 => to_unsigned(1654, 12), 1648 => to_unsigned(411, 12), 1649 => to_unsigned(2993, 12), 1650 => to_unsigned(642, 12), 1651 => to_unsigned(622, 12), 1652 => to_unsigned(3252, 12), 1653 => to_unsigned(3879, 12), 1654 => to_unsigned(1024, 12), 1655 => to_unsigned(737, 12), 1656 => to_unsigned(684, 12), 1657 => to_unsigned(1201, 12), 1658 => to_unsigned(1682, 12), 1659 => to_unsigned(3611, 12), 1660 => to_unsigned(1188, 12), 1661 => to_unsigned(1538, 12), 1662 => to_unsigned(3146, 12), 1663 => to_unsigned(450, 12), 1664 => to_unsigned(913, 12), 1665 => to_unsigned(101, 12), 1666 => to_unsigned(2723, 12), 1667 => to_unsigned(1292, 12), 1668 => to_unsigned(499, 12), 1669 => to_unsigned(95, 12), 1670 => to_unsigned(3487, 12), 1671 => to_unsigned(3636, 12), 1672 => to_unsigned(3789, 12), 1673 => to_unsigned(2381, 12), 1674 => to_unsigned(1638, 12), 1675 => to_unsigned(279, 12), 1676 => to_unsigned(336, 12), 1677 => to_unsigned(989, 12), 1678 => to_unsigned(3848, 12), 1679 => to_unsigned(3798, 12), 1680 => to_unsigned(1364, 12), 1681 => to_unsigned(3849, 12), 1682 => to_unsigned(3017, 12), 1683 => to_unsigned(1795, 12), 1684 => to_unsigned(3431, 12), 1685 => to_unsigned(31, 12), 1686 => to_unsigned(3930, 12), 1687 => to_unsigned(928, 12), 1688 => to_unsigned(1671, 12), 1689 => to_unsigned(1833, 12), 1690 => to_unsigned(3716, 12), 1691 => to_unsigned(877, 12), 1692 => to_unsigned(114, 12), 1693 => to_unsigned(1422, 12), 1694 => to_unsigned(3855, 12), 1695 => to_unsigned(1002, 12), 1696 => to_unsigned(1741, 12), 1697 => to_unsigned(1087, 12), 1698 => to_unsigned(3254, 12), 1699 => to_unsigned(2712, 12), 1700 => to_unsigned(657, 12), 1701 => to_unsigned(2412, 12), 1702 => to_unsigned(3717, 12), 1703 => to_unsigned(3828, 12), 1704 => to_unsigned(2029, 12), 1705 => to_unsigned(3005, 12), 1706 => to_unsigned(3705, 12), 1707 => to_unsigned(125, 12), 1708 => to_unsigned(1318, 12), 1709 => to_unsigned(2853, 12), 1710 => to_unsigned(3410, 12), 1711 => to_unsigned(3500, 12), 1712 => to_unsigned(3548, 12), 1713 => to_unsigned(3390, 12), 1714 => to_unsigned(3441, 12), 1715 => to_unsigned(3011, 12), 1716 => to_unsigned(3308, 12), 1717 => to_unsigned(934, 12), 1718 => to_unsigned(3044, 12), 1719 => to_unsigned(1323, 12), 1720 => to_unsigned(3331, 12), 1721 => to_unsigned(3590, 12), 1722 => to_unsigned(2159, 12), 1723 => to_unsigned(1713, 12), 1724 => to_unsigned(2060, 12), 1725 => to_unsigned(21, 12), 1726 => to_unsigned(2448, 12), 1727 => to_unsigned(2412, 12), 1728 => to_unsigned(1721, 12), 1729 => to_unsigned(3954, 12), 1730 => to_unsigned(1545, 12), 1731 => to_unsigned(677, 12), 1732 => to_unsigned(3461, 12), 1733 => to_unsigned(73, 12), 1734 => to_unsigned(2043, 12), 1735 => to_unsigned(1269, 12), 1736 => to_unsigned(2887, 12), 1737 => to_unsigned(2417, 12), 1738 => to_unsigned(2536, 12), 1739 => to_unsigned(3650, 12), 1740 => to_unsigned(1250, 12), 1741 => to_unsigned(2726, 12), 1742 => to_unsigned(3709, 12), 1743 => to_unsigned(3771, 12), 1744 => to_unsigned(1912, 12), 1745 => to_unsigned(3348, 12), 1746 => to_unsigned(2093, 12), 1747 => to_unsigned(1807, 12), 1748 => to_unsigned(3857, 12), 1749 => to_unsigned(3882, 12), 1750 => to_unsigned(2292, 12), 1751 => to_unsigned(3776, 12), 1752 => to_unsigned(1764, 12), 1753 => to_unsigned(2053, 12), 1754 => to_unsigned(2010, 12), 1755 => to_unsigned(2186, 12), 1756 => to_unsigned(3164, 12), 1757 => to_unsigned(1678, 12), 1758 => to_unsigned(1577, 12), 1759 => to_unsigned(3955, 12), 1760 => to_unsigned(3823, 12), 1761 => to_unsigned(3914, 12), 1762 => to_unsigned(2067, 12), 1763 => to_unsigned(1822, 12), 1764 => to_unsigned(2531, 12), 1765 => to_unsigned(896, 12), 1766 => to_unsigned(489, 12), 1767 => to_unsigned(1720, 12), 1768 => to_unsigned(2456, 12), 1769 => to_unsigned(3269, 12), 1770 => to_unsigned(3728, 12), 1771 => to_unsigned(316, 12), 1772 => to_unsigned(1914, 12), 1773 => to_unsigned(244, 12), 1774 => to_unsigned(2259, 12), 1775 => to_unsigned(3564, 12), 1776 => to_unsigned(108, 12), 1777 => to_unsigned(3746, 12), 1778 => to_unsigned(3633, 12), 1779 => to_unsigned(3779, 12), 1780 => to_unsigned(303, 12), 1781 => to_unsigned(1070, 12), 1782 => to_unsigned(1000, 12), 1783 => to_unsigned(4027, 12), 1784 => to_unsigned(2478, 12), 1785 => to_unsigned(986, 12), 1786 => to_unsigned(1986, 12), 1787 => to_unsigned(1298, 12), 1788 => to_unsigned(19, 12), 1789 => to_unsigned(229, 12), 1790 => to_unsigned(3303, 12), 1791 => to_unsigned(1977, 12), 1792 => to_unsigned(2248, 12), 1793 => to_unsigned(440, 12), 1794 => to_unsigned(2666, 12), 1795 => to_unsigned(3928, 12), 1796 => to_unsigned(2108, 12), 1797 => to_unsigned(3944, 12), 1798 => to_unsigned(2286, 12), 1799 => to_unsigned(1411, 12), 1800 => to_unsigned(4059, 12), 1801 => to_unsigned(3729, 12), 1802 => to_unsigned(1689, 12), 1803 => to_unsigned(1935, 12), 1804 => to_unsigned(779, 12), 1805 => to_unsigned(2276, 12), 1806 => to_unsigned(2041, 12), 1807 => to_unsigned(203, 12), 1808 => to_unsigned(3277, 12), 1809 => to_unsigned(1852, 12), 1810 => to_unsigned(469, 12), 1811 => to_unsigned(423, 12), 1812 => to_unsigned(3145, 12), 1813 => to_unsigned(228, 12), 1814 => to_unsigned(877, 12), 1815 => to_unsigned(1138, 12), 1816 => to_unsigned(2859, 12), 1817 => to_unsigned(3121, 12), 1818 => to_unsigned(2215, 12), 1819 => to_unsigned(2688, 12), 1820 => to_unsigned(1311, 12), 1821 => to_unsigned(791, 12), 1822 => to_unsigned(1645, 12), 1823 => to_unsigned(2029, 12), 1824 => to_unsigned(3978, 12), 1825 => to_unsigned(671, 12), 1826 => to_unsigned(336, 12), 1827 => to_unsigned(3199, 12), 1828 => to_unsigned(3436, 12), 1829 => to_unsigned(1906, 12), 1830 => to_unsigned(2381, 12), 1831 => to_unsigned(2938, 12), 1832 => to_unsigned(1243, 12), 1833 => to_unsigned(2470, 12), 1834 => to_unsigned(290, 12), 1835 => to_unsigned(1419, 12), 1836 => to_unsigned(325, 12), 1837 => to_unsigned(38, 12), 1838 => to_unsigned(3320, 12), 1839 => to_unsigned(2501, 12), 1840 => to_unsigned(2928, 12), 1841 => to_unsigned(504, 12), 1842 => to_unsigned(2709, 12), 1843 => to_unsigned(3617, 12), 1844 => to_unsigned(693, 12), 1845 => to_unsigned(2336, 12), 1846 => to_unsigned(3761, 12), 1847 => to_unsigned(682, 12), 1848 => to_unsigned(569, 12), 1849 => to_unsigned(3937, 12), 1850 => to_unsigned(3214, 12), 1851 => to_unsigned(4093, 12), 1852 => to_unsigned(552, 12), 1853 => to_unsigned(2938, 12), 1854 => to_unsigned(3224, 12), 1855 => to_unsigned(1550, 12), 1856 => to_unsigned(2061, 12), 1857 => to_unsigned(116, 12), 1858 => to_unsigned(978, 12), 1859 => to_unsigned(3153, 12), 1860 => to_unsigned(2917, 12), 1861 => to_unsigned(2760, 12), 1862 => to_unsigned(1050, 12), 1863 => to_unsigned(2130, 12), 1864 => to_unsigned(3580, 12), 1865 => to_unsigned(117, 12), 1866 => to_unsigned(1306, 12), 1867 => to_unsigned(679, 12), 1868 => to_unsigned(1982, 12), 1869 => to_unsigned(2336, 12), 1870 => to_unsigned(101, 12), 1871 => to_unsigned(2773, 12), 1872 => to_unsigned(2823, 12), 1873 => to_unsigned(3815, 12), 1874 => to_unsigned(3430, 12), 1875 => to_unsigned(273, 12), 1876 => to_unsigned(599, 12), 1877 => to_unsigned(2101, 12), 1878 => to_unsigned(1787, 12), 1879 => to_unsigned(2963, 12), 1880 => to_unsigned(2724, 12), 1881 => to_unsigned(1480, 12), 1882 => to_unsigned(585, 12), 1883 => to_unsigned(561, 12), 1884 => to_unsigned(893, 12), 1885 => to_unsigned(2977, 12), 1886 => to_unsigned(2219, 12), 1887 => to_unsigned(2693, 12), 1888 => to_unsigned(17, 12), 1889 => to_unsigned(3259, 12), 1890 => to_unsigned(3060, 12), 1891 => to_unsigned(3663, 12), 1892 => to_unsigned(2016, 12), 1893 => to_unsigned(1591, 12), 1894 => to_unsigned(1290, 12), 1895 => to_unsigned(1482, 12), 1896 => to_unsigned(1966, 12), 1897 => to_unsigned(3061, 12), 1898 => to_unsigned(1189, 12), 1899 => to_unsigned(614, 12), 1900 => to_unsigned(2000, 12), 1901 => to_unsigned(4, 12), 1902 => to_unsigned(2469, 12), 1903 => to_unsigned(2729, 12), 1904 => to_unsigned(310, 12), 1905 => to_unsigned(169, 12), 1906 => to_unsigned(3150, 12), 1907 => to_unsigned(1177, 12), 1908 => to_unsigned(1317, 12), 1909 => to_unsigned(1714, 12), 1910 => to_unsigned(628, 12), 1911 => to_unsigned(2940, 12), 1912 => to_unsigned(870, 12), 1913 => to_unsigned(2096, 12), 1914 => to_unsigned(3867, 12), 1915 => to_unsigned(857, 12), 1916 => to_unsigned(756, 12), 1917 => to_unsigned(2627, 12), 1918 => to_unsigned(559, 12), 1919 => to_unsigned(2227, 12), 1920 => to_unsigned(1176, 12), 1921 => to_unsigned(3344, 12), 1922 => to_unsigned(2073, 12), 1923 => to_unsigned(1132, 12), 1924 => to_unsigned(1633, 12), 1925 => to_unsigned(1204, 12), 1926 => to_unsigned(3235, 12), 1927 => to_unsigned(2835, 12), 1928 => to_unsigned(2043, 12), 1929 => to_unsigned(642, 12), 1930 => to_unsigned(633, 12), 1931 => to_unsigned(2764, 12), 1932 => to_unsigned(3954, 12), 1933 => to_unsigned(4030, 12), 1934 => to_unsigned(2721, 12), 1935 => to_unsigned(3000, 12), 1936 => to_unsigned(2572, 12), 1937 => to_unsigned(2888, 12), 1938 => to_unsigned(3131, 12), 1939 => to_unsigned(1750, 12), 1940 => to_unsigned(1597, 12), 1941 => to_unsigned(1391, 12), 1942 => to_unsigned(240, 12), 1943 => to_unsigned(1993, 12), 1944 => to_unsigned(3752, 12), 1945 => to_unsigned(2844, 12), 1946 => to_unsigned(123, 12), 1947 => to_unsigned(1881, 12), 1948 => to_unsigned(414, 12), 1949 => to_unsigned(1528, 12), 1950 => to_unsigned(3878, 12), 1951 => to_unsigned(895, 12), 1952 => to_unsigned(502, 12), 1953 => to_unsigned(3651, 12), 1954 => to_unsigned(3914, 12), 1955 => to_unsigned(3337, 12), 1956 => to_unsigned(63, 12), 1957 => to_unsigned(2173, 12), 1958 => to_unsigned(1011, 12), 1959 => to_unsigned(760, 12), 1960 => to_unsigned(2077, 12), 1961 => to_unsigned(623, 12), 1962 => to_unsigned(2436, 12), 1963 => to_unsigned(162, 12), 1964 => to_unsigned(3517, 12), 1965 => to_unsigned(2158, 12), 1966 => to_unsigned(1127, 12), 1967 => to_unsigned(2343, 12), 1968 => to_unsigned(2338, 12), 1969 => to_unsigned(3056, 12), 1970 => to_unsigned(1032, 12), 1971 => to_unsigned(3671, 12), 1972 => to_unsigned(683, 12), 1973 => to_unsigned(602, 12), 1974 => to_unsigned(3629, 12), 1975 => to_unsigned(2235, 12), 1976 => to_unsigned(1666, 12), 1977 => to_unsigned(295, 12), 1978 => to_unsigned(2462, 12), 1979 => to_unsigned(65, 12), 1980 => to_unsigned(3605, 12), 1981 => to_unsigned(2122, 12), 1982 => to_unsigned(1195, 12), 1983 => to_unsigned(3591, 12), 1984 => to_unsigned(1064, 12), 1985 => to_unsigned(1761, 12), 1986 => to_unsigned(2625, 12), 1987 => to_unsigned(3177, 12), 1988 => to_unsigned(3018, 12), 1989 => to_unsigned(2175, 12), 1990 => to_unsigned(1954, 12), 1991 => to_unsigned(2074, 12), 1992 => to_unsigned(2378, 12), 1993 => to_unsigned(3481, 12), 1994 => to_unsigned(2456, 12), 1995 => to_unsigned(3670, 12), 1996 => to_unsigned(3502, 12), 1997 => to_unsigned(510, 12), 1998 => to_unsigned(907, 12), 1999 => to_unsigned(1689, 12), 2000 => to_unsigned(3356, 12), 2001 => to_unsigned(2017, 12), 2002 => to_unsigned(204, 12), 2003 => to_unsigned(573, 12), 2004 => to_unsigned(164, 12), 2005 => to_unsigned(3125, 12), 2006 => to_unsigned(2865, 12), 2007 => to_unsigned(3503, 12), 2008 => to_unsigned(1534, 12), 2009 => to_unsigned(2358, 12), 2010 => to_unsigned(3320, 12), 2011 => to_unsigned(1249, 12), 2012 => to_unsigned(1492, 12), 2013 => to_unsigned(919, 12), 2014 => to_unsigned(674, 12), 2015 => to_unsigned(710, 12), 2016 => to_unsigned(3899, 12), 2017 => to_unsigned(1949, 12), 2018 => to_unsigned(1190, 12), 2019 => to_unsigned(3737, 12), 2020 => to_unsigned(2959, 12), 2021 => to_unsigned(3274, 12), 2022 => to_unsigned(647, 12), 2023 => to_unsigned(1524, 12), 2024 => to_unsigned(195, 12), 2025 => to_unsigned(3562, 12), 2026 => to_unsigned(2628, 12), 2027 => to_unsigned(2871, 12), 2028 => to_unsigned(800, 12), 2029 => to_unsigned(3037, 12), 2030 => to_unsigned(2916, 12), 2031 => to_unsigned(1270, 12), 2032 => to_unsigned(50, 12), 2033 => to_unsigned(250, 12), 2034 => to_unsigned(3332, 12), 2035 => to_unsigned(3753, 12), 2036 => to_unsigned(2921, 12), 2037 => to_unsigned(2827, 12), 2038 => to_unsigned(1548, 12), 2039 => to_unsigned(3334, 12), 2040 => to_unsigned(793, 12), 2041 => to_unsigned(1231, 12), 2042 => to_unsigned(1888, 12), 2043 => to_unsigned(3118, 12), 2044 => to_unsigned(2390, 12), 2045 => to_unsigned(1463, 12), 2046 => to_unsigned(448, 12), 2047 => to_unsigned(3445, 12)),
            3 => (0 => to_unsigned(2219, 12), 1 => to_unsigned(649, 12), 2 => to_unsigned(594, 12), 3 => to_unsigned(357, 12), 4 => to_unsigned(2285, 12), 5 => to_unsigned(2947, 12), 6 => to_unsigned(3994, 12), 7 => to_unsigned(1572, 12), 8 => to_unsigned(3080, 12), 9 => to_unsigned(3154, 12), 10 => to_unsigned(1246, 12), 11 => to_unsigned(3920, 12), 12 => to_unsigned(2796, 12), 13 => to_unsigned(1448, 12), 14 => to_unsigned(2215, 12), 15 => to_unsigned(1261, 12), 16 => to_unsigned(3508, 12), 17 => to_unsigned(2485, 12), 18 => to_unsigned(542, 12), 19 => to_unsigned(2215, 12), 20 => to_unsigned(2122, 12), 21 => to_unsigned(1771, 12), 22 => to_unsigned(1522, 12), 23 => to_unsigned(2196, 12), 24 => to_unsigned(546, 12), 25 => to_unsigned(873, 12), 26 => to_unsigned(3650, 12), 27 => to_unsigned(3679, 12), 28 => to_unsigned(518, 12), 29 => to_unsigned(1468, 12), 30 => to_unsigned(327, 12), 31 => to_unsigned(864, 12), 32 => to_unsigned(2726, 12), 33 => to_unsigned(1125, 12), 34 => to_unsigned(2860, 12), 35 => to_unsigned(708, 12), 36 => to_unsigned(3573, 12), 37 => to_unsigned(1468, 12), 38 => to_unsigned(1265, 12), 39 => to_unsigned(23, 12), 40 => to_unsigned(2989, 12), 41 => to_unsigned(3237, 12), 42 => to_unsigned(664, 12), 43 => to_unsigned(3258, 12), 44 => to_unsigned(3550, 12), 45 => to_unsigned(52, 12), 46 => to_unsigned(2149, 12), 47 => to_unsigned(322, 12), 48 => to_unsigned(3070, 12), 49 => to_unsigned(348, 12), 50 => to_unsigned(1982, 12), 51 => to_unsigned(1226, 12), 52 => to_unsigned(967, 12), 53 => to_unsigned(1798, 12), 54 => to_unsigned(2008, 12), 55 => to_unsigned(452, 12), 56 => to_unsigned(3718, 12), 57 => to_unsigned(906, 12), 58 => to_unsigned(962, 12), 59 => to_unsigned(473, 12), 60 => to_unsigned(1778, 12), 61 => to_unsigned(1628, 12), 62 => to_unsigned(160, 12), 63 => to_unsigned(591, 12), 64 => to_unsigned(2877, 12), 65 => to_unsigned(3022, 12), 66 => to_unsigned(1793, 12), 67 => to_unsigned(3852, 12), 68 => to_unsigned(1363, 12), 69 => to_unsigned(2073, 12), 70 => to_unsigned(2637, 12), 71 => to_unsigned(1091, 12), 72 => to_unsigned(2027, 12), 73 => to_unsigned(846, 12), 74 => to_unsigned(1814, 12), 75 => to_unsigned(234, 12), 76 => to_unsigned(1843, 12), 77 => to_unsigned(799, 12), 78 => to_unsigned(274, 12), 79 => to_unsigned(3120, 12), 80 => to_unsigned(1413, 12), 81 => to_unsigned(1675, 12), 82 => to_unsigned(3701, 12), 83 => to_unsigned(1731, 12), 84 => to_unsigned(1658, 12), 85 => to_unsigned(3379, 12), 86 => to_unsigned(2343, 12), 87 => to_unsigned(1996, 12), 88 => to_unsigned(3975, 12), 89 => to_unsigned(888, 12), 90 => to_unsigned(3522, 12), 91 => to_unsigned(2153, 12), 92 => to_unsigned(2745, 12), 93 => to_unsigned(699, 12), 94 => to_unsigned(2221, 12), 95 => to_unsigned(169, 12), 96 => to_unsigned(591, 12), 97 => to_unsigned(3865, 12), 98 => to_unsigned(3512, 12), 99 => to_unsigned(2040, 12), 100 => to_unsigned(27, 12), 101 => to_unsigned(2712, 12), 102 => to_unsigned(1277, 12), 103 => to_unsigned(2630, 12), 104 => to_unsigned(2601, 12), 105 => to_unsigned(1838, 12), 106 => to_unsigned(489, 12), 107 => to_unsigned(2883, 12), 108 => to_unsigned(68, 12), 109 => to_unsigned(2613, 12), 110 => to_unsigned(3856, 12), 111 => to_unsigned(3156, 12), 112 => to_unsigned(938, 12), 113 => to_unsigned(1262, 12), 114 => to_unsigned(1642, 12), 115 => to_unsigned(224, 12), 116 => to_unsigned(2820, 12), 117 => to_unsigned(2561, 12), 118 => to_unsigned(1875, 12), 119 => to_unsigned(2906, 12), 120 => to_unsigned(2577, 12), 121 => to_unsigned(2957, 12), 122 => to_unsigned(872, 12), 123 => to_unsigned(1048, 12), 124 => to_unsigned(1261, 12), 125 => to_unsigned(1873, 12), 126 => to_unsigned(1136, 12), 127 => to_unsigned(1287, 12), 128 => to_unsigned(3769, 12), 129 => to_unsigned(1420, 12), 130 => to_unsigned(932, 12), 131 => to_unsigned(4040, 12), 132 => to_unsigned(2322, 12), 133 => to_unsigned(2254, 12), 134 => to_unsigned(3448, 12), 135 => to_unsigned(2225, 12), 136 => to_unsigned(3525, 12), 137 => to_unsigned(250, 12), 138 => to_unsigned(1542, 12), 139 => to_unsigned(983, 12), 140 => to_unsigned(2760, 12), 141 => to_unsigned(845, 12), 142 => to_unsigned(916, 12), 143 => to_unsigned(3303, 12), 144 => to_unsigned(1648, 12), 145 => to_unsigned(1739, 12), 146 => to_unsigned(2521, 12), 147 => to_unsigned(756, 12), 148 => to_unsigned(3149, 12), 149 => to_unsigned(705, 12), 150 => to_unsigned(3589, 12), 151 => to_unsigned(2755, 12), 152 => to_unsigned(2812, 12), 153 => to_unsigned(528, 12), 154 => to_unsigned(878, 12), 155 => to_unsigned(2170, 12), 156 => to_unsigned(4064, 12), 157 => to_unsigned(3156, 12), 158 => to_unsigned(2475, 12), 159 => to_unsigned(2668, 12), 160 => to_unsigned(2273, 12), 161 => to_unsigned(2560, 12), 162 => to_unsigned(1263, 12), 163 => to_unsigned(2349, 12), 164 => to_unsigned(15, 12), 165 => to_unsigned(3472, 12), 166 => to_unsigned(4010, 12), 167 => to_unsigned(2306, 12), 168 => to_unsigned(2576, 12), 169 => to_unsigned(3540, 12), 170 => to_unsigned(2085, 12), 171 => to_unsigned(172, 12), 172 => to_unsigned(165, 12), 173 => to_unsigned(2346, 12), 174 => to_unsigned(3201, 12), 175 => to_unsigned(2918, 12), 176 => to_unsigned(754, 12), 177 => to_unsigned(58, 12), 178 => to_unsigned(642, 12), 179 => to_unsigned(1422, 12), 180 => to_unsigned(233, 12), 181 => to_unsigned(716, 12), 182 => to_unsigned(4058, 12), 183 => to_unsigned(160, 12), 184 => to_unsigned(1903, 12), 185 => to_unsigned(4059, 12), 186 => to_unsigned(198, 12), 187 => to_unsigned(2474, 12), 188 => to_unsigned(2107, 12), 189 => to_unsigned(1256, 12), 190 => to_unsigned(1501, 12), 191 => to_unsigned(871, 12), 192 => to_unsigned(1771, 12), 193 => to_unsigned(3367, 12), 194 => to_unsigned(4049, 12), 195 => to_unsigned(1326, 12), 196 => to_unsigned(232, 12), 197 => to_unsigned(605, 12), 198 => to_unsigned(436, 12), 199 => to_unsigned(560, 12), 200 => to_unsigned(3273, 12), 201 => to_unsigned(245, 12), 202 => to_unsigned(2897, 12), 203 => to_unsigned(1727, 12), 204 => to_unsigned(2762, 12), 205 => to_unsigned(396, 12), 206 => to_unsigned(1405, 12), 207 => to_unsigned(1519, 12), 208 => to_unsigned(3710, 12), 209 => to_unsigned(991, 12), 210 => to_unsigned(641, 12), 211 => to_unsigned(2329, 12), 212 => to_unsigned(152, 12), 213 => to_unsigned(589, 12), 214 => to_unsigned(233, 12), 215 => to_unsigned(222, 12), 216 => to_unsigned(241, 12), 217 => to_unsigned(3884, 12), 218 => to_unsigned(3639, 12), 219 => to_unsigned(3946, 12), 220 => to_unsigned(1960, 12), 221 => to_unsigned(3061, 12), 222 => to_unsigned(236, 12), 223 => to_unsigned(2334, 12), 224 => to_unsigned(1465, 12), 225 => to_unsigned(1555, 12), 226 => to_unsigned(2780, 12), 227 => to_unsigned(944, 12), 228 => to_unsigned(3334, 12), 229 => to_unsigned(3948, 12), 230 => to_unsigned(2122, 12), 231 => to_unsigned(1270, 12), 232 => to_unsigned(680, 12), 233 => to_unsigned(2003, 12), 234 => to_unsigned(1648, 12), 235 => to_unsigned(2872, 12), 236 => to_unsigned(1286, 12), 237 => to_unsigned(3621, 12), 238 => to_unsigned(3024, 12), 239 => to_unsigned(5, 12), 240 => to_unsigned(3490, 12), 241 => to_unsigned(908, 12), 242 => to_unsigned(861, 12), 243 => to_unsigned(882, 12), 244 => to_unsigned(1812, 12), 245 => to_unsigned(2141, 12), 246 => to_unsigned(2314, 12), 247 => to_unsigned(3547, 12), 248 => to_unsigned(3378, 12), 249 => to_unsigned(1788, 12), 250 => to_unsigned(1249, 12), 251 => to_unsigned(2538, 12), 252 => to_unsigned(1482, 12), 253 => to_unsigned(1245, 12), 254 => to_unsigned(3594, 12), 255 => to_unsigned(3983, 12), 256 => to_unsigned(2230, 12), 257 => to_unsigned(2705, 12), 258 => to_unsigned(3421, 12), 259 => to_unsigned(3920, 12), 260 => to_unsigned(2872, 12), 261 => to_unsigned(76, 12), 262 => to_unsigned(3036, 12), 263 => to_unsigned(772, 12), 264 => to_unsigned(1286, 12), 265 => to_unsigned(3693, 12), 266 => to_unsigned(958, 12), 267 => to_unsigned(1399, 12), 268 => to_unsigned(3122, 12), 269 => to_unsigned(2609, 12), 270 => to_unsigned(3884, 12), 271 => to_unsigned(170, 12), 272 => to_unsigned(3230, 12), 273 => to_unsigned(2387, 12), 274 => to_unsigned(1682, 12), 275 => to_unsigned(4002, 12), 276 => to_unsigned(285, 12), 277 => to_unsigned(2894, 12), 278 => to_unsigned(2958, 12), 279 => to_unsigned(2540, 12), 280 => to_unsigned(1786, 12), 281 => to_unsigned(2178, 12), 282 => to_unsigned(1274, 12), 283 => to_unsigned(2241, 12), 284 => to_unsigned(2951, 12), 285 => to_unsigned(369, 12), 286 => to_unsigned(2338, 12), 287 => to_unsigned(3544, 12), 288 => to_unsigned(3999, 12), 289 => to_unsigned(109, 12), 290 => to_unsigned(1729, 12), 291 => to_unsigned(1404, 12), 292 => to_unsigned(2404, 12), 293 => to_unsigned(325, 12), 294 => to_unsigned(2212, 12), 295 => to_unsigned(521, 12), 296 => to_unsigned(3511, 12), 297 => to_unsigned(1095, 12), 298 => to_unsigned(54, 12), 299 => to_unsigned(195, 12), 300 => to_unsigned(2449, 12), 301 => to_unsigned(2658, 12), 302 => to_unsigned(3690, 12), 303 => to_unsigned(2904, 12), 304 => to_unsigned(1853, 12), 305 => to_unsigned(2735, 12), 306 => to_unsigned(1886, 12), 307 => to_unsigned(868, 12), 308 => to_unsigned(3880, 12), 309 => to_unsigned(1695, 12), 310 => to_unsigned(9, 12), 311 => to_unsigned(363, 12), 312 => to_unsigned(3088, 12), 313 => to_unsigned(2002, 12), 314 => to_unsigned(1430, 12), 315 => to_unsigned(2633, 12), 316 => to_unsigned(2175, 12), 317 => to_unsigned(1053, 12), 318 => to_unsigned(2883, 12), 319 => to_unsigned(196, 12), 320 => to_unsigned(905, 12), 321 => to_unsigned(1781, 12), 322 => to_unsigned(464, 12), 323 => to_unsigned(4058, 12), 324 => to_unsigned(671, 12), 325 => to_unsigned(1223, 12), 326 => to_unsigned(536, 12), 327 => to_unsigned(2129, 12), 328 => to_unsigned(1638, 12), 329 => to_unsigned(3329, 12), 330 => to_unsigned(3813, 12), 331 => to_unsigned(1307, 12), 332 => to_unsigned(2724, 12), 333 => to_unsigned(1862, 12), 334 => to_unsigned(3642, 12), 335 => to_unsigned(3405, 12), 336 => to_unsigned(2053, 12), 337 => to_unsigned(3312, 12), 338 => to_unsigned(951, 12), 339 => to_unsigned(2840, 12), 340 => to_unsigned(3590, 12), 341 => to_unsigned(3054, 12), 342 => to_unsigned(1386, 12), 343 => to_unsigned(2801, 12), 344 => to_unsigned(3958, 12), 345 => to_unsigned(3537, 12), 346 => to_unsigned(3068, 12), 347 => to_unsigned(3762, 12), 348 => to_unsigned(3405, 12), 349 => to_unsigned(486, 12), 350 => to_unsigned(837, 12), 351 => to_unsigned(1640, 12), 352 => to_unsigned(2310, 12), 353 => to_unsigned(852, 12), 354 => to_unsigned(307, 12), 355 => to_unsigned(2460, 12), 356 => to_unsigned(1197, 12), 357 => to_unsigned(1757, 12), 358 => to_unsigned(2481, 12), 359 => to_unsigned(1823, 12), 360 => to_unsigned(376, 12), 361 => to_unsigned(1001, 12), 362 => to_unsigned(293, 12), 363 => to_unsigned(2431, 12), 364 => to_unsigned(3291, 12), 365 => to_unsigned(2744, 12), 366 => to_unsigned(3008, 12), 367 => to_unsigned(42, 12), 368 => to_unsigned(2773, 12), 369 => to_unsigned(3752, 12), 370 => to_unsigned(3787, 12), 371 => to_unsigned(1541, 12), 372 => to_unsigned(2921, 12), 373 => to_unsigned(10, 12), 374 => to_unsigned(930, 12), 375 => to_unsigned(2008, 12), 376 => to_unsigned(779, 12), 377 => to_unsigned(1442, 12), 378 => to_unsigned(3743, 12), 379 => to_unsigned(2244, 12), 380 => to_unsigned(3483, 12), 381 => to_unsigned(3111, 12), 382 => to_unsigned(3988, 12), 383 => to_unsigned(1433, 12), 384 => to_unsigned(3522, 12), 385 => to_unsigned(1281, 12), 386 => to_unsigned(2281, 12), 387 => to_unsigned(1935, 12), 388 => to_unsigned(915, 12), 389 => to_unsigned(1326, 12), 390 => to_unsigned(2388, 12), 391 => to_unsigned(2016, 12), 392 => to_unsigned(974, 12), 393 => to_unsigned(3116, 12), 394 => to_unsigned(873, 12), 395 => to_unsigned(1159, 12), 396 => to_unsigned(1161, 12), 397 => to_unsigned(908, 12), 398 => to_unsigned(851, 12), 399 => to_unsigned(2360, 12), 400 => to_unsigned(2342, 12), 401 => to_unsigned(3885, 12), 402 => to_unsigned(739, 12), 403 => to_unsigned(1966, 12), 404 => to_unsigned(688, 12), 405 => to_unsigned(2873, 12), 406 => to_unsigned(1682, 12), 407 => to_unsigned(3506, 12), 408 => to_unsigned(1187, 12), 409 => to_unsigned(2312, 12), 410 => to_unsigned(3070, 12), 411 => to_unsigned(3558, 12), 412 => to_unsigned(3543, 12), 413 => to_unsigned(16, 12), 414 => to_unsigned(2312, 12), 415 => to_unsigned(2747, 12), 416 => to_unsigned(373, 12), 417 => to_unsigned(3308, 12), 418 => to_unsigned(3635, 12), 419 => to_unsigned(280, 12), 420 => to_unsigned(1932, 12), 421 => to_unsigned(1576, 12), 422 => to_unsigned(2581, 12), 423 => to_unsigned(475, 12), 424 => to_unsigned(921, 12), 425 => to_unsigned(1953, 12), 426 => to_unsigned(3916, 12), 427 => to_unsigned(756, 12), 428 => to_unsigned(3435, 12), 429 => to_unsigned(2537, 12), 430 => to_unsigned(3586, 12), 431 => to_unsigned(1059, 12), 432 => to_unsigned(408, 12), 433 => to_unsigned(839, 12), 434 => to_unsigned(1291, 12), 435 => to_unsigned(312, 12), 436 => to_unsigned(2087, 12), 437 => to_unsigned(3407, 12), 438 => to_unsigned(808, 12), 439 => to_unsigned(3019, 12), 440 => to_unsigned(2274, 12), 441 => to_unsigned(3425, 12), 442 => to_unsigned(1318, 12), 443 => to_unsigned(2544, 12), 444 => to_unsigned(3716, 12), 445 => to_unsigned(460, 12), 446 => to_unsigned(3746, 12), 447 => to_unsigned(3228, 12), 448 => to_unsigned(2413, 12), 449 => to_unsigned(4045, 12), 450 => to_unsigned(111, 12), 451 => to_unsigned(677, 12), 452 => to_unsigned(1354, 12), 453 => to_unsigned(482, 12), 454 => to_unsigned(955, 12), 455 => to_unsigned(2275, 12), 456 => to_unsigned(837, 12), 457 => to_unsigned(215, 12), 458 => to_unsigned(1138, 12), 459 => to_unsigned(3097, 12), 460 => to_unsigned(2070, 12), 461 => to_unsigned(414, 12), 462 => to_unsigned(2138, 12), 463 => to_unsigned(1971, 12), 464 => to_unsigned(2989, 12), 465 => to_unsigned(1214, 12), 466 => to_unsigned(354, 12), 467 => to_unsigned(1431, 12), 468 => to_unsigned(3186, 12), 469 => to_unsigned(112, 12), 470 => to_unsigned(3491, 12), 471 => to_unsigned(654, 12), 472 => to_unsigned(2461, 12), 473 => to_unsigned(1358, 12), 474 => to_unsigned(1107, 12), 475 => to_unsigned(2338, 12), 476 => to_unsigned(45, 12), 477 => to_unsigned(1334, 12), 478 => to_unsigned(1121, 12), 479 => to_unsigned(1853, 12), 480 => to_unsigned(1626, 12), 481 => to_unsigned(3908, 12), 482 => to_unsigned(467, 12), 483 => to_unsigned(1133, 12), 484 => to_unsigned(3487, 12), 485 => to_unsigned(1910, 12), 486 => to_unsigned(2846, 12), 487 => to_unsigned(1518, 12), 488 => to_unsigned(3490, 12), 489 => to_unsigned(2423, 12), 490 => to_unsigned(3184, 12), 491 => to_unsigned(545, 12), 492 => to_unsigned(1539, 12), 493 => to_unsigned(3743, 12), 494 => to_unsigned(2962, 12), 495 => to_unsigned(509, 12), 496 => to_unsigned(2160, 12), 497 => to_unsigned(669, 12), 498 => to_unsigned(3873, 12), 499 => to_unsigned(983, 12), 500 => to_unsigned(2237, 12), 501 => to_unsigned(1487, 12), 502 => to_unsigned(861, 12), 503 => to_unsigned(2373, 12), 504 => to_unsigned(389, 12), 505 => to_unsigned(1277, 12), 506 => to_unsigned(2692, 12), 507 => to_unsigned(2957, 12), 508 => to_unsigned(3750, 12), 509 => to_unsigned(1505, 12), 510 => to_unsigned(979, 12), 511 => to_unsigned(1907, 12), 512 => to_unsigned(2462, 12), 513 => to_unsigned(2548, 12), 514 => to_unsigned(3971, 12), 515 => to_unsigned(637, 12), 516 => to_unsigned(477, 12), 517 => to_unsigned(2060, 12), 518 => to_unsigned(2323, 12), 519 => to_unsigned(1551, 12), 520 => to_unsigned(2061, 12), 521 => to_unsigned(2402, 12), 522 => to_unsigned(340, 12), 523 => to_unsigned(283, 12), 524 => to_unsigned(1491, 12), 525 => to_unsigned(350, 12), 526 => to_unsigned(237, 12), 527 => to_unsigned(2131, 12), 528 => to_unsigned(1246, 12), 529 => to_unsigned(3297, 12), 530 => to_unsigned(2547, 12), 531 => to_unsigned(3605, 12), 532 => to_unsigned(2513, 12), 533 => to_unsigned(2371, 12), 534 => to_unsigned(3991, 12), 535 => to_unsigned(2446, 12), 536 => to_unsigned(116, 12), 537 => to_unsigned(55, 12), 538 => to_unsigned(2786, 12), 539 => to_unsigned(3857, 12), 540 => to_unsigned(101, 12), 541 => to_unsigned(2882, 12), 542 => to_unsigned(2774, 12), 543 => to_unsigned(57, 12), 544 => to_unsigned(319, 12), 545 => to_unsigned(2063, 12), 546 => to_unsigned(1542, 12), 547 => to_unsigned(1764, 12), 548 => to_unsigned(1493, 12), 549 => to_unsigned(1227, 12), 550 => to_unsigned(2891, 12), 551 => to_unsigned(3891, 12), 552 => to_unsigned(3182, 12), 553 => to_unsigned(4038, 12), 554 => to_unsigned(3415, 12), 555 => to_unsigned(3986, 12), 556 => to_unsigned(2829, 12), 557 => to_unsigned(1651, 12), 558 => to_unsigned(3191, 12), 559 => to_unsigned(2136, 12), 560 => to_unsigned(327, 12), 561 => to_unsigned(3959, 12), 562 => to_unsigned(3237, 12), 563 => to_unsigned(1250, 12), 564 => to_unsigned(2307, 12), 565 => to_unsigned(3837, 12), 566 => to_unsigned(1714, 12), 567 => to_unsigned(1490, 12), 568 => to_unsigned(919, 12), 569 => to_unsigned(4065, 12), 570 => to_unsigned(2613, 12), 571 => to_unsigned(1093, 12), 572 => to_unsigned(431, 12), 573 => to_unsigned(2270, 12), 574 => to_unsigned(1945, 12), 575 => to_unsigned(2741, 12), 576 => to_unsigned(2289, 12), 577 => to_unsigned(3459, 12), 578 => to_unsigned(1160, 12), 579 => to_unsigned(2697, 12), 580 => to_unsigned(894, 12), 581 => to_unsigned(2136, 12), 582 => to_unsigned(561, 12), 583 => to_unsigned(4012, 12), 584 => to_unsigned(30, 12), 585 => to_unsigned(1483, 12), 586 => to_unsigned(1214, 12), 587 => to_unsigned(1410, 12), 588 => to_unsigned(432, 12), 589 => to_unsigned(2388, 12), 590 => to_unsigned(1199, 12), 591 => to_unsigned(1291, 12), 592 => to_unsigned(1248, 12), 593 => to_unsigned(3868, 12), 594 => to_unsigned(2291, 12), 595 => to_unsigned(613, 12), 596 => to_unsigned(235, 12), 597 => to_unsigned(165, 12), 598 => to_unsigned(2342, 12), 599 => to_unsigned(1974, 12), 600 => to_unsigned(1827, 12), 601 => to_unsigned(2954, 12), 602 => to_unsigned(1471, 12), 603 => to_unsigned(1689, 12), 604 => to_unsigned(2869, 12), 605 => to_unsigned(91, 12), 606 => to_unsigned(2516, 12), 607 => to_unsigned(2106, 12), 608 => to_unsigned(2047, 12), 609 => to_unsigned(973, 12), 610 => to_unsigned(2138, 12), 611 => to_unsigned(406, 12), 612 => to_unsigned(3254, 12), 613 => to_unsigned(3523, 12), 614 => to_unsigned(1558, 12), 615 => to_unsigned(2717, 12), 616 => to_unsigned(2879, 12), 617 => to_unsigned(697, 12), 618 => to_unsigned(2671, 12), 619 => to_unsigned(2802, 12), 620 => to_unsigned(2917, 12), 621 => to_unsigned(1708, 12), 622 => to_unsigned(768, 12), 623 => to_unsigned(2790, 12), 624 => to_unsigned(204, 12), 625 => to_unsigned(207, 12), 626 => to_unsigned(2954, 12), 627 => to_unsigned(492, 12), 628 => to_unsigned(3531, 12), 629 => to_unsigned(3045, 12), 630 => to_unsigned(365, 12), 631 => to_unsigned(2551, 12), 632 => to_unsigned(3793, 12), 633 => to_unsigned(1863, 12), 634 => to_unsigned(277, 12), 635 => to_unsigned(2071, 12), 636 => to_unsigned(2915, 12), 637 => to_unsigned(2570, 12), 638 => to_unsigned(3246, 12), 639 => to_unsigned(1397, 12), 640 => to_unsigned(1809, 12), 641 => to_unsigned(523, 12), 642 => to_unsigned(39, 12), 643 => to_unsigned(1576, 12), 644 => to_unsigned(191, 12), 645 => to_unsigned(1416, 12), 646 => to_unsigned(183, 12), 647 => to_unsigned(3986, 12), 648 => to_unsigned(44, 12), 649 => to_unsigned(1926, 12), 650 => to_unsigned(1508, 12), 651 => to_unsigned(3053, 12), 652 => to_unsigned(2399, 12), 653 => to_unsigned(1553, 12), 654 => to_unsigned(1388, 12), 655 => to_unsigned(1282, 12), 656 => to_unsigned(818, 12), 657 => to_unsigned(2183, 12), 658 => to_unsigned(2133, 12), 659 => to_unsigned(1025, 12), 660 => to_unsigned(2319, 12), 661 => to_unsigned(3526, 12), 662 => to_unsigned(879, 12), 663 => to_unsigned(394, 12), 664 => to_unsigned(4026, 12), 665 => to_unsigned(2761, 12), 666 => to_unsigned(4008, 12), 667 => to_unsigned(1654, 12), 668 => to_unsigned(2104, 12), 669 => to_unsigned(845, 12), 670 => to_unsigned(1094, 12), 671 => to_unsigned(3834, 12), 672 => to_unsigned(3736, 12), 673 => to_unsigned(1034, 12), 674 => to_unsigned(498, 12), 675 => to_unsigned(122, 12), 676 => to_unsigned(430, 12), 677 => to_unsigned(2466, 12), 678 => to_unsigned(704, 12), 679 => to_unsigned(2909, 12), 680 => to_unsigned(3057, 12), 681 => to_unsigned(3613, 12), 682 => to_unsigned(1653, 12), 683 => to_unsigned(3531, 12), 684 => to_unsigned(1497, 12), 685 => to_unsigned(3164, 12), 686 => to_unsigned(2712, 12), 687 => to_unsigned(3023, 12), 688 => to_unsigned(1832, 12), 689 => to_unsigned(1822, 12), 690 => to_unsigned(240, 12), 691 => to_unsigned(1760, 12), 692 => to_unsigned(1148, 12), 693 => to_unsigned(551, 12), 694 => to_unsigned(491, 12), 695 => to_unsigned(1981, 12), 696 => to_unsigned(1889, 12), 697 => to_unsigned(1377, 12), 698 => to_unsigned(2909, 12), 699 => to_unsigned(495, 12), 700 => to_unsigned(1423, 12), 701 => to_unsigned(3957, 12), 702 => to_unsigned(2574, 12), 703 => to_unsigned(1466, 12), 704 => to_unsigned(246, 12), 705 => to_unsigned(3511, 12), 706 => to_unsigned(972, 12), 707 => to_unsigned(277, 12), 708 => to_unsigned(573, 12), 709 => to_unsigned(2180, 12), 710 => to_unsigned(897, 12), 711 => to_unsigned(4051, 12), 712 => to_unsigned(3728, 12), 713 => to_unsigned(279, 12), 714 => to_unsigned(2034, 12), 715 => to_unsigned(2706, 12), 716 => to_unsigned(1019, 12), 717 => to_unsigned(3756, 12), 718 => to_unsigned(1944, 12), 719 => to_unsigned(2648, 12), 720 => to_unsigned(3280, 12), 721 => to_unsigned(3743, 12), 722 => to_unsigned(3232, 12), 723 => to_unsigned(1887, 12), 724 => to_unsigned(1871, 12), 725 => to_unsigned(1428, 12), 726 => to_unsigned(3108, 12), 727 => to_unsigned(3128, 12), 728 => to_unsigned(2974, 12), 729 => to_unsigned(232, 12), 730 => to_unsigned(989, 12), 731 => to_unsigned(2795, 12), 732 => to_unsigned(1909, 12), 733 => to_unsigned(3504, 12), 734 => to_unsigned(3486, 12), 735 => to_unsigned(340, 12), 736 => to_unsigned(176, 12), 737 => to_unsigned(3568, 12), 738 => to_unsigned(307, 12), 739 => to_unsigned(3121, 12), 740 => to_unsigned(1244, 12), 741 => to_unsigned(3832, 12), 742 => to_unsigned(1754, 12), 743 => to_unsigned(3537, 12), 744 => to_unsigned(70, 12), 745 => to_unsigned(1565, 12), 746 => to_unsigned(947, 12), 747 => to_unsigned(897, 12), 748 => to_unsigned(1030, 12), 749 => to_unsigned(950, 12), 750 => to_unsigned(1845, 12), 751 => to_unsigned(2165, 12), 752 => to_unsigned(1581, 12), 753 => to_unsigned(503, 12), 754 => to_unsigned(2433, 12), 755 => to_unsigned(1876, 12), 756 => to_unsigned(1725, 12), 757 => to_unsigned(733, 12), 758 => to_unsigned(1905, 12), 759 => to_unsigned(1257, 12), 760 => to_unsigned(3570, 12), 761 => to_unsigned(145, 12), 762 => to_unsigned(2589, 12), 763 => to_unsigned(614, 12), 764 => to_unsigned(1143, 12), 765 => to_unsigned(1723, 12), 766 => to_unsigned(1351, 12), 767 => to_unsigned(1236, 12), 768 => to_unsigned(987, 12), 769 => to_unsigned(2265, 12), 770 => to_unsigned(776, 12), 771 => to_unsigned(204, 12), 772 => to_unsigned(3031, 12), 773 => to_unsigned(2245, 12), 774 => to_unsigned(509, 12), 775 => to_unsigned(3550, 12), 776 => to_unsigned(3363, 12), 777 => to_unsigned(539, 12), 778 => to_unsigned(249, 12), 779 => to_unsigned(3293, 12), 780 => to_unsigned(1519, 12), 781 => to_unsigned(2780, 12), 782 => to_unsigned(2328, 12), 783 => to_unsigned(458, 12), 784 => to_unsigned(1943, 12), 785 => to_unsigned(3540, 12), 786 => to_unsigned(3836, 12), 787 => to_unsigned(641, 12), 788 => to_unsigned(743, 12), 789 => to_unsigned(262, 12), 790 => to_unsigned(1141, 12), 791 => to_unsigned(3938, 12), 792 => to_unsigned(2265, 12), 793 => to_unsigned(1822, 12), 794 => to_unsigned(654, 12), 795 => to_unsigned(3436, 12), 796 => to_unsigned(3111, 12), 797 => to_unsigned(1898, 12), 798 => to_unsigned(3998, 12), 799 => to_unsigned(146, 12), 800 => to_unsigned(1026, 12), 801 => to_unsigned(147, 12), 802 => to_unsigned(1271, 12), 803 => to_unsigned(3321, 12), 804 => to_unsigned(3901, 12), 805 => to_unsigned(1888, 12), 806 => to_unsigned(1040, 12), 807 => to_unsigned(3815, 12), 808 => to_unsigned(1594, 12), 809 => to_unsigned(3813, 12), 810 => to_unsigned(1064, 12), 811 => to_unsigned(3043, 12), 812 => to_unsigned(1994, 12), 813 => to_unsigned(47, 12), 814 => to_unsigned(97, 12), 815 => to_unsigned(2627, 12), 816 => to_unsigned(2901, 12), 817 => to_unsigned(2189, 12), 818 => to_unsigned(3304, 12), 819 => to_unsigned(292, 12), 820 => to_unsigned(2398, 12), 821 => to_unsigned(3499, 12), 822 => to_unsigned(2641, 12), 823 => to_unsigned(2685, 12), 824 => to_unsigned(2810, 12), 825 => to_unsigned(169, 12), 826 => to_unsigned(3100, 12), 827 => to_unsigned(1900, 12), 828 => to_unsigned(1570, 12), 829 => to_unsigned(1850, 12), 830 => to_unsigned(1530, 12), 831 => to_unsigned(1486, 12), 832 => to_unsigned(892, 12), 833 => to_unsigned(710, 12), 834 => to_unsigned(2007, 12), 835 => to_unsigned(895, 12), 836 => to_unsigned(793, 12), 837 => to_unsigned(1820, 12), 838 => to_unsigned(4084, 12), 839 => to_unsigned(3235, 12), 840 => to_unsigned(1733, 12), 841 => to_unsigned(511, 12), 842 => to_unsigned(3829, 12), 843 => to_unsigned(1769, 12), 844 => to_unsigned(3840, 12), 845 => to_unsigned(2436, 12), 846 => to_unsigned(836, 12), 847 => to_unsigned(2531, 12), 848 => to_unsigned(713, 12), 849 => to_unsigned(3228, 12), 850 => to_unsigned(2285, 12), 851 => to_unsigned(1538, 12), 852 => to_unsigned(2738, 12), 853 => to_unsigned(686, 12), 854 => to_unsigned(2962, 12), 855 => to_unsigned(1751, 12), 856 => to_unsigned(1905, 12), 857 => to_unsigned(375, 12), 858 => to_unsigned(3159, 12), 859 => to_unsigned(37, 12), 860 => to_unsigned(3887, 12), 861 => to_unsigned(2021, 12), 862 => to_unsigned(2982, 12), 863 => to_unsigned(3120, 12), 864 => to_unsigned(1502, 12), 865 => to_unsigned(1968, 12), 866 => to_unsigned(1285, 12), 867 => to_unsigned(3909, 12), 868 => to_unsigned(514, 12), 869 => to_unsigned(1426, 12), 870 => to_unsigned(1043, 12), 871 => to_unsigned(743, 12), 872 => to_unsigned(2076, 12), 873 => to_unsigned(1006, 12), 874 => to_unsigned(1289, 12), 875 => to_unsigned(1018, 12), 876 => to_unsigned(2382, 12), 877 => to_unsigned(3776, 12), 878 => to_unsigned(3851, 12), 879 => to_unsigned(137, 12), 880 => to_unsigned(3262, 12), 881 => to_unsigned(3507, 12), 882 => to_unsigned(2779, 12), 883 => to_unsigned(1483, 12), 884 => to_unsigned(1474, 12), 885 => to_unsigned(2531, 12), 886 => to_unsigned(2764, 12), 887 => to_unsigned(3218, 12), 888 => to_unsigned(1159, 12), 889 => to_unsigned(2113, 12), 890 => to_unsigned(3961, 12), 891 => to_unsigned(3358, 12), 892 => to_unsigned(1927, 12), 893 => to_unsigned(78, 12), 894 => to_unsigned(160, 12), 895 => to_unsigned(1895, 12), 896 => to_unsigned(3425, 12), 897 => to_unsigned(2762, 12), 898 => to_unsigned(1884, 12), 899 => to_unsigned(999, 12), 900 => to_unsigned(1041, 12), 901 => to_unsigned(258, 12), 902 => to_unsigned(3191, 12), 903 => to_unsigned(3479, 12), 904 => to_unsigned(804, 12), 905 => to_unsigned(2410, 12), 906 => to_unsigned(847, 12), 907 => to_unsigned(3334, 12), 908 => to_unsigned(662, 12), 909 => to_unsigned(461, 12), 910 => to_unsigned(2938, 12), 911 => to_unsigned(2264, 12), 912 => to_unsigned(3263, 12), 913 => to_unsigned(1849, 12), 914 => to_unsigned(2138, 12), 915 => to_unsigned(1276, 12), 916 => to_unsigned(2335, 12), 917 => to_unsigned(2325, 12), 918 => to_unsigned(3592, 12), 919 => to_unsigned(1256, 12), 920 => to_unsigned(3141, 12), 921 => to_unsigned(246, 12), 922 => to_unsigned(2585, 12), 923 => to_unsigned(1083, 12), 924 => to_unsigned(585, 12), 925 => to_unsigned(4081, 12), 926 => to_unsigned(1930, 12), 927 => to_unsigned(2575, 12), 928 => to_unsigned(935, 12), 929 => to_unsigned(798, 12), 930 => to_unsigned(1988, 12), 931 => to_unsigned(2792, 12), 932 => to_unsigned(1804, 12), 933 => to_unsigned(2547, 12), 934 => to_unsigned(3909, 12), 935 => to_unsigned(3816, 12), 936 => to_unsigned(3592, 12), 937 => to_unsigned(2909, 12), 938 => to_unsigned(1617, 12), 939 => to_unsigned(3469, 12), 940 => to_unsigned(3018, 12), 941 => to_unsigned(525, 12), 942 => to_unsigned(1283, 12), 943 => to_unsigned(2732, 12), 944 => to_unsigned(1351, 12), 945 => to_unsigned(2890, 12), 946 => to_unsigned(1628, 12), 947 => to_unsigned(1970, 12), 948 => to_unsigned(669, 12), 949 => to_unsigned(339, 12), 950 => to_unsigned(2450, 12), 951 => to_unsigned(1568, 12), 952 => to_unsigned(2787, 12), 953 => to_unsigned(3572, 12), 954 => to_unsigned(3129, 12), 955 => to_unsigned(1746, 12), 956 => to_unsigned(259, 12), 957 => to_unsigned(3283, 12), 958 => to_unsigned(3756, 12), 959 => to_unsigned(242, 12), 960 => to_unsigned(641, 12), 961 => to_unsigned(1307, 12), 962 => to_unsigned(3931, 12), 963 => to_unsigned(3352, 12), 964 => to_unsigned(2356, 12), 965 => to_unsigned(931, 12), 966 => to_unsigned(1757, 12), 967 => to_unsigned(3112, 12), 968 => to_unsigned(1107, 12), 969 => to_unsigned(19, 12), 970 => to_unsigned(3706, 12), 971 => to_unsigned(156, 12), 972 => to_unsigned(2188, 12), 973 => to_unsigned(46, 12), 974 => to_unsigned(2269, 12), 975 => to_unsigned(2116, 12), 976 => to_unsigned(1179, 12), 977 => to_unsigned(1142, 12), 978 => to_unsigned(2877, 12), 979 => to_unsigned(2011, 12), 980 => to_unsigned(3372, 12), 981 => to_unsigned(3792, 12), 982 => to_unsigned(1112, 12), 983 => to_unsigned(2217, 12), 984 => to_unsigned(3909, 12), 985 => to_unsigned(2653, 12), 986 => to_unsigned(3014, 12), 987 => to_unsigned(2312, 12), 988 => to_unsigned(3446, 12), 989 => to_unsigned(3043, 12), 990 => to_unsigned(3055, 12), 991 => to_unsigned(446, 12), 992 => to_unsigned(1417, 12), 993 => to_unsigned(163, 12), 994 => to_unsigned(3661, 12), 995 => to_unsigned(154, 12), 996 => to_unsigned(1736, 12), 997 => to_unsigned(1852, 12), 998 => to_unsigned(637, 12), 999 => to_unsigned(4068, 12), 1000 => to_unsigned(3975, 12), 1001 => to_unsigned(42, 12), 1002 => to_unsigned(2722, 12), 1003 => to_unsigned(1135, 12), 1004 => to_unsigned(987, 12), 1005 => to_unsigned(2359, 12), 1006 => to_unsigned(2036, 12), 1007 => to_unsigned(1614, 12), 1008 => to_unsigned(2455, 12), 1009 => to_unsigned(4057, 12), 1010 => to_unsigned(1317, 12), 1011 => to_unsigned(712, 12), 1012 => to_unsigned(341, 12), 1013 => to_unsigned(1828, 12), 1014 => to_unsigned(2711, 12), 1015 => to_unsigned(2535, 12), 1016 => to_unsigned(2973, 12), 1017 => to_unsigned(140, 12), 1018 => to_unsigned(320, 12), 1019 => to_unsigned(3046, 12), 1020 => to_unsigned(1576, 12), 1021 => to_unsigned(3192, 12), 1022 => to_unsigned(93, 12), 1023 => to_unsigned(1795, 12), 1024 => to_unsigned(2047, 12), 1025 => to_unsigned(2631, 12), 1026 => to_unsigned(2466, 12), 1027 => to_unsigned(1215, 12), 1028 => to_unsigned(3719, 12), 1029 => to_unsigned(3508, 12), 1030 => to_unsigned(2677, 12), 1031 => to_unsigned(3600, 12), 1032 => to_unsigned(114, 12), 1033 => to_unsigned(2640, 12), 1034 => to_unsigned(1313, 12), 1035 => to_unsigned(2346, 12), 1036 => to_unsigned(290, 12), 1037 => to_unsigned(254, 12), 1038 => to_unsigned(2304, 12), 1039 => to_unsigned(3022, 12), 1040 => to_unsigned(1583, 12), 1041 => to_unsigned(38, 12), 1042 => to_unsigned(256, 12), 1043 => to_unsigned(3209, 12), 1044 => to_unsigned(1147, 12), 1045 => to_unsigned(497, 12), 1046 => to_unsigned(1289, 12), 1047 => to_unsigned(682, 12), 1048 => to_unsigned(640, 12), 1049 => to_unsigned(632, 12), 1050 => to_unsigned(574, 12), 1051 => to_unsigned(823, 12), 1052 => to_unsigned(386, 12), 1053 => to_unsigned(1996, 12), 1054 => to_unsigned(2718, 12), 1055 => to_unsigned(44, 12), 1056 => to_unsigned(3278, 12), 1057 => to_unsigned(1693, 12), 1058 => to_unsigned(2819, 12), 1059 => to_unsigned(3492, 12), 1060 => to_unsigned(3500, 12), 1061 => to_unsigned(1108, 12), 1062 => to_unsigned(1896, 12), 1063 => to_unsigned(2251, 12), 1064 => to_unsigned(3063, 12), 1065 => to_unsigned(2444, 12), 1066 => to_unsigned(2771, 12), 1067 => to_unsigned(1407, 12), 1068 => to_unsigned(3530, 12), 1069 => to_unsigned(1436, 12), 1070 => to_unsigned(4034, 12), 1071 => to_unsigned(2588, 12), 1072 => to_unsigned(2650, 12), 1073 => to_unsigned(3262, 12), 1074 => to_unsigned(893, 12), 1075 => to_unsigned(2445, 12), 1076 => to_unsigned(2055, 12), 1077 => to_unsigned(3808, 12), 1078 => to_unsigned(3553, 12), 1079 => to_unsigned(252, 12), 1080 => to_unsigned(2500, 12), 1081 => to_unsigned(1842, 12), 1082 => to_unsigned(113, 12), 1083 => to_unsigned(1538, 12), 1084 => to_unsigned(1217, 12), 1085 => to_unsigned(497, 12), 1086 => to_unsigned(954, 12), 1087 => to_unsigned(2995, 12), 1088 => to_unsigned(2344, 12), 1089 => to_unsigned(767, 12), 1090 => to_unsigned(577, 12), 1091 => to_unsigned(2143, 12), 1092 => to_unsigned(528, 12), 1093 => to_unsigned(3543, 12), 1094 => to_unsigned(383, 12), 1095 => to_unsigned(1628, 12), 1096 => to_unsigned(3485, 12), 1097 => to_unsigned(2602, 12), 1098 => to_unsigned(2825, 12), 1099 => to_unsigned(1497, 12), 1100 => to_unsigned(3435, 12), 1101 => to_unsigned(1652, 12), 1102 => to_unsigned(616, 12), 1103 => to_unsigned(3449, 12), 1104 => to_unsigned(2887, 12), 1105 => to_unsigned(3044, 12), 1106 => to_unsigned(3954, 12), 1107 => to_unsigned(2342, 12), 1108 => to_unsigned(3407, 12), 1109 => to_unsigned(3729, 12), 1110 => to_unsigned(2729, 12), 1111 => to_unsigned(3775, 12), 1112 => to_unsigned(274, 12), 1113 => to_unsigned(1163, 12), 1114 => to_unsigned(3455, 12), 1115 => to_unsigned(1498, 12), 1116 => to_unsigned(2732, 12), 1117 => to_unsigned(1461, 12), 1118 => to_unsigned(2261, 12), 1119 => to_unsigned(3433, 12), 1120 => to_unsigned(2401, 12), 1121 => to_unsigned(2917, 12), 1122 => to_unsigned(2710, 12), 1123 => to_unsigned(623, 12), 1124 => to_unsigned(2583, 12), 1125 => to_unsigned(2539, 12), 1126 => to_unsigned(3730, 12), 1127 => to_unsigned(3909, 12), 1128 => to_unsigned(2297, 12), 1129 => to_unsigned(2946, 12), 1130 => to_unsigned(179, 12), 1131 => to_unsigned(3189, 12), 1132 => to_unsigned(884, 12), 1133 => to_unsigned(1454, 12), 1134 => to_unsigned(3161, 12), 1135 => to_unsigned(2899, 12), 1136 => to_unsigned(2533, 12), 1137 => to_unsigned(3145, 12), 1138 => to_unsigned(152, 12), 1139 => to_unsigned(546, 12), 1140 => to_unsigned(4016, 12), 1141 => to_unsigned(1727, 12), 1142 => to_unsigned(1751, 12), 1143 => to_unsigned(212, 12), 1144 => to_unsigned(1377, 12), 1145 => to_unsigned(721, 12), 1146 => to_unsigned(246, 12), 1147 => to_unsigned(210, 12), 1148 => to_unsigned(1730, 12), 1149 => to_unsigned(1733, 12), 1150 => to_unsigned(4051, 12), 1151 => to_unsigned(1079, 12), 1152 => to_unsigned(2389, 12), 1153 => to_unsigned(177, 12), 1154 => to_unsigned(3574, 12), 1155 => to_unsigned(3680, 12), 1156 => to_unsigned(2637, 12), 1157 => to_unsigned(2742, 12), 1158 => to_unsigned(3179, 12), 1159 => to_unsigned(1608, 12), 1160 => to_unsigned(44, 12), 1161 => to_unsigned(3455, 12), 1162 => to_unsigned(3928, 12), 1163 => to_unsigned(1774, 12), 1164 => to_unsigned(2447, 12), 1165 => to_unsigned(646, 12), 1166 => to_unsigned(693, 12), 1167 => to_unsigned(138, 12), 1168 => to_unsigned(986, 12), 1169 => to_unsigned(2935, 12), 1170 => to_unsigned(2535, 12), 1171 => to_unsigned(1488, 12), 1172 => to_unsigned(4036, 12), 1173 => to_unsigned(2652, 12), 1174 => to_unsigned(2185, 12), 1175 => to_unsigned(757, 12), 1176 => to_unsigned(2158, 12), 1177 => to_unsigned(312, 12), 1178 => to_unsigned(308, 12), 1179 => to_unsigned(3288, 12), 1180 => to_unsigned(1431, 12), 1181 => to_unsigned(1579, 12), 1182 => to_unsigned(1163, 12), 1183 => to_unsigned(3780, 12), 1184 => to_unsigned(244, 12), 1185 => to_unsigned(2844, 12), 1186 => to_unsigned(2914, 12), 1187 => to_unsigned(1430, 12), 1188 => to_unsigned(1247, 12), 1189 => to_unsigned(2599, 12), 1190 => to_unsigned(4050, 12), 1191 => to_unsigned(1880, 12), 1192 => to_unsigned(508, 12), 1193 => to_unsigned(2220, 12), 1194 => to_unsigned(2980, 12), 1195 => to_unsigned(4032, 12), 1196 => to_unsigned(1002, 12), 1197 => to_unsigned(1660, 12), 1198 => to_unsigned(2956, 12), 1199 => to_unsigned(331, 12), 1200 => to_unsigned(3182, 12), 1201 => to_unsigned(1642, 12), 1202 => to_unsigned(1784, 12), 1203 => to_unsigned(4024, 12), 1204 => to_unsigned(2428, 12), 1205 => to_unsigned(2020, 12), 1206 => to_unsigned(1129, 12), 1207 => to_unsigned(168, 12), 1208 => to_unsigned(1611, 12), 1209 => to_unsigned(2275, 12), 1210 => to_unsigned(3813, 12), 1211 => to_unsigned(3443, 12), 1212 => to_unsigned(520, 12), 1213 => to_unsigned(3725, 12), 1214 => to_unsigned(2284, 12), 1215 => to_unsigned(2082, 12), 1216 => to_unsigned(3871, 12), 1217 => to_unsigned(3117, 12), 1218 => to_unsigned(1090, 12), 1219 => to_unsigned(797, 12), 1220 => to_unsigned(880, 12), 1221 => to_unsigned(2246, 12), 1222 => to_unsigned(1913, 12), 1223 => to_unsigned(1856, 12), 1224 => to_unsigned(1021, 12), 1225 => to_unsigned(2045, 12), 1226 => to_unsigned(1521, 12), 1227 => to_unsigned(1599, 12), 1228 => to_unsigned(3283, 12), 1229 => to_unsigned(3864, 12), 1230 => to_unsigned(3579, 12), 1231 => to_unsigned(1952, 12), 1232 => to_unsigned(1570, 12), 1233 => to_unsigned(123, 12), 1234 => to_unsigned(1339, 12), 1235 => to_unsigned(380, 12), 1236 => to_unsigned(950, 12), 1237 => to_unsigned(683, 12), 1238 => to_unsigned(2775, 12), 1239 => to_unsigned(3149, 12), 1240 => to_unsigned(3750, 12), 1241 => to_unsigned(427, 12), 1242 => to_unsigned(1268, 12), 1243 => to_unsigned(3704, 12), 1244 => to_unsigned(929, 12), 1245 => to_unsigned(17, 12), 1246 => to_unsigned(769, 12), 1247 => to_unsigned(2981, 12), 1248 => to_unsigned(2877, 12), 1249 => to_unsigned(2000, 12), 1250 => to_unsigned(2646, 12), 1251 => to_unsigned(2169, 12), 1252 => to_unsigned(2738, 12), 1253 => to_unsigned(224, 12), 1254 => to_unsigned(2779, 12), 1255 => to_unsigned(2190, 12), 1256 => to_unsigned(3658, 12), 1257 => to_unsigned(3222, 12), 1258 => to_unsigned(140, 12), 1259 => to_unsigned(2364, 12), 1260 => to_unsigned(110, 12), 1261 => to_unsigned(74, 12), 1262 => to_unsigned(2339, 12), 1263 => to_unsigned(2149, 12), 1264 => to_unsigned(474, 12), 1265 => to_unsigned(3281, 12), 1266 => to_unsigned(4007, 12), 1267 => to_unsigned(1279, 12), 1268 => to_unsigned(1573, 12), 1269 => to_unsigned(225, 12), 1270 => to_unsigned(2581, 12), 1271 => to_unsigned(2769, 12), 1272 => to_unsigned(3509, 12), 1273 => to_unsigned(3176, 12), 1274 => to_unsigned(1651, 12), 1275 => to_unsigned(337, 12), 1276 => to_unsigned(2188, 12), 1277 => to_unsigned(2022, 12), 1278 => to_unsigned(1871, 12), 1279 => to_unsigned(2567, 12), 1280 => to_unsigned(2337, 12), 1281 => to_unsigned(4095, 12), 1282 => to_unsigned(540, 12), 1283 => to_unsigned(3333, 12), 1284 => to_unsigned(1573, 12), 1285 => to_unsigned(611, 12), 1286 => to_unsigned(175, 12), 1287 => to_unsigned(3134, 12), 1288 => to_unsigned(233, 12), 1289 => to_unsigned(2969, 12), 1290 => to_unsigned(2321, 12), 1291 => to_unsigned(266, 12), 1292 => to_unsigned(1562, 12), 1293 => to_unsigned(541, 12), 1294 => to_unsigned(657, 12), 1295 => to_unsigned(3946, 12), 1296 => to_unsigned(2115, 12), 1297 => to_unsigned(261, 12), 1298 => to_unsigned(3285, 12), 1299 => to_unsigned(833, 12), 1300 => to_unsigned(179, 12), 1301 => to_unsigned(2926, 12), 1302 => to_unsigned(3055, 12), 1303 => to_unsigned(167, 12), 1304 => to_unsigned(3423, 12), 1305 => to_unsigned(3064, 12), 1306 => to_unsigned(486, 12), 1307 => to_unsigned(3505, 12), 1308 => to_unsigned(3220, 12), 1309 => to_unsigned(1543, 12), 1310 => to_unsigned(1112, 12), 1311 => to_unsigned(1384, 12), 1312 => to_unsigned(2787, 12), 1313 => to_unsigned(2499, 12), 1314 => to_unsigned(567, 12), 1315 => to_unsigned(334, 12), 1316 => to_unsigned(3867, 12), 1317 => to_unsigned(1043, 12), 1318 => to_unsigned(229, 12), 1319 => to_unsigned(69, 12), 1320 => to_unsigned(157, 12), 1321 => to_unsigned(2622, 12), 1322 => to_unsigned(2399, 12), 1323 => to_unsigned(3248, 12), 1324 => to_unsigned(1512, 12), 1325 => to_unsigned(3907, 12), 1326 => to_unsigned(3132, 12), 1327 => to_unsigned(1058, 12), 1328 => to_unsigned(3101, 12), 1329 => to_unsigned(3632, 12), 1330 => to_unsigned(1960, 12), 1331 => to_unsigned(3379, 12), 1332 => to_unsigned(3797, 12), 1333 => to_unsigned(1025, 12), 1334 => to_unsigned(2417, 12), 1335 => to_unsigned(1844, 12), 1336 => to_unsigned(1483, 12), 1337 => to_unsigned(2017, 12), 1338 => to_unsigned(993, 12), 1339 => to_unsigned(3789, 12), 1340 => to_unsigned(38, 12), 1341 => to_unsigned(2790, 12), 1342 => to_unsigned(3308, 12), 1343 => to_unsigned(1029, 12), 1344 => to_unsigned(2951, 12), 1345 => to_unsigned(794, 12), 1346 => to_unsigned(1483, 12), 1347 => to_unsigned(497, 12), 1348 => to_unsigned(3668, 12), 1349 => to_unsigned(3575, 12), 1350 => to_unsigned(3557, 12), 1351 => to_unsigned(1539, 12), 1352 => to_unsigned(2136, 12), 1353 => to_unsigned(2936, 12), 1354 => to_unsigned(3242, 12), 1355 => to_unsigned(2391, 12), 1356 => to_unsigned(2187, 12), 1357 => to_unsigned(2106, 12), 1358 => to_unsigned(3868, 12), 1359 => to_unsigned(2402, 12), 1360 => to_unsigned(2750, 12), 1361 => to_unsigned(2617, 12), 1362 => to_unsigned(356, 12), 1363 => to_unsigned(2845, 12), 1364 => to_unsigned(2920, 12), 1365 => to_unsigned(1595, 12), 1366 => to_unsigned(2473, 12), 1367 => to_unsigned(290, 12), 1368 => to_unsigned(1024, 12), 1369 => to_unsigned(3111, 12), 1370 => to_unsigned(1625, 12), 1371 => to_unsigned(508, 12), 1372 => to_unsigned(2978, 12), 1373 => to_unsigned(3636, 12), 1374 => to_unsigned(1513, 12), 1375 => to_unsigned(3526, 12), 1376 => to_unsigned(3843, 12), 1377 => to_unsigned(1220, 12), 1378 => to_unsigned(3323, 12), 1379 => to_unsigned(3878, 12), 1380 => to_unsigned(1162, 12), 1381 => to_unsigned(398, 12), 1382 => to_unsigned(95, 12), 1383 => to_unsigned(1393, 12), 1384 => to_unsigned(2724, 12), 1385 => to_unsigned(3912, 12), 1386 => to_unsigned(1262, 12), 1387 => to_unsigned(1951, 12), 1388 => to_unsigned(2144, 12), 1389 => to_unsigned(57, 12), 1390 => to_unsigned(3542, 12), 1391 => to_unsigned(782, 12), 1392 => to_unsigned(3613, 12), 1393 => to_unsigned(2063, 12), 1394 => to_unsigned(3570, 12), 1395 => to_unsigned(1557, 12), 1396 => to_unsigned(4010, 12), 1397 => to_unsigned(3229, 12), 1398 => to_unsigned(3072, 12), 1399 => to_unsigned(2658, 12), 1400 => to_unsigned(1459, 12), 1401 => to_unsigned(1361, 12), 1402 => to_unsigned(3150, 12), 1403 => to_unsigned(4081, 12), 1404 => to_unsigned(3516, 12), 1405 => to_unsigned(2708, 12), 1406 => to_unsigned(4007, 12), 1407 => to_unsigned(2305, 12), 1408 => to_unsigned(3677, 12), 1409 => to_unsigned(3687, 12), 1410 => to_unsigned(671, 12), 1411 => to_unsigned(667, 12), 1412 => to_unsigned(3018, 12), 1413 => to_unsigned(2111, 12), 1414 => to_unsigned(582, 12), 1415 => to_unsigned(3776, 12), 1416 => to_unsigned(42, 12), 1417 => to_unsigned(2331, 12), 1418 => to_unsigned(102, 12), 1419 => to_unsigned(2194, 12), 1420 => to_unsigned(3634, 12), 1421 => to_unsigned(2214, 12), 1422 => to_unsigned(2591, 12), 1423 => to_unsigned(1330, 12), 1424 => to_unsigned(3056, 12), 1425 => to_unsigned(437, 12), 1426 => to_unsigned(52, 12), 1427 => to_unsigned(3421, 12), 1428 => to_unsigned(3521, 12), 1429 => to_unsigned(3755, 12), 1430 => to_unsigned(3498, 12), 1431 => to_unsigned(932, 12), 1432 => to_unsigned(2258, 12), 1433 => to_unsigned(3225, 12), 1434 => to_unsigned(4085, 12), 1435 => to_unsigned(318, 12), 1436 => to_unsigned(3136, 12), 1437 => to_unsigned(169, 12), 1438 => to_unsigned(1371, 12), 1439 => to_unsigned(374, 12), 1440 => to_unsigned(4026, 12), 1441 => to_unsigned(1113, 12), 1442 => to_unsigned(3175, 12), 1443 => to_unsigned(1826, 12), 1444 => to_unsigned(386, 12), 1445 => to_unsigned(1784, 12), 1446 => to_unsigned(3993, 12), 1447 => to_unsigned(1056, 12), 1448 => to_unsigned(4027, 12), 1449 => to_unsigned(3797, 12), 1450 => to_unsigned(637, 12), 1451 => to_unsigned(3973, 12), 1452 => to_unsigned(2345, 12), 1453 => to_unsigned(3553, 12), 1454 => to_unsigned(2754, 12), 1455 => to_unsigned(1272, 12), 1456 => to_unsigned(848, 12), 1457 => to_unsigned(2821, 12), 1458 => to_unsigned(2857, 12), 1459 => to_unsigned(1659, 12), 1460 => to_unsigned(3844, 12), 1461 => to_unsigned(19, 12), 1462 => to_unsigned(1728, 12), 1463 => to_unsigned(2104, 12), 1464 => to_unsigned(3671, 12), 1465 => to_unsigned(2504, 12), 1466 => to_unsigned(3470, 12), 1467 => to_unsigned(3962, 12), 1468 => to_unsigned(702, 12), 1469 => to_unsigned(3894, 12), 1470 => to_unsigned(932, 12), 1471 => to_unsigned(1617, 12), 1472 => to_unsigned(2745, 12), 1473 => to_unsigned(1529, 12), 1474 => to_unsigned(1557, 12), 1475 => to_unsigned(3786, 12), 1476 => to_unsigned(997, 12), 1477 => to_unsigned(1922, 12), 1478 => to_unsigned(2588, 12), 1479 => to_unsigned(1012, 12), 1480 => to_unsigned(3693, 12), 1481 => to_unsigned(927, 12), 1482 => to_unsigned(1441, 12), 1483 => to_unsigned(1401, 12), 1484 => to_unsigned(3143, 12), 1485 => to_unsigned(865, 12), 1486 => to_unsigned(196, 12), 1487 => to_unsigned(2568, 12), 1488 => to_unsigned(1488, 12), 1489 => to_unsigned(3539, 12), 1490 => to_unsigned(3113, 12), 1491 => to_unsigned(3546, 12), 1492 => to_unsigned(1398, 12), 1493 => to_unsigned(3396, 12), 1494 => to_unsigned(1069, 12), 1495 => to_unsigned(2236, 12), 1496 => to_unsigned(540, 12), 1497 => to_unsigned(3850, 12), 1498 => to_unsigned(1049, 12), 1499 => to_unsigned(121, 12), 1500 => to_unsigned(1238, 12), 1501 => to_unsigned(3409, 12), 1502 => to_unsigned(1137, 12), 1503 => to_unsigned(339, 12), 1504 => to_unsigned(1835, 12), 1505 => to_unsigned(2043, 12), 1506 => to_unsigned(3763, 12), 1507 => to_unsigned(2708, 12), 1508 => to_unsigned(985, 12), 1509 => to_unsigned(3359, 12), 1510 => to_unsigned(3648, 12), 1511 => to_unsigned(2625, 12), 1512 => to_unsigned(2164, 12), 1513 => to_unsigned(963, 12), 1514 => to_unsigned(424, 12), 1515 => to_unsigned(3081, 12), 1516 => to_unsigned(2488, 12), 1517 => to_unsigned(475, 12), 1518 => to_unsigned(1904, 12), 1519 => to_unsigned(2916, 12), 1520 => to_unsigned(2640, 12), 1521 => to_unsigned(925, 12), 1522 => to_unsigned(3589, 12), 1523 => to_unsigned(1034, 12), 1524 => to_unsigned(3639, 12), 1525 => to_unsigned(2826, 12), 1526 => to_unsigned(2561, 12), 1527 => to_unsigned(3475, 12), 1528 => to_unsigned(2337, 12), 1529 => to_unsigned(2425, 12), 1530 => to_unsigned(296, 12), 1531 => to_unsigned(1600, 12), 1532 => to_unsigned(1455, 12), 1533 => to_unsigned(1050, 12), 1534 => to_unsigned(756, 12), 1535 => to_unsigned(436, 12), 1536 => to_unsigned(153, 12), 1537 => to_unsigned(2611, 12), 1538 => to_unsigned(3033, 12), 1539 => to_unsigned(711, 12), 1540 => to_unsigned(3379, 12), 1541 => to_unsigned(1180, 12), 1542 => to_unsigned(656, 12), 1543 => to_unsigned(2336, 12), 1544 => to_unsigned(1536, 12), 1545 => to_unsigned(3479, 12), 1546 => to_unsigned(3160, 12), 1547 => to_unsigned(1718, 12), 1548 => to_unsigned(1073, 12), 1549 => to_unsigned(247, 12), 1550 => to_unsigned(2880, 12), 1551 => to_unsigned(2521, 12), 1552 => to_unsigned(2319, 12), 1553 => to_unsigned(3376, 12), 1554 => to_unsigned(928, 12), 1555 => to_unsigned(1339, 12), 1556 => to_unsigned(3995, 12), 1557 => to_unsigned(3884, 12), 1558 => to_unsigned(54, 12), 1559 => to_unsigned(2583, 12), 1560 => to_unsigned(2979, 12), 1561 => to_unsigned(589, 12), 1562 => to_unsigned(2096, 12), 1563 => to_unsigned(1284, 12), 1564 => to_unsigned(185, 12), 1565 => to_unsigned(1402, 12), 1566 => to_unsigned(3257, 12), 1567 => to_unsigned(3162, 12), 1568 => to_unsigned(3149, 12), 1569 => to_unsigned(2680, 12), 1570 => to_unsigned(791, 12), 1571 => to_unsigned(3373, 12), 1572 => to_unsigned(731, 12), 1573 => to_unsigned(327, 12), 1574 => to_unsigned(2466, 12), 1575 => to_unsigned(2158, 12), 1576 => to_unsigned(2364, 12), 1577 => to_unsigned(3647, 12), 1578 => to_unsigned(2548, 12), 1579 => to_unsigned(3426, 12), 1580 => to_unsigned(1878, 12), 1581 => to_unsigned(2239, 12), 1582 => to_unsigned(1164, 12), 1583 => to_unsigned(2798, 12), 1584 => to_unsigned(208, 12), 1585 => to_unsigned(3806, 12), 1586 => to_unsigned(2697, 12), 1587 => to_unsigned(291, 12), 1588 => to_unsigned(2972, 12), 1589 => to_unsigned(655, 12), 1590 => to_unsigned(3514, 12), 1591 => to_unsigned(3643, 12), 1592 => to_unsigned(1952, 12), 1593 => to_unsigned(2877, 12), 1594 => to_unsigned(1997, 12), 1595 => to_unsigned(3718, 12), 1596 => to_unsigned(416, 12), 1597 => to_unsigned(706, 12), 1598 => to_unsigned(2009, 12), 1599 => to_unsigned(422, 12), 1600 => to_unsigned(2180, 12), 1601 => to_unsigned(2174, 12), 1602 => to_unsigned(214, 12), 1603 => to_unsigned(2169, 12), 1604 => to_unsigned(2144, 12), 1605 => to_unsigned(93, 12), 1606 => to_unsigned(1952, 12), 1607 => to_unsigned(3498, 12), 1608 => to_unsigned(2840, 12), 1609 => to_unsigned(3797, 12), 1610 => to_unsigned(896, 12), 1611 => to_unsigned(1609, 12), 1612 => to_unsigned(2070, 12), 1613 => to_unsigned(2016, 12), 1614 => to_unsigned(998, 12), 1615 => to_unsigned(411, 12), 1616 => to_unsigned(2410, 12), 1617 => to_unsigned(379, 12), 1618 => to_unsigned(1607, 12), 1619 => to_unsigned(3958, 12), 1620 => to_unsigned(1306, 12), 1621 => to_unsigned(3322, 12), 1622 => to_unsigned(316, 12), 1623 => to_unsigned(1924, 12), 1624 => to_unsigned(3662, 12), 1625 => to_unsigned(3511, 12), 1626 => to_unsigned(2872, 12), 1627 => to_unsigned(2543, 12), 1628 => to_unsigned(2197, 12), 1629 => to_unsigned(1975, 12), 1630 => to_unsigned(3554, 12), 1631 => to_unsigned(1395, 12), 1632 => to_unsigned(1629, 12), 1633 => to_unsigned(623, 12), 1634 => to_unsigned(2603, 12), 1635 => to_unsigned(2357, 12), 1636 => to_unsigned(2720, 12), 1637 => to_unsigned(861, 12), 1638 => to_unsigned(763, 12), 1639 => to_unsigned(547, 12), 1640 => to_unsigned(463, 12), 1641 => to_unsigned(2085, 12), 1642 => to_unsigned(1206, 12), 1643 => to_unsigned(3798, 12), 1644 => to_unsigned(3364, 12), 1645 => to_unsigned(548, 12), 1646 => to_unsigned(1435, 12), 1647 => to_unsigned(1997, 12), 1648 => to_unsigned(3967, 12), 1649 => to_unsigned(3834, 12), 1650 => to_unsigned(643, 12), 1651 => to_unsigned(166, 12), 1652 => to_unsigned(2546, 12), 1653 => to_unsigned(4000, 12), 1654 => to_unsigned(3422, 12), 1655 => to_unsigned(3788, 12), 1656 => to_unsigned(163, 12), 1657 => to_unsigned(1225, 12), 1658 => to_unsigned(434, 12), 1659 => to_unsigned(686, 12), 1660 => to_unsigned(2526, 12), 1661 => to_unsigned(116, 12), 1662 => to_unsigned(3673, 12), 1663 => to_unsigned(3447, 12), 1664 => to_unsigned(3390, 12), 1665 => to_unsigned(2829, 12), 1666 => to_unsigned(1795, 12), 1667 => to_unsigned(3104, 12), 1668 => to_unsigned(942, 12), 1669 => to_unsigned(3660, 12), 1670 => to_unsigned(1647, 12), 1671 => to_unsigned(2231, 12), 1672 => to_unsigned(2024, 12), 1673 => to_unsigned(3836, 12), 1674 => to_unsigned(892, 12), 1675 => to_unsigned(2107, 12), 1676 => to_unsigned(433, 12), 1677 => to_unsigned(1953, 12), 1678 => to_unsigned(1450, 12), 1679 => to_unsigned(2082, 12), 1680 => to_unsigned(1371, 12), 1681 => to_unsigned(2910, 12), 1682 => to_unsigned(3101, 12), 1683 => to_unsigned(2847, 12), 1684 => to_unsigned(588, 12), 1685 => to_unsigned(3112, 12), 1686 => to_unsigned(3425, 12), 1687 => to_unsigned(2055, 12), 1688 => to_unsigned(1449, 12), 1689 => to_unsigned(1780, 12), 1690 => to_unsigned(536, 12), 1691 => to_unsigned(2592, 12), 1692 => to_unsigned(3977, 12), 1693 => to_unsigned(743, 12), 1694 => to_unsigned(3745, 12), 1695 => to_unsigned(2993, 12), 1696 => to_unsigned(2795, 12), 1697 => to_unsigned(1632, 12), 1698 => to_unsigned(1348, 12), 1699 => to_unsigned(4076, 12), 1700 => to_unsigned(1754, 12), 1701 => to_unsigned(327, 12), 1702 => to_unsigned(2546, 12), 1703 => to_unsigned(1971, 12), 1704 => to_unsigned(838, 12), 1705 => to_unsigned(3477, 12), 1706 => to_unsigned(3629, 12), 1707 => to_unsigned(1179, 12), 1708 => to_unsigned(8, 12), 1709 => to_unsigned(3389, 12), 1710 => to_unsigned(3068, 12), 1711 => to_unsigned(2142, 12), 1712 => to_unsigned(3587, 12), 1713 => to_unsigned(2116, 12), 1714 => to_unsigned(780, 12), 1715 => to_unsigned(645, 12), 1716 => to_unsigned(1205, 12), 1717 => to_unsigned(278, 12), 1718 => to_unsigned(1525, 12), 1719 => to_unsigned(3694, 12), 1720 => to_unsigned(2082, 12), 1721 => to_unsigned(3131, 12), 1722 => to_unsigned(1313, 12), 1723 => to_unsigned(4092, 12), 1724 => to_unsigned(3895, 12), 1725 => to_unsigned(1334, 12), 1726 => to_unsigned(485, 12), 1727 => to_unsigned(1569, 12), 1728 => to_unsigned(3961, 12), 1729 => to_unsigned(3530, 12), 1730 => to_unsigned(1541, 12), 1731 => to_unsigned(1147, 12), 1732 => to_unsigned(479, 12), 1733 => to_unsigned(3892, 12), 1734 => to_unsigned(2166, 12), 1735 => to_unsigned(866, 12), 1736 => to_unsigned(2738, 12), 1737 => to_unsigned(2017, 12), 1738 => to_unsigned(1258, 12), 1739 => to_unsigned(187, 12), 1740 => to_unsigned(3483, 12), 1741 => to_unsigned(1028, 12), 1742 => to_unsigned(993, 12), 1743 => to_unsigned(3680, 12), 1744 => to_unsigned(1931, 12), 1745 => to_unsigned(1073, 12), 1746 => to_unsigned(1639, 12), 1747 => to_unsigned(505, 12), 1748 => to_unsigned(2027, 12), 1749 => to_unsigned(3941, 12), 1750 => to_unsigned(2047, 12), 1751 => to_unsigned(1771, 12), 1752 => to_unsigned(3339, 12), 1753 => to_unsigned(1572, 12), 1754 => to_unsigned(3776, 12), 1755 => to_unsigned(3943, 12), 1756 => to_unsigned(964, 12), 1757 => to_unsigned(641, 12), 1758 => to_unsigned(557, 12), 1759 => to_unsigned(3069, 12), 1760 => to_unsigned(152, 12), 1761 => to_unsigned(3749, 12), 1762 => to_unsigned(2904, 12), 1763 => to_unsigned(47, 12), 1764 => to_unsigned(277, 12), 1765 => to_unsigned(2104, 12), 1766 => to_unsigned(630, 12), 1767 => to_unsigned(2738, 12), 1768 => to_unsigned(3328, 12), 1769 => to_unsigned(664, 12), 1770 => to_unsigned(736, 12), 1771 => to_unsigned(4053, 12), 1772 => to_unsigned(1182, 12), 1773 => to_unsigned(210, 12), 1774 => to_unsigned(3643, 12), 1775 => to_unsigned(1135, 12), 1776 => to_unsigned(2748, 12), 1777 => to_unsigned(3985, 12), 1778 => to_unsigned(704, 12), 1779 => to_unsigned(402, 12), 1780 => to_unsigned(3060, 12), 1781 => to_unsigned(2746, 12), 1782 => to_unsigned(2381, 12), 1783 => to_unsigned(842, 12), 1784 => to_unsigned(3911, 12), 1785 => to_unsigned(1873, 12), 1786 => to_unsigned(2312, 12), 1787 => to_unsigned(554, 12), 1788 => to_unsigned(603, 12), 1789 => to_unsigned(1098, 12), 1790 => to_unsigned(958, 12), 1791 => to_unsigned(2096, 12), 1792 => to_unsigned(1576, 12), 1793 => to_unsigned(3613, 12), 1794 => to_unsigned(3819, 12), 1795 => to_unsigned(26, 12), 1796 => to_unsigned(3070, 12), 1797 => to_unsigned(3289, 12), 1798 => to_unsigned(3952, 12), 1799 => to_unsigned(822, 12), 1800 => to_unsigned(1739, 12), 1801 => to_unsigned(2341, 12), 1802 => to_unsigned(1690, 12), 1803 => to_unsigned(420, 12), 1804 => to_unsigned(2192, 12), 1805 => to_unsigned(1645, 12), 1806 => to_unsigned(200, 12), 1807 => to_unsigned(901, 12), 1808 => to_unsigned(1484, 12), 1809 => to_unsigned(1285, 12), 1810 => to_unsigned(1189, 12), 1811 => to_unsigned(515, 12), 1812 => to_unsigned(2426, 12), 1813 => to_unsigned(1935, 12), 1814 => to_unsigned(1975, 12), 1815 => to_unsigned(2403, 12), 1816 => to_unsigned(2410, 12), 1817 => to_unsigned(3917, 12), 1818 => to_unsigned(412, 12), 1819 => to_unsigned(1879, 12), 1820 => to_unsigned(3637, 12), 1821 => to_unsigned(230, 12), 1822 => to_unsigned(1785, 12), 1823 => to_unsigned(2918, 12), 1824 => to_unsigned(3180, 12), 1825 => to_unsigned(1176, 12), 1826 => to_unsigned(1207, 12), 1827 => to_unsigned(365, 12), 1828 => to_unsigned(3629, 12), 1829 => to_unsigned(3901, 12), 1830 => to_unsigned(1602, 12), 1831 => to_unsigned(3881, 12), 1832 => to_unsigned(1074, 12), 1833 => to_unsigned(1434, 12), 1834 => to_unsigned(2379, 12), 1835 => to_unsigned(42, 12), 1836 => to_unsigned(1793, 12), 1837 => to_unsigned(2661, 12), 1838 => to_unsigned(2137, 12), 1839 => to_unsigned(988, 12), 1840 => to_unsigned(3775, 12), 1841 => to_unsigned(556, 12), 1842 => to_unsigned(1208, 12), 1843 => to_unsigned(1885, 12), 1844 => to_unsigned(2853, 12), 1845 => to_unsigned(1128, 12), 1846 => to_unsigned(863, 12), 1847 => to_unsigned(741, 12), 1848 => to_unsigned(1845, 12), 1849 => to_unsigned(2772, 12), 1850 => to_unsigned(2623, 12), 1851 => to_unsigned(2119, 12), 1852 => to_unsigned(1029, 12), 1853 => to_unsigned(1475, 12), 1854 => to_unsigned(1296, 12), 1855 => to_unsigned(1556, 12), 1856 => to_unsigned(451, 12), 1857 => to_unsigned(1634, 12), 1858 => to_unsigned(2426, 12), 1859 => to_unsigned(3229, 12), 1860 => to_unsigned(1403, 12), 1861 => to_unsigned(2778, 12), 1862 => to_unsigned(843, 12), 1863 => to_unsigned(3759, 12), 1864 => to_unsigned(2939, 12), 1865 => to_unsigned(2067, 12), 1866 => to_unsigned(2023, 12), 1867 => to_unsigned(939, 12), 1868 => to_unsigned(1403, 12), 1869 => to_unsigned(168, 12), 1870 => to_unsigned(160, 12), 1871 => to_unsigned(4031, 12), 1872 => to_unsigned(2805, 12), 1873 => to_unsigned(137, 12), 1874 => to_unsigned(692, 12), 1875 => to_unsigned(2481, 12), 1876 => to_unsigned(2884, 12), 1877 => to_unsigned(2890, 12), 1878 => to_unsigned(4052, 12), 1879 => to_unsigned(2237, 12), 1880 => to_unsigned(3923, 12), 1881 => to_unsigned(1259, 12), 1882 => to_unsigned(4040, 12), 1883 => to_unsigned(1982, 12), 1884 => to_unsigned(1437, 12), 1885 => to_unsigned(2031, 12), 1886 => to_unsigned(179, 12), 1887 => to_unsigned(1091, 12), 1888 => to_unsigned(3764, 12), 1889 => to_unsigned(776, 12), 1890 => to_unsigned(3315, 12), 1891 => to_unsigned(1703, 12), 1892 => to_unsigned(315, 12), 1893 => to_unsigned(893, 12), 1894 => to_unsigned(578, 12), 1895 => to_unsigned(59, 12), 1896 => to_unsigned(1125, 12), 1897 => to_unsigned(3480, 12), 1898 => to_unsigned(1380, 12), 1899 => to_unsigned(29, 12), 1900 => to_unsigned(2398, 12), 1901 => to_unsigned(2384, 12), 1902 => to_unsigned(1673, 12), 1903 => to_unsigned(2439, 12), 1904 => to_unsigned(1593, 12), 1905 => to_unsigned(497, 12), 1906 => to_unsigned(3969, 12), 1907 => to_unsigned(223, 12), 1908 => to_unsigned(522, 12), 1909 => to_unsigned(2441, 12), 1910 => to_unsigned(168, 12), 1911 => to_unsigned(31, 12), 1912 => to_unsigned(855, 12), 1913 => to_unsigned(2182, 12), 1914 => to_unsigned(3963, 12), 1915 => to_unsigned(860, 12), 1916 => to_unsigned(1785, 12), 1917 => to_unsigned(2689, 12), 1918 => to_unsigned(2063, 12), 1919 => to_unsigned(3934, 12), 1920 => to_unsigned(3851, 12), 1921 => to_unsigned(2164, 12), 1922 => to_unsigned(956, 12), 1923 => to_unsigned(1247, 12), 1924 => to_unsigned(1582, 12), 1925 => to_unsigned(693, 12), 1926 => to_unsigned(1256, 12), 1927 => to_unsigned(2641, 12), 1928 => to_unsigned(1346, 12), 1929 => to_unsigned(3983, 12), 1930 => to_unsigned(2096, 12), 1931 => to_unsigned(2537, 12), 1932 => to_unsigned(3025, 12), 1933 => to_unsigned(2802, 12), 1934 => to_unsigned(1195, 12), 1935 => to_unsigned(2941, 12), 1936 => to_unsigned(3764, 12), 1937 => to_unsigned(3982, 12), 1938 => to_unsigned(552, 12), 1939 => to_unsigned(1723, 12), 1940 => to_unsigned(3556, 12), 1941 => to_unsigned(2134, 12), 1942 => to_unsigned(1597, 12), 1943 => to_unsigned(2457, 12), 1944 => to_unsigned(1094, 12), 1945 => to_unsigned(4022, 12), 1946 => to_unsigned(495, 12), 1947 => to_unsigned(823, 12), 1948 => to_unsigned(2161, 12), 1949 => to_unsigned(3220, 12), 1950 => to_unsigned(1756, 12), 1951 => to_unsigned(3948, 12), 1952 => to_unsigned(3590, 12), 1953 => to_unsigned(517, 12), 1954 => to_unsigned(1562, 12), 1955 => to_unsigned(1962, 12), 1956 => to_unsigned(2029, 12), 1957 => to_unsigned(1594, 12), 1958 => to_unsigned(1521, 12), 1959 => to_unsigned(754, 12), 1960 => to_unsigned(3728, 12), 1961 => to_unsigned(2391, 12), 1962 => to_unsigned(3611, 12), 1963 => to_unsigned(3193, 12), 1964 => to_unsigned(2585, 12), 1965 => to_unsigned(1701, 12), 1966 => to_unsigned(3289, 12), 1967 => to_unsigned(314, 12), 1968 => to_unsigned(3698, 12), 1969 => to_unsigned(758, 12), 1970 => to_unsigned(871, 12), 1971 => to_unsigned(1216, 12), 1972 => to_unsigned(338, 12), 1973 => to_unsigned(3033, 12), 1974 => to_unsigned(3298, 12), 1975 => to_unsigned(2895, 12), 1976 => to_unsigned(1804, 12), 1977 => to_unsigned(1545, 12), 1978 => to_unsigned(3911, 12), 1979 => to_unsigned(2522, 12), 1980 => to_unsigned(3481, 12), 1981 => to_unsigned(258, 12), 1982 => to_unsigned(3948, 12), 1983 => to_unsigned(2035, 12), 1984 => to_unsigned(2045, 12), 1985 => to_unsigned(2232, 12), 1986 => to_unsigned(867, 12), 1987 => to_unsigned(1576, 12), 1988 => to_unsigned(1991, 12), 1989 => to_unsigned(1567, 12), 1990 => to_unsigned(2514, 12), 1991 => to_unsigned(3019, 12), 1992 => to_unsigned(1019, 12), 1993 => to_unsigned(2943, 12), 1994 => to_unsigned(2988, 12), 1995 => to_unsigned(1407, 12), 1996 => to_unsigned(172, 12), 1997 => to_unsigned(1100, 12), 1998 => to_unsigned(1579, 12), 1999 => to_unsigned(2415, 12), 2000 => to_unsigned(1260, 12), 2001 => to_unsigned(2554, 12), 2002 => to_unsigned(2482, 12), 2003 => to_unsigned(1478, 12), 2004 => to_unsigned(46, 12), 2005 => to_unsigned(3950, 12), 2006 => to_unsigned(4047, 12), 2007 => to_unsigned(607, 12), 2008 => to_unsigned(1480, 12), 2009 => to_unsigned(3097, 12), 2010 => to_unsigned(1391, 12), 2011 => to_unsigned(1908, 12), 2012 => to_unsigned(3196, 12), 2013 => to_unsigned(1831, 12), 2014 => to_unsigned(1198, 12), 2015 => to_unsigned(2835, 12), 2016 => to_unsigned(4037, 12), 2017 => to_unsigned(1738, 12), 2018 => to_unsigned(220, 12), 2019 => to_unsigned(1094, 12), 2020 => to_unsigned(2780, 12), 2021 => to_unsigned(1657, 12), 2022 => to_unsigned(42, 12), 2023 => to_unsigned(3907, 12), 2024 => to_unsigned(314, 12), 2025 => to_unsigned(599, 12), 2026 => to_unsigned(706, 12), 2027 => to_unsigned(1483, 12), 2028 => to_unsigned(674, 12), 2029 => to_unsigned(2229, 12), 2030 => to_unsigned(1223, 12), 2031 => to_unsigned(2469, 12), 2032 => to_unsigned(3900, 12), 2033 => to_unsigned(3560, 12), 2034 => to_unsigned(3045, 12), 2035 => to_unsigned(3000, 12), 2036 => to_unsigned(462, 12), 2037 => to_unsigned(196, 12), 2038 => to_unsigned(3640, 12), 2039 => to_unsigned(2983, 12), 2040 => to_unsigned(760, 12), 2041 => to_unsigned(124, 12), 2042 => to_unsigned(2511, 12), 2043 => to_unsigned(958, 12), 2044 => to_unsigned(2349, 12), 2045 => to_unsigned(539, 12), 2046 => to_unsigned(2316, 12), 2047 => to_unsigned(360, 12)),
            4 => (0 => to_unsigned(3274, 12), 1 => to_unsigned(2212, 12), 2 => to_unsigned(635, 12), 3 => to_unsigned(834, 12), 4 => to_unsigned(135, 12), 5 => to_unsigned(1765, 12), 6 => to_unsigned(1326, 12), 7 => to_unsigned(417, 12), 8 => to_unsigned(1317, 12), 9 => to_unsigned(745, 12), 10 => to_unsigned(535, 12), 11 => to_unsigned(849, 12), 12 => to_unsigned(1688, 12), 13 => to_unsigned(2745, 12), 14 => to_unsigned(1209, 12), 15 => to_unsigned(2356, 12), 16 => to_unsigned(1329, 12), 17 => to_unsigned(2380, 12), 18 => to_unsigned(3686, 12), 19 => to_unsigned(4053, 12), 20 => to_unsigned(3421, 12), 21 => to_unsigned(1181, 12), 22 => to_unsigned(3641, 12), 23 => to_unsigned(740, 12), 24 => to_unsigned(1068, 12), 25 => to_unsigned(1194, 12), 26 => to_unsigned(2894, 12), 27 => to_unsigned(3298, 12), 28 => to_unsigned(2430, 12), 29 => to_unsigned(837, 12), 30 => to_unsigned(2314, 12), 31 => to_unsigned(1819, 12), 32 => to_unsigned(477, 12), 33 => to_unsigned(3215, 12), 34 => to_unsigned(1755, 12), 35 => to_unsigned(2072, 12), 36 => to_unsigned(1199, 12), 37 => to_unsigned(3421, 12), 38 => to_unsigned(693, 12), 39 => to_unsigned(3052, 12), 40 => to_unsigned(2957, 12), 41 => to_unsigned(1882, 12), 42 => to_unsigned(1711, 12), 43 => to_unsigned(4017, 12), 44 => to_unsigned(3101, 12), 45 => to_unsigned(1916, 12), 46 => to_unsigned(1929, 12), 47 => to_unsigned(3577, 12), 48 => to_unsigned(3155, 12), 49 => to_unsigned(2475, 12), 50 => to_unsigned(3782, 12), 51 => to_unsigned(1458, 12), 52 => to_unsigned(1569, 12), 53 => to_unsigned(1075, 12), 54 => to_unsigned(2202, 12), 55 => to_unsigned(3414, 12), 56 => to_unsigned(949, 12), 57 => to_unsigned(45, 12), 58 => to_unsigned(2156, 12), 59 => to_unsigned(3800, 12), 60 => to_unsigned(3163, 12), 61 => to_unsigned(2001, 12), 62 => to_unsigned(2956, 12), 63 => to_unsigned(1676, 12), 64 => to_unsigned(748, 12), 65 => to_unsigned(673, 12), 66 => to_unsigned(1229, 12), 67 => to_unsigned(923, 12), 68 => to_unsigned(2316, 12), 69 => to_unsigned(865, 12), 70 => to_unsigned(3652, 12), 71 => to_unsigned(743, 12), 72 => to_unsigned(1993, 12), 73 => to_unsigned(3427, 12), 74 => to_unsigned(1157, 12), 75 => to_unsigned(3058, 12), 76 => to_unsigned(3156, 12), 77 => to_unsigned(866, 12), 78 => to_unsigned(3855, 12), 79 => to_unsigned(2175, 12), 80 => to_unsigned(1555, 12), 81 => to_unsigned(2877, 12), 82 => to_unsigned(670, 12), 83 => to_unsigned(1988, 12), 84 => to_unsigned(1157, 12), 85 => to_unsigned(1729, 12), 86 => to_unsigned(2854, 12), 87 => to_unsigned(213, 12), 88 => to_unsigned(1354, 12), 89 => to_unsigned(1102, 12), 90 => to_unsigned(51, 12), 91 => to_unsigned(1740, 12), 92 => to_unsigned(2336, 12), 93 => to_unsigned(3324, 12), 94 => to_unsigned(3373, 12), 95 => to_unsigned(2061, 12), 96 => to_unsigned(486, 12), 97 => to_unsigned(3905, 12), 98 => to_unsigned(3574, 12), 99 => to_unsigned(265, 12), 100 => to_unsigned(3250, 12), 101 => to_unsigned(1257, 12), 102 => to_unsigned(1181, 12), 103 => to_unsigned(2783, 12), 104 => to_unsigned(4040, 12), 105 => to_unsigned(47, 12), 106 => to_unsigned(2063, 12), 107 => to_unsigned(2086, 12), 108 => to_unsigned(132, 12), 109 => to_unsigned(3885, 12), 110 => to_unsigned(3278, 12), 111 => to_unsigned(1795, 12), 112 => to_unsigned(2263, 12), 113 => to_unsigned(3004, 12), 114 => to_unsigned(856, 12), 115 => to_unsigned(1764, 12), 116 => to_unsigned(1431, 12), 117 => to_unsigned(3753, 12), 118 => to_unsigned(1804, 12), 119 => to_unsigned(531, 12), 120 => to_unsigned(1284, 12), 121 => to_unsigned(3506, 12), 122 => to_unsigned(2292, 12), 123 => to_unsigned(2515, 12), 124 => to_unsigned(913, 12), 125 => to_unsigned(3302, 12), 126 => to_unsigned(304, 12), 127 => to_unsigned(2242, 12), 128 => to_unsigned(2290, 12), 129 => to_unsigned(1963, 12), 130 => to_unsigned(1630, 12), 131 => to_unsigned(4061, 12), 132 => to_unsigned(3176, 12), 133 => to_unsigned(2583, 12), 134 => to_unsigned(3256, 12), 135 => to_unsigned(318, 12), 136 => to_unsigned(2934, 12), 137 => to_unsigned(3396, 12), 138 => to_unsigned(3283, 12), 139 => to_unsigned(1783, 12), 140 => to_unsigned(1047, 12), 141 => to_unsigned(400, 12), 142 => to_unsigned(3143, 12), 143 => to_unsigned(1556, 12), 144 => to_unsigned(973, 12), 145 => to_unsigned(1782, 12), 146 => to_unsigned(1265, 12), 147 => to_unsigned(2533, 12), 148 => to_unsigned(2847, 12), 149 => to_unsigned(3747, 12), 150 => to_unsigned(3131, 12), 151 => to_unsigned(103, 12), 152 => to_unsigned(835, 12), 153 => to_unsigned(2424, 12), 154 => to_unsigned(3284, 12), 155 => to_unsigned(792, 12), 156 => to_unsigned(2412, 12), 157 => to_unsigned(960, 12), 158 => to_unsigned(2862, 12), 159 => to_unsigned(1676, 12), 160 => to_unsigned(1679, 12), 161 => to_unsigned(1500, 12), 162 => to_unsigned(2470, 12), 163 => to_unsigned(3325, 12), 164 => to_unsigned(1628, 12), 165 => to_unsigned(1547, 12), 166 => to_unsigned(542, 12), 167 => to_unsigned(3411, 12), 168 => to_unsigned(3644, 12), 169 => to_unsigned(3810, 12), 170 => to_unsigned(1512, 12), 171 => to_unsigned(2523, 12), 172 => to_unsigned(2658, 12), 173 => to_unsigned(2232, 12), 174 => to_unsigned(860, 12), 175 => to_unsigned(3947, 12), 176 => to_unsigned(3750, 12), 177 => to_unsigned(2652, 12), 178 => to_unsigned(1505, 12), 179 => to_unsigned(1865, 12), 180 => to_unsigned(3172, 12), 181 => to_unsigned(3887, 12), 182 => to_unsigned(4019, 12), 183 => to_unsigned(3846, 12), 184 => to_unsigned(392, 12), 185 => to_unsigned(2319, 12), 186 => to_unsigned(1271, 12), 187 => to_unsigned(2964, 12), 188 => to_unsigned(845, 12), 189 => to_unsigned(3969, 12), 190 => to_unsigned(1654, 12), 191 => to_unsigned(3633, 12), 192 => to_unsigned(2649, 12), 193 => to_unsigned(1633, 12), 194 => to_unsigned(2222, 12), 195 => to_unsigned(304, 12), 196 => to_unsigned(3281, 12), 197 => to_unsigned(1995, 12), 198 => to_unsigned(1329, 12), 199 => to_unsigned(466, 12), 200 => to_unsigned(227, 12), 201 => to_unsigned(2789, 12), 202 => to_unsigned(3599, 12), 203 => to_unsigned(2221, 12), 204 => to_unsigned(391, 12), 205 => to_unsigned(72, 12), 206 => to_unsigned(195, 12), 207 => to_unsigned(1187, 12), 208 => to_unsigned(3446, 12), 209 => to_unsigned(366, 12), 210 => to_unsigned(613, 12), 211 => to_unsigned(1853, 12), 212 => to_unsigned(2608, 12), 213 => to_unsigned(624, 12), 214 => to_unsigned(2732, 12), 215 => to_unsigned(3827, 12), 216 => to_unsigned(707, 12), 217 => to_unsigned(3783, 12), 218 => to_unsigned(106, 12), 219 => to_unsigned(3078, 12), 220 => to_unsigned(130, 12), 221 => to_unsigned(1591, 12), 222 => to_unsigned(2048, 12), 223 => to_unsigned(3843, 12), 224 => to_unsigned(703, 12), 225 => to_unsigned(1472, 12), 226 => to_unsigned(1389, 12), 227 => to_unsigned(489, 12), 228 => to_unsigned(3259, 12), 229 => to_unsigned(3641, 12), 230 => to_unsigned(2469, 12), 231 => to_unsigned(3428, 12), 232 => to_unsigned(1547, 12), 233 => to_unsigned(2409, 12), 234 => to_unsigned(1417, 12), 235 => to_unsigned(1966, 12), 236 => to_unsigned(629, 12), 237 => to_unsigned(1024, 12), 238 => to_unsigned(2049, 12), 239 => to_unsigned(3467, 12), 240 => to_unsigned(870, 12), 241 => to_unsigned(1519, 12), 242 => to_unsigned(3619, 12), 243 => to_unsigned(518, 12), 244 => to_unsigned(3259, 12), 245 => to_unsigned(2552, 12), 246 => to_unsigned(3813, 12), 247 => to_unsigned(3288, 12), 248 => to_unsigned(3138, 12), 249 => to_unsigned(2105, 12), 250 => to_unsigned(2330, 12), 251 => to_unsigned(2161, 12), 252 => to_unsigned(215, 12), 253 => to_unsigned(346, 12), 254 => to_unsigned(1413, 12), 255 => to_unsigned(2456, 12), 256 => to_unsigned(2423, 12), 257 => to_unsigned(3178, 12), 258 => to_unsigned(2014, 12), 259 => to_unsigned(427, 12), 260 => to_unsigned(3464, 12), 261 => to_unsigned(2680, 12), 262 => to_unsigned(2278, 12), 263 => to_unsigned(1783, 12), 264 => to_unsigned(2237, 12), 265 => to_unsigned(1436, 12), 266 => to_unsigned(2125, 12), 267 => to_unsigned(3939, 12), 268 => to_unsigned(3185, 12), 269 => to_unsigned(3292, 12), 270 => to_unsigned(106, 12), 271 => to_unsigned(552, 12), 272 => to_unsigned(677, 12), 273 => to_unsigned(597, 12), 274 => to_unsigned(3595, 12), 275 => to_unsigned(3367, 12), 276 => to_unsigned(944, 12), 277 => to_unsigned(1113, 12), 278 => to_unsigned(2285, 12), 279 => to_unsigned(1435, 12), 280 => to_unsigned(3924, 12), 281 => to_unsigned(1498, 12), 282 => to_unsigned(2272, 12), 283 => to_unsigned(1978, 12), 284 => to_unsigned(1756, 12), 285 => to_unsigned(4086, 12), 286 => to_unsigned(575, 12), 287 => to_unsigned(1559, 12), 288 => to_unsigned(31, 12), 289 => to_unsigned(1349, 12), 290 => to_unsigned(4027, 12), 291 => to_unsigned(3610, 12), 292 => to_unsigned(1999, 12), 293 => to_unsigned(2147, 12), 294 => to_unsigned(1198, 12), 295 => to_unsigned(3677, 12), 296 => to_unsigned(3278, 12), 297 => to_unsigned(1211, 12), 298 => to_unsigned(2439, 12), 299 => to_unsigned(1590, 12), 300 => to_unsigned(1438, 12), 301 => to_unsigned(3592, 12), 302 => to_unsigned(2537, 12), 303 => to_unsigned(3255, 12), 304 => to_unsigned(1556, 12), 305 => to_unsigned(678, 12), 306 => to_unsigned(2918, 12), 307 => to_unsigned(4024, 12), 308 => to_unsigned(42, 12), 309 => to_unsigned(467, 12), 310 => to_unsigned(1625, 12), 311 => to_unsigned(2789, 12), 312 => to_unsigned(1258, 12), 313 => to_unsigned(3064, 12), 314 => to_unsigned(1741, 12), 315 => to_unsigned(1459, 12), 316 => to_unsigned(691, 12), 317 => to_unsigned(1839, 12), 318 => to_unsigned(3752, 12), 319 => to_unsigned(3638, 12), 320 => to_unsigned(532, 12), 321 => to_unsigned(4020, 12), 322 => to_unsigned(884, 12), 323 => to_unsigned(274, 12), 324 => to_unsigned(1917, 12), 325 => to_unsigned(61, 12), 326 => to_unsigned(2957, 12), 327 => to_unsigned(3959, 12), 328 => to_unsigned(2312, 12), 329 => to_unsigned(2345, 12), 330 => to_unsigned(3321, 12), 331 => to_unsigned(67, 12), 332 => to_unsigned(319, 12), 333 => to_unsigned(3990, 12), 334 => to_unsigned(2133, 12), 335 => to_unsigned(1747, 12), 336 => to_unsigned(3346, 12), 337 => to_unsigned(3154, 12), 338 => to_unsigned(726, 12), 339 => to_unsigned(1310, 12), 340 => to_unsigned(3251, 12), 341 => to_unsigned(2941, 12), 342 => to_unsigned(3579, 12), 343 => to_unsigned(749, 12), 344 => to_unsigned(1148, 12), 345 => to_unsigned(3666, 12), 346 => to_unsigned(939, 12), 347 => to_unsigned(1619, 12), 348 => to_unsigned(2422, 12), 349 => to_unsigned(153, 12), 350 => to_unsigned(1861, 12), 351 => to_unsigned(1435, 12), 352 => to_unsigned(2344, 12), 353 => to_unsigned(1214, 12), 354 => to_unsigned(3189, 12), 355 => to_unsigned(2499, 12), 356 => to_unsigned(880, 12), 357 => to_unsigned(1131, 12), 358 => to_unsigned(3144, 12), 359 => to_unsigned(816, 12), 360 => to_unsigned(3597, 12), 361 => to_unsigned(2334, 12), 362 => to_unsigned(2366, 12), 363 => to_unsigned(2420, 12), 364 => to_unsigned(2716, 12), 365 => to_unsigned(3696, 12), 366 => to_unsigned(2069, 12), 367 => to_unsigned(3964, 12), 368 => to_unsigned(1015, 12), 369 => to_unsigned(1596, 12), 370 => to_unsigned(72, 12), 371 => to_unsigned(3135, 12), 372 => to_unsigned(2954, 12), 373 => to_unsigned(1662, 12), 374 => to_unsigned(152, 12), 375 => to_unsigned(2209, 12), 376 => to_unsigned(2661, 12), 377 => to_unsigned(1348, 12), 378 => to_unsigned(686, 12), 379 => to_unsigned(1238, 12), 380 => to_unsigned(533, 12), 381 => to_unsigned(164, 12), 382 => to_unsigned(42, 12), 383 => to_unsigned(2926, 12), 384 => to_unsigned(70, 12), 385 => to_unsigned(839, 12), 386 => to_unsigned(2614, 12), 387 => to_unsigned(1738, 12), 388 => to_unsigned(2600, 12), 389 => to_unsigned(865, 12), 390 => to_unsigned(1307, 12), 391 => to_unsigned(2826, 12), 392 => to_unsigned(3449, 12), 393 => to_unsigned(2289, 12), 394 => to_unsigned(2046, 12), 395 => to_unsigned(2208, 12), 396 => to_unsigned(85, 12), 397 => to_unsigned(1625, 12), 398 => to_unsigned(3717, 12), 399 => to_unsigned(2629, 12), 400 => to_unsigned(466, 12), 401 => to_unsigned(2893, 12), 402 => to_unsigned(2274, 12), 403 => to_unsigned(1519, 12), 404 => to_unsigned(2094, 12), 405 => to_unsigned(3300, 12), 406 => to_unsigned(640, 12), 407 => to_unsigned(2455, 12), 408 => to_unsigned(1223, 12), 409 => to_unsigned(1464, 12), 410 => to_unsigned(1728, 12), 411 => to_unsigned(252, 12), 412 => to_unsigned(1936, 12), 413 => to_unsigned(2477, 12), 414 => to_unsigned(3811, 12), 415 => to_unsigned(874, 12), 416 => to_unsigned(4082, 12), 417 => to_unsigned(2113, 12), 418 => to_unsigned(2576, 12), 419 => to_unsigned(1800, 12), 420 => to_unsigned(3049, 12), 421 => to_unsigned(1148, 12), 422 => to_unsigned(3353, 12), 423 => to_unsigned(745, 12), 424 => to_unsigned(1413, 12), 425 => to_unsigned(389, 12), 426 => to_unsigned(3698, 12), 427 => to_unsigned(2128, 12), 428 => to_unsigned(547, 12), 429 => to_unsigned(955, 12), 430 => to_unsigned(716, 12), 431 => to_unsigned(3620, 12), 432 => to_unsigned(3688, 12), 433 => to_unsigned(2791, 12), 434 => to_unsigned(2237, 12), 435 => to_unsigned(3017, 12), 436 => to_unsigned(506, 12), 437 => to_unsigned(2114, 12), 438 => to_unsigned(413, 12), 439 => to_unsigned(1933, 12), 440 => to_unsigned(2328, 12), 441 => to_unsigned(2044, 12), 442 => to_unsigned(2035, 12), 443 => to_unsigned(2244, 12), 444 => to_unsigned(2365, 12), 445 => to_unsigned(2559, 12), 446 => to_unsigned(1362, 12), 447 => to_unsigned(3079, 12), 448 => to_unsigned(2868, 12), 449 => to_unsigned(61, 12), 450 => to_unsigned(2007, 12), 451 => to_unsigned(3109, 12), 452 => to_unsigned(147, 12), 453 => to_unsigned(3049, 12), 454 => to_unsigned(2560, 12), 455 => to_unsigned(646, 12), 456 => to_unsigned(1436, 12), 457 => to_unsigned(823, 12), 458 => to_unsigned(2300, 12), 459 => to_unsigned(1321, 12), 460 => to_unsigned(1256, 12), 461 => to_unsigned(383, 12), 462 => to_unsigned(2397, 12), 463 => to_unsigned(1951, 12), 464 => to_unsigned(431, 12), 465 => to_unsigned(77, 12), 466 => to_unsigned(1278, 12), 467 => to_unsigned(3800, 12), 468 => to_unsigned(4088, 12), 469 => to_unsigned(3281, 12), 470 => to_unsigned(3977, 12), 471 => to_unsigned(2965, 12), 472 => to_unsigned(3020, 12), 473 => to_unsigned(3679, 12), 474 => to_unsigned(1652, 12), 475 => to_unsigned(2882, 12), 476 => to_unsigned(3883, 12), 477 => to_unsigned(2705, 12), 478 => to_unsigned(480, 12), 479 => to_unsigned(3285, 12), 480 => to_unsigned(2652, 12), 481 => to_unsigned(3699, 12), 482 => to_unsigned(2794, 12), 483 => to_unsigned(2232, 12), 484 => to_unsigned(2051, 12), 485 => to_unsigned(604, 12), 486 => to_unsigned(2705, 12), 487 => to_unsigned(2176, 12), 488 => to_unsigned(1543, 12), 489 => to_unsigned(3614, 12), 490 => to_unsigned(1518, 12), 491 => to_unsigned(2665, 12), 492 => to_unsigned(3796, 12), 493 => to_unsigned(3173, 12), 494 => to_unsigned(1736, 12), 495 => to_unsigned(1648, 12), 496 => to_unsigned(3372, 12), 497 => to_unsigned(3923, 12), 498 => to_unsigned(1494, 12), 499 => to_unsigned(3463, 12), 500 => to_unsigned(2121, 12), 501 => to_unsigned(1580, 12), 502 => to_unsigned(2579, 12), 503 => to_unsigned(963, 12), 504 => to_unsigned(918, 12), 505 => to_unsigned(2784, 12), 506 => to_unsigned(3249, 12), 507 => to_unsigned(2305, 12), 508 => to_unsigned(1957, 12), 509 => to_unsigned(529, 12), 510 => to_unsigned(183, 12), 511 => to_unsigned(3916, 12), 512 => to_unsigned(817, 12), 513 => to_unsigned(3722, 12), 514 => to_unsigned(3640, 12), 515 => to_unsigned(1811, 12), 516 => to_unsigned(1153, 12), 517 => to_unsigned(2227, 12), 518 => to_unsigned(2988, 12), 519 => to_unsigned(1804, 12), 520 => to_unsigned(1999, 12), 521 => to_unsigned(2546, 12), 522 => to_unsigned(3094, 12), 523 => to_unsigned(1082, 12), 524 => to_unsigned(237, 12), 525 => to_unsigned(1458, 12), 526 => to_unsigned(475, 12), 527 => to_unsigned(2228, 12), 528 => to_unsigned(2188, 12), 529 => to_unsigned(25, 12), 530 => to_unsigned(3685, 12), 531 => to_unsigned(2819, 12), 532 => to_unsigned(3584, 12), 533 => to_unsigned(1533, 12), 534 => to_unsigned(1492, 12), 535 => to_unsigned(280, 12), 536 => to_unsigned(3448, 12), 537 => to_unsigned(2802, 12), 538 => to_unsigned(3511, 12), 539 => to_unsigned(2701, 12), 540 => to_unsigned(1842, 12), 541 => to_unsigned(1843, 12), 542 => to_unsigned(1946, 12), 543 => to_unsigned(3302, 12), 544 => to_unsigned(1918, 12), 545 => to_unsigned(1088, 12), 546 => to_unsigned(1142, 12), 547 => to_unsigned(346, 12), 548 => to_unsigned(1120, 12), 549 => to_unsigned(3968, 12), 550 => to_unsigned(1540, 12), 551 => to_unsigned(2724, 12), 552 => to_unsigned(829, 12), 553 => to_unsigned(609, 12), 554 => to_unsigned(102, 12), 555 => to_unsigned(132, 12), 556 => to_unsigned(3507, 12), 557 => to_unsigned(2833, 12), 558 => to_unsigned(3552, 12), 559 => to_unsigned(2250, 12), 560 => to_unsigned(547, 12), 561 => to_unsigned(2099, 12), 562 => to_unsigned(3071, 12), 563 => to_unsigned(4029, 12), 564 => to_unsigned(59, 12), 565 => to_unsigned(1189, 12), 566 => to_unsigned(3124, 12), 567 => to_unsigned(164, 12), 568 => to_unsigned(3286, 12), 569 => to_unsigned(789, 12), 570 => to_unsigned(1240, 12), 571 => to_unsigned(2988, 12), 572 => to_unsigned(2096, 12), 573 => to_unsigned(2813, 12), 574 => to_unsigned(2892, 12), 575 => to_unsigned(3554, 12), 576 => to_unsigned(179, 12), 577 => to_unsigned(508, 12), 578 => to_unsigned(2492, 12), 579 => to_unsigned(1197, 12), 580 => to_unsigned(2283, 12), 581 => to_unsigned(179, 12), 582 => to_unsigned(3174, 12), 583 => to_unsigned(2497, 12), 584 => to_unsigned(1844, 12), 585 => to_unsigned(3536, 12), 586 => to_unsigned(800, 12), 587 => to_unsigned(1106, 12), 588 => to_unsigned(3103, 12), 589 => to_unsigned(616, 12), 590 => to_unsigned(3253, 12), 591 => to_unsigned(346, 12), 592 => to_unsigned(183, 12), 593 => to_unsigned(1934, 12), 594 => to_unsigned(1911, 12), 595 => to_unsigned(1372, 12), 596 => to_unsigned(2098, 12), 597 => to_unsigned(1952, 12), 598 => to_unsigned(451, 12), 599 => to_unsigned(3563, 12), 600 => to_unsigned(1586, 12), 601 => to_unsigned(516, 12), 602 => to_unsigned(2423, 12), 603 => to_unsigned(2240, 12), 604 => to_unsigned(54, 12), 605 => to_unsigned(2258, 12), 606 => to_unsigned(3782, 12), 607 => to_unsigned(2683, 12), 608 => to_unsigned(2810, 12), 609 => to_unsigned(3810, 12), 610 => to_unsigned(2123, 12), 611 => to_unsigned(219, 12), 612 => to_unsigned(2959, 12), 613 => to_unsigned(1537, 12), 614 => to_unsigned(2916, 12), 615 => to_unsigned(1655, 12), 616 => to_unsigned(993, 12), 617 => to_unsigned(3241, 12), 618 => to_unsigned(3857, 12), 619 => to_unsigned(3829, 12), 620 => to_unsigned(2244, 12), 621 => to_unsigned(456, 12), 622 => to_unsigned(3731, 12), 623 => to_unsigned(1859, 12), 624 => to_unsigned(2512, 12), 625 => to_unsigned(931, 12), 626 => to_unsigned(2440, 12), 627 => to_unsigned(906, 12), 628 => to_unsigned(3618, 12), 629 => to_unsigned(1954, 12), 630 => to_unsigned(3762, 12), 631 => to_unsigned(3294, 12), 632 => to_unsigned(2526, 12), 633 => to_unsigned(278, 12), 634 => to_unsigned(1089, 12), 635 => to_unsigned(2185, 12), 636 => to_unsigned(554, 12), 637 => to_unsigned(1297, 12), 638 => to_unsigned(705, 12), 639 => to_unsigned(3960, 12), 640 => to_unsigned(2902, 12), 641 => to_unsigned(2797, 12), 642 => to_unsigned(2440, 12), 643 => to_unsigned(20, 12), 644 => to_unsigned(190, 12), 645 => to_unsigned(1421, 12), 646 => to_unsigned(1184, 12), 647 => to_unsigned(1123, 12), 648 => to_unsigned(1705, 12), 649 => to_unsigned(2253, 12), 650 => to_unsigned(3826, 12), 651 => to_unsigned(3751, 12), 652 => to_unsigned(175, 12), 653 => to_unsigned(3531, 12), 654 => to_unsigned(2966, 12), 655 => to_unsigned(2093, 12), 656 => to_unsigned(2543, 12), 657 => to_unsigned(2985, 12), 658 => to_unsigned(1080, 12), 659 => to_unsigned(3513, 12), 660 => to_unsigned(2096, 12), 661 => to_unsigned(1761, 12), 662 => to_unsigned(3023, 12), 663 => to_unsigned(2573, 12), 664 => to_unsigned(3600, 12), 665 => to_unsigned(1763, 12), 666 => to_unsigned(2415, 12), 667 => to_unsigned(2363, 12), 668 => to_unsigned(886, 12), 669 => to_unsigned(889, 12), 670 => to_unsigned(2059, 12), 671 => to_unsigned(3678, 12), 672 => to_unsigned(3989, 12), 673 => to_unsigned(2020, 12), 674 => to_unsigned(1767, 12), 675 => to_unsigned(1869, 12), 676 => to_unsigned(2182, 12), 677 => to_unsigned(2971, 12), 678 => to_unsigned(1554, 12), 679 => to_unsigned(813, 12), 680 => to_unsigned(977, 12), 681 => to_unsigned(4029, 12), 682 => to_unsigned(2207, 12), 683 => to_unsigned(3930, 12), 684 => to_unsigned(1045, 12), 685 => to_unsigned(3679, 12), 686 => to_unsigned(1608, 12), 687 => to_unsigned(1963, 12), 688 => to_unsigned(1413, 12), 689 => to_unsigned(3141, 12), 690 => to_unsigned(272, 12), 691 => to_unsigned(1792, 12), 692 => to_unsigned(3031, 12), 693 => to_unsigned(4033, 12), 694 => to_unsigned(3384, 12), 695 => to_unsigned(1701, 12), 696 => to_unsigned(3382, 12), 697 => to_unsigned(967, 12), 698 => to_unsigned(3005, 12), 699 => to_unsigned(3659, 12), 700 => to_unsigned(1507, 12), 701 => to_unsigned(3693, 12), 702 => to_unsigned(932, 12), 703 => to_unsigned(2013, 12), 704 => to_unsigned(851, 12), 705 => to_unsigned(3625, 12), 706 => to_unsigned(698, 12), 707 => to_unsigned(1611, 12), 708 => to_unsigned(1927, 12), 709 => to_unsigned(142, 12), 710 => to_unsigned(1179, 12), 711 => to_unsigned(2098, 12), 712 => to_unsigned(1637, 12), 713 => to_unsigned(2373, 12), 714 => to_unsigned(776, 12), 715 => to_unsigned(1460, 12), 716 => to_unsigned(1348, 12), 717 => to_unsigned(46, 12), 718 => to_unsigned(2256, 12), 719 => to_unsigned(2253, 12), 720 => to_unsigned(3798, 12), 721 => to_unsigned(1721, 12), 722 => to_unsigned(1962, 12), 723 => to_unsigned(3282, 12), 724 => to_unsigned(785, 12), 725 => to_unsigned(893, 12), 726 => to_unsigned(2793, 12), 727 => to_unsigned(1923, 12), 728 => to_unsigned(1237, 12), 729 => to_unsigned(2808, 12), 730 => to_unsigned(1103, 12), 731 => to_unsigned(3628, 12), 732 => to_unsigned(3260, 12), 733 => to_unsigned(3021, 12), 734 => to_unsigned(1043, 12), 735 => to_unsigned(1881, 12), 736 => to_unsigned(1412, 12), 737 => to_unsigned(7, 12), 738 => to_unsigned(1383, 12), 739 => to_unsigned(981, 12), 740 => to_unsigned(2194, 12), 741 => to_unsigned(1397, 12), 742 => to_unsigned(1343, 12), 743 => to_unsigned(2403, 12), 744 => to_unsigned(3679, 12), 745 => to_unsigned(244, 12), 746 => to_unsigned(1433, 12), 747 => to_unsigned(2080, 12), 748 => to_unsigned(2257, 12), 749 => to_unsigned(1485, 12), 750 => to_unsigned(2813, 12), 751 => to_unsigned(3191, 12), 752 => to_unsigned(1143, 12), 753 => to_unsigned(499, 12), 754 => to_unsigned(3099, 12), 755 => to_unsigned(3061, 12), 756 => to_unsigned(336, 12), 757 => to_unsigned(3932, 12), 758 => to_unsigned(2350, 12), 759 => to_unsigned(1791, 12), 760 => to_unsigned(2706, 12), 761 => to_unsigned(2914, 12), 762 => to_unsigned(2999, 12), 763 => to_unsigned(64, 12), 764 => to_unsigned(283, 12), 765 => to_unsigned(3867, 12), 766 => to_unsigned(2843, 12), 767 => to_unsigned(32, 12), 768 => to_unsigned(1450, 12), 769 => to_unsigned(3602, 12), 770 => to_unsigned(3412, 12), 771 => to_unsigned(1393, 12), 772 => to_unsigned(2058, 12), 773 => to_unsigned(3067, 12), 774 => to_unsigned(1715, 12), 775 => to_unsigned(3656, 12), 776 => to_unsigned(44, 12), 777 => to_unsigned(2127, 12), 778 => to_unsigned(1314, 12), 779 => to_unsigned(3307, 12), 780 => to_unsigned(3192, 12), 781 => to_unsigned(3010, 12), 782 => to_unsigned(2209, 12), 783 => to_unsigned(1222, 12), 784 => to_unsigned(1183, 12), 785 => to_unsigned(3621, 12), 786 => to_unsigned(1281, 12), 787 => to_unsigned(2956, 12), 788 => to_unsigned(732, 12), 789 => to_unsigned(2296, 12), 790 => to_unsigned(1012, 12), 791 => to_unsigned(1117, 12), 792 => to_unsigned(3443, 12), 793 => to_unsigned(1957, 12), 794 => to_unsigned(4092, 12), 795 => to_unsigned(1646, 12), 796 => to_unsigned(2613, 12), 797 => to_unsigned(2320, 12), 798 => to_unsigned(2360, 12), 799 => to_unsigned(1023, 12), 800 => to_unsigned(835, 12), 801 => to_unsigned(1620, 12), 802 => to_unsigned(2490, 12), 803 => to_unsigned(498, 12), 804 => to_unsigned(201, 12), 805 => to_unsigned(61, 12), 806 => to_unsigned(2181, 12), 807 => to_unsigned(855, 12), 808 => to_unsigned(3811, 12), 809 => to_unsigned(2045, 12), 810 => to_unsigned(3023, 12), 811 => to_unsigned(1251, 12), 812 => to_unsigned(1662, 12), 813 => to_unsigned(3199, 12), 814 => to_unsigned(728, 12), 815 => to_unsigned(657, 12), 816 => to_unsigned(14, 12), 817 => to_unsigned(2395, 12), 818 => to_unsigned(3322, 12), 819 => to_unsigned(1240, 12), 820 => to_unsigned(2285, 12), 821 => to_unsigned(972, 12), 822 => to_unsigned(2294, 12), 823 => to_unsigned(658, 12), 824 => to_unsigned(287, 12), 825 => to_unsigned(1790, 12), 826 => to_unsigned(113, 12), 827 => to_unsigned(2732, 12), 828 => to_unsigned(1907, 12), 829 => to_unsigned(56, 12), 830 => to_unsigned(1655, 12), 831 => to_unsigned(3094, 12), 832 => to_unsigned(2912, 12), 833 => to_unsigned(959, 12), 834 => to_unsigned(2062, 12), 835 => to_unsigned(1148, 12), 836 => to_unsigned(113, 12), 837 => to_unsigned(369, 12), 838 => to_unsigned(2035, 12), 839 => to_unsigned(1945, 12), 840 => to_unsigned(1828, 12), 841 => to_unsigned(3561, 12), 842 => to_unsigned(1853, 12), 843 => to_unsigned(960, 12), 844 => to_unsigned(2161, 12), 845 => to_unsigned(536, 12), 846 => to_unsigned(2085, 12), 847 => to_unsigned(3984, 12), 848 => to_unsigned(2607, 12), 849 => to_unsigned(526, 12), 850 => to_unsigned(2537, 12), 851 => to_unsigned(3169, 12), 852 => to_unsigned(1078, 12), 853 => to_unsigned(3196, 12), 854 => to_unsigned(3169, 12), 855 => to_unsigned(3780, 12), 856 => to_unsigned(3538, 12), 857 => to_unsigned(809, 12), 858 => to_unsigned(2464, 12), 859 => to_unsigned(2627, 12), 860 => to_unsigned(1395, 12), 861 => to_unsigned(3828, 12), 862 => to_unsigned(1409, 12), 863 => to_unsigned(3308, 12), 864 => to_unsigned(3565, 12), 865 => to_unsigned(2522, 12), 866 => to_unsigned(824, 12), 867 => to_unsigned(917, 12), 868 => to_unsigned(2811, 12), 869 => to_unsigned(2323, 12), 870 => to_unsigned(858, 12), 871 => to_unsigned(1415, 12), 872 => to_unsigned(1873, 12), 873 => to_unsigned(139, 12), 874 => to_unsigned(618, 12), 875 => to_unsigned(366, 12), 876 => to_unsigned(2049, 12), 877 => to_unsigned(687, 12), 878 => to_unsigned(3375, 12), 879 => to_unsigned(2315, 12), 880 => to_unsigned(1401, 12), 881 => to_unsigned(1722, 12), 882 => to_unsigned(2063, 12), 883 => to_unsigned(483, 12), 884 => to_unsigned(858, 12), 885 => to_unsigned(3199, 12), 886 => to_unsigned(1109, 12), 887 => to_unsigned(3491, 12), 888 => to_unsigned(1246, 12), 889 => to_unsigned(9, 12), 890 => to_unsigned(111, 12), 891 => to_unsigned(2036, 12), 892 => to_unsigned(3394, 12), 893 => to_unsigned(3832, 12), 894 => to_unsigned(1405, 12), 895 => to_unsigned(2538, 12), 896 => to_unsigned(3904, 12), 897 => to_unsigned(894, 12), 898 => to_unsigned(375, 12), 899 => to_unsigned(2570, 12), 900 => to_unsigned(2317, 12), 901 => to_unsigned(3341, 12), 902 => to_unsigned(3732, 12), 903 => to_unsigned(168, 12), 904 => to_unsigned(3744, 12), 905 => to_unsigned(79, 12), 906 => to_unsigned(3822, 12), 907 => to_unsigned(1441, 12), 908 => to_unsigned(1049, 12), 909 => to_unsigned(2549, 12), 910 => to_unsigned(3821, 12), 911 => to_unsigned(3327, 12), 912 => to_unsigned(889, 12), 913 => to_unsigned(3782, 12), 914 => to_unsigned(289, 12), 915 => to_unsigned(1510, 12), 916 => to_unsigned(1976, 12), 917 => to_unsigned(2715, 12), 918 => to_unsigned(3569, 12), 919 => to_unsigned(2895, 12), 920 => to_unsigned(2992, 12), 921 => to_unsigned(2411, 12), 922 => to_unsigned(3629, 12), 923 => to_unsigned(2114, 12), 924 => to_unsigned(667, 12), 925 => to_unsigned(184, 12), 926 => to_unsigned(3559, 12), 927 => to_unsigned(2657, 12), 928 => to_unsigned(1480, 12), 929 => to_unsigned(521, 12), 930 => to_unsigned(1571, 12), 931 => to_unsigned(2267, 12), 932 => to_unsigned(2738, 12), 933 => to_unsigned(1682, 12), 934 => to_unsigned(1730, 12), 935 => to_unsigned(3977, 12), 936 => to_unsigned(971, 12), 937 => to_unsigned(353, 12), 938 => to_unsigned(4009, 12), 939 => to_unsigned(162, 12), 940 => to_unsigned(1229, 12), 941 => to_unsigned(2085, 12), 942 => to_unsigned(590, 12), 943 => to_unsigned(3139, 12), 944 => to_unsigned(648, 12), 945 => to_unsigned(3396, 12), 946 => to_unsigned(3360, 12), 947 => to_unsigned(507, 12), 948 => to_unsigned(1446, 12), 949 => to_unsigned(739, 12), 950 => to_unsigned(1162, 12), 951 => to_unsigned(1939, 12), 952 => to_unsigned(990, 12), 953 => to_unsigned(927, 12), 954 => to_unsigned(1861, 12), 955 => to_unsigned(3216, 12), 956 => to_unsigned(3455, 12), 957 => to_unsigned(2892, 12), 958 => to_unsigned(3813, 12), 959 => to_unsigned(2647, 12), 960 => to_unsigned(2550, 12), 961 => to_unsigned(1636, 12), 962 => to_unsigned(2988, 12), 963 => to_unsigned(2964, 12), 964 => to_unsigned(2223, 12), 965 => to_unsigned(2889, 12), 966 => to_unsigned(2974, 12), 967 => to_unsigned(2603, 12), 968 => to_unsigned(3118, 12), 969 => to_unsigned(1862, 12), 970 => to_unsigned(115, 12), 971 => to_unsigned(1607, 12), 972 => to_unsigned(4027, 12), 973 => to_unsigned(113, 12), 974 => to_unsigned(993, 12), 975 => to_unsigned(495, 12), 976 => to_unsigned(3132, 12), 977 => to_unsigned(2740, 12), 978 => to_unsigned(3242, 12), 979 => to_unsigned(1268, 12), 980 => to_unsigned(2593, 12), 981 => to_unsigned(1092, 12), 982 => to_unsigned(2234, 12), 983 => to_unsigned(451, 12), 984 => to_unsigned(2452, 12), 985 => to_unsigned(2559, 12), 986 => to_unsigned(124, 12), 987 => to_unsigned(3559, 12), 988 => to_unsigned(3066, 12), 989 => to_unsigned(1276, 12), 990 => to_unsigned(1677, 12), 991 => to_unsigned(377, 12), 992 => to_unsigned(2751, 12), 993 => to_unsigned(2539, 12), 994 => to_unsigned(4005, 12), 995 => to_unsigned(1467, 12), 996 => to_unsigned(910, 12), 997 => to_unsigned(1827, 12), 998 => to_unsigned(440, 12), 999 => to_unsigned(2199, 12), 1000 => to_unsigned(3770, 12), 1001 => to_unsigned(2114, 12), 1002 => to_unsigned(1508, 12), 1003 => to_unsigned(1071, 12), 1004 => to_unsigned(933, 12), 1005 => to_unsigned(337, 12), 1006 => to_unsigned(3537, 12), 1007 => to_unsigned(2585, 12), 1008 => to_unsigned(722, 12), 1009 => to_unsigned(342, 12), 1010 => to_unsigned(841, 12), 1011 => to_unsigned(3762, 12), 1012 => to_unsigned(2941, 12), 1013 => to_unsigned(1068, 12), 1014 => to_unsigned(186, 12), 1015 => to_unsigned(3944, 12), 1016 => to_unsigned(16, 12), 1017 => to_unsigned(2073, 12), 1018 => to_unsigned(2309, 12), 1019 => to_unsigned(2787, 12), 1020 => to_unsigned(124, 12), 1021 => to_unsigned(3440, 12), 1022 => to_unsigned(839, 12), 1023 => to_unsigned(2021, 12), 1024 => to_unsigned(604, 12), 1025 => to_unsigned(1663, 12), 1026 => to_unsigned(1730, 12), 1027 => to_unsigned(2310, 12), 1028 => to_unsigned(1022, 12), 1029 => to_unsigned(150, 12), 1030 => to_unsigned(1256, 12), 1031 => to_unsigned(3056, 12), 1032 => to_unsigned(1024, 12), 1033 => to_unsigned(2721, 12), 1034 => to_unsigned(200, 12), 1035 => to_unsigned(4080, 12), 1036 => to_unsigned(1137, 12), 1037 => to_unsigned(329, 12), 1038 => to_unsigned(1190, 12), 1039 => to_unsigned(3105, 12), 1040 => to_unsigned(3825, 12), 1041 => to_unsigned(2975, 12), 1042 => to_unsigned(2160, 12), 1043 => to_unsigned(2381, 12), 1044 => to_unsigned(2406, 12), 1045 => to_unsigned(2128, 12), 1046 => to_unsigned(246, 12), 1047 => to_unsigned(1524, 12), 1048 => to_unsigned(2897, 12), 1049 => to_unsigned(1217, 12), 1050 => to_unsigned(2376, 12), 1051 => to_unsigned(2003, 12), 1052 => to_unsigned(951, 12), 1053 => to_unsigned(3187, 12), 1054 => to_unsigned(3343, 12), 1055 => to_unsigned(3070, 12), 1056 => to_unsigned(3168, 12), 1057 => to_unsigned(4011, 12), 1058 => to_unsigned(1420, 12), 1059 => to_unsigned(2381, 12), 1060 => to_unsigned(3949, 12), 1061 => to_unsigned(3545, 12), 1062 => to_unsigned(426, 12), 1063 => to_unsigned(1916, 12), 1064 => to_unsigned(2291, 12), 1065 => to_unsigned(1917, 12), 1066 => to_unsigned(644, 12), 1067 => to_unsigned(3397, 12), 1068 => to_unsigned(2528, 12), 1069 => to_unsigned(3533, 12), 1070 => to_unsigned(2240, 12), 1071 => to_unsigned(2169, 12), 1072 => to_unsigned(1952, 12), 1073 => to_unsigned(1952, 12), 1074 => to_unsigned(2839, 12), 1075 => to_unsigned(2883, 12), 1076 => to_unsigned(1804, 12), 1077 => to_unsigned(3466, 12), 1078 => to_unsigned(94, 12), 1079 => to_unsigned(1592, 12), 1080 => to_unsigned(2453, 12), 1081 => to_unsigned(938, 12), 1082 => to_unsigned(2549, 12), 1083 => to_unsigned(2173, 12), 1084 => to_unsigned(707, 12), 1085 => to_unsigned(1563, 12), 1086 => to_unsigned(1185, 12), 1087 => to_unsigned(3803, 12), 1088 => to_unsigned(421, 12), 1089 => to_unsigned(2411, 12), 1090 => to_unsigned(515, 12), 1091 => to_unsigned(1892, 12), 1092 => to_unsigned(793, 12), 1093 => to_unsigned(1634, 12), 1094 => to_unsigned(1336, 12), 1095 => to_unsigned(3008, 12), 1096 => to_unsigned(844, 12), 1097 => to_unsigned(1036, 12), 1098 => to_unsigned(2155, 12), 1099 => to_unsigned(2573, 12), 1100 => to_unsigned(259, 12), 1101 => to_unsigned(3277, 12), 1102 => to_unsigned(968, 12), 1103 => to_unsigned(1809, 12), 1104 => to_unsigned(3999, 12), 1105 => to_unsigned(1056, 12), 1106 => to_unsigned(1768, 12), 1107 => to_unsigned(3665, 12), 1108 => to_unsigned(1138, 12), 1109 => to_unsigned(2310, 12), 1110 => to_unsigned(4081, 12), 1111 => to_unsigned(3394, 12), 1112 => to_unsigned(802, 12), 1113 => to_unsigned(1612, 12), 1114 => to_unsigned(1489, 12), 1115 => to_unsigned(1559, 12), 1116 => to_unsigned(680, 12), 1117 => to_unsigned(3954, 12), 1118 => to_unsigned(3663, 12), 1119 => to_unsigned(162, 12), 1120 => to_unsigned(1827, 12), 1121 => to_unsigned(2012, 12), 1122 => to_unsigned(670, 12), 1123 => to_unsigned(3109, 12), 1124 => to_unsigned(1321, 12), 1125 => to_unsigned(3303, 12), 1126 => to_unsigned(3709, 12), 1127 => to_unsigned(2738, 12), 1128 => to_unsigned(2904, 12), 1129 => to_unsigned(2501, 12), 1130 => to_unsigned(2209, 12), 1131 => to_unsigned(2520, 12), 1132 => to_unsigned(215, 12), 1133 => to_unsigned(3689, 12), 1134 => to_unsigned(862, 12), 1135 => to_unsigned(1897, 12), 1136 => to_unsigned(3761, 12), 1137 => to_unsigned(4059, 12), 1138 => to_unsigned(2203, 12), 1139 => to_unsigned(1533, 12), 1140 => to_unsigned(3681, 12), 1141 => to_unsigned(1884, 12), 1142 => to_unsigned(1962, 12), 1143 => to_unsigned(2791, 12), 1144 => to_unsigned(1846, 12), 1145 => to_unsigned(3794, 12), 1146 => to_unsigned(3699, 12), 1147 => to_unsigned(1176, 12), 1148 => to_unsigned(1644, 12), 1149 => to_unsigned(4043, 12), 1150 => to_unsigned(3662, 12), 1151 => to_unsigned(1082, 12), 1152 => to_unsigned(4084, 12), 1153 => to_unsigned(2373, 12), 1154 => to_unsigned(1138, 12), 1155 => to_unsigned(1395, 12), 1156 => to_unsigned(2660, 12), 1157 => to_unsigned(1345, 12), 1158 => to_unsigned(1169, 12), 1159 => to_unsigned(3901, 12), 1160 => to_unsigned(1105, 12), 1161 => to_unsigned(3305, 12), 1162 => to_unsigned(3642, 12), 1163 => to_unsigned(1156, 12), 1164 => to_unsigned(992, 12), 1165 => to_unsigned(1975, 12), 1166 => to_unsigned(1979, 12), 1167 => to_unsigned(1388, 12), 1168 => to_unsigned(3665, 12), 1169 => to_unsigned(1571, 12), 1170 => to_unsigned(68, 12), 1171 => to_unsigned(2209, 12), 1172 => to_unsigned(7, 12), 1173 => to_unsigned(3596, 12), 1174 => to_unsigned(749, 12), 1175 => to_unsigned(1808, 12), 1176 => to_unsigned(1387, 12), 1177 => to_unsigned(754, 12), 1178 => to_unsigned(2661, 12), 1179 => to_unsigned(1234, 12), 1180 => to_unsigned(2457, 12), 1181 => to_unsigned(343, 12), 1182 => to_unsigned(3559, 12), 1183 => to_unsigned(19, 12), 1184 => to_unsigned(3158, 12), 1185 => to_unsigned(48, 12), 1186 => to_unsigned(3183, 12), 1187 => to_unsigned(988, 12), 1188 => to_unsigned(3566, 12), 1189 => to_unsigned(3408, 12), 1190 => to_unsigned(3574, 12), 1191 => to_unsigned(540, 12), 1192 => to_unsigned(3163, 12), 1193 => to_unsigned(96, 12), 1194 => to_unsigned(1918, 12), 1195 => to_unsigned(2148, 12), 1196 => to_unsigned(1063, 12), 1197 => to_unsigned(979, 12), 1198 => to_unsigned(193, 12), 1199 => to_unsigned(3449, 12), 1200 => to_unsigned(1501, 12), 1201 => to_unsigned(551, 12), 1202 => to_unsigned(3724, 12), 1203 => to_unsigned(1313, 12), 1204 => to_unsigned(3065, 12), 1205 => to_unsigned(2569, 12), 1206 => to_unsigned(3683, 12), 1207 => to_unsigned(1784, 12), 1208 => to_unsigned(807, 12), 1209 => to_unsigned(1861, 12), 1210 => to_unsigned(3469, 12), 1211 => to_unsigned(2123, 12), 1212 => to_unsigned(1625, 12), 1213 => to_unsigned(2795, 12), 1214 => to_unsigned(1845, 12), 1215 => to_unsigned(3745, 12), 1216 => to_unsigned(178, 12), 1217 => to_unsigned(3868, 12), 1218 => to_unsigned(3310, 12), 1219 => to_unsigned(1562, 12), 1220 => to_unsigned(207, 12), 1221 => to_unsigned(770, 12), 1222 => to_unsigned(1645, 12), 1223 => to_unsigned(2010, 12), 1224 => to_unsigned(2095, 12), 1225 => to_unsigned(1606, 12), 1226 => to_unsigned(1557, 12), 1227 => to_unsigned(1289, 12), 1228 => to_unsigned(1744, 12), 1229 => to_unsigned(1573, 12), 1230 => to_unsigned(757, 12), 1231 => to_unsigned(535, 12), 1232 => to_unsigned(493, 12), 1233 => to_unsigned(602, 12), 1234 => to_unsigned(3590, 12), 1235 => to_unsigned(3778, 12), 1236 => to_unsigned(3357, 12), 1237 => to_unsigned(2853, 12), 1238 => to_unsigned(2471, 12), 1239 => to_unsigned(1049, 12), 1240 => to_unsigned(619, 12), 1241 => to_unsigned(432, 12), 1242 => to_unsigned(3858, 12), 1243 => to_unsigned(2490, 12), 1244 => to_unsigned(592, 12), 1245 => to_unsigned(1970, 12), 1246 => to_unsigned(430, 12), 1247 => to_unsigned(2897, 12), 1248 => to_unsigned(749, 12), 1249 => to_unsigned(638, 12), 1250 => to_unsigned(2555, 12), 1251 => to_unsigned(400, 12), 1252 => to_unsigned(1304, 12), 1253 => to_unsigned(3884, 12), 1254 => to_unsigned(3212, 12), 1255 => to_unsigned(2217, 12), 1256 => to_unsigned(1748, 12), 1257 => to_unsigned(3130, 12), 1258 => to_unsigned(155, 12), 1259 => to_unsigned(1296, 12), 1260 => to_unsigned(2340, 12), 1261 => to_unsigned(1503, 12), 1262 => to_unsigned(3324, 12), 1263 => to_unsigned(2316, 12), 1264 => to_unsigned(3333, 12), 1265 => to_unsigned(3341, 12), 1266 => to_unsigned(2477, 12), 1267 => to_unsigned(3945, 12), 1268 => to_unsigned(1394, 12), 1269 => to_unsigned(994, 12), 1270 => to_unsigned(79, 12), 1271 => to_unsigned(1137, 12), 1272 => to_unsigned(293, 12), 1273 => to_unsigned(547, 12), 1274 => to_unsigned(3296, 12), 1275 => to_unsigned(104, 12), 1276 => to_unsigned(1023, 12), 1277 => to_unsigned(3849, 12), 1278 => to_unsigned(367, 12), 1279 => to_unsigned(2429, 12), 1280 => to_unsigned(2088, 12), 1281 => to_unsigned(3086, 12), 1282 => to_unsigned(2819, 12), 1283 => to_unsigned(2961, 12), 1284 => to_unsigned(1451, 12), 1285 => to_unsigned(710, 12), 1286 => to_unsigned(2007, 12), 1287 => to_unsigned(3354, 12), 1288 => to_unsigned(1324, 12), 1289 => to_unsigned(2972, 12), 1290 => to_unsigned(1253, 12), 1291 => to_unsigned(1916, 12), 1292 => to_unsigned(650, 12), 1293 => to_unsigned(3506, 12), 1294 => to_unsigned(253, 12), 1295 => to_unsigned(2578, 12), 1296 => to_unsigned(492, 12), 1297 => to_unsigned(723, 12), 1298 => to_unsigned(861, 12), 1299 => to_unsigned(2947, 12), 1300 => to_unsigned(2820, 12), 1301 => to_unsigned(687, 12), 1302 => to_unsigned(2734, 12), 1303 => to_unsigned(3919, 12), 1304 => to_unsigned(2000, 12), 1305 => to_unsigned(587, 12), 1306 => to_unsigned(2989, 12), 1307 => to_unsigned(3947, 12), 1308 => to_unsigned(2827, 12), 1309 => to_unsigned(3839, 12), 1310 => to_unsigned(639, 12), 1311 => to_unsigned(3228, 12), 1312 => to_unsigned(1026, 12), 1313 => to_unsigned(1061, 12), 1314 => to_unsigned(327, 12), 1315 => to_unsigned(1606, 12), 1316 => to_unsigned(3564, 12), 1317 => to_unsigned(15, 12), 1318 => to_unsigned(3675, 12), 1319 => to_unsigned(93, 12), 1320 => to_unsigned(3811, 12), 1321 => to_unsigned(1157, 12), 1322 => to_unsigned(516, 12), 1323 => to_unsigned(1580, 12), 1324 => to_unsigned(2022, 12), 1325 => to_unsigned(2130, 12), 1326 => to_unsigned(3833, 12), 1327 => to_unsigned(2269, 12), 1328 => to_unsigned(1294, 12), 1329 => to_unsigned(4008, 12), 1330 => to_unsigned(1114, 12), 1331 => to_unsigned(871, 12), 1332 => to_unsigned(3106, 12), 1333 => to_unsigned(2072, 12), 1334 => to_unsigned(2443, 12), 1335 => to_unsigned(2214, 12), 1336 => to_unsigned(2100, 12), 1337 => to_unsigned(2329, 12), 1338 => to_unsigned(692, 12), 1339 => to_unsigned(2606, 12), 1340 => to_unsigned(1464, 12), 1341 => to_unsigned(3049, 12), 1342 => to_unsigned(46, 12), 1343 => to_unsigned(3262, 12), 1344 => to_unsigned(1402, 12), 1345 => to_unsigned(958, 12), 1346 => to_unsigned(2390, 12), 1347 => to_unsigned(2984, 12), 1348 => to_unsigned(2771, 12), 1349 => to_unsigned(4089, 12), 1350 => to_unsigned(2940, 12), 1351 => to_unsigned(1871, 12), 1352 => to_unsigned(1926, 12), 1353 => to_unsigned(2176, 12), 1354 => to_unsigned(2938, 12), 1355 => to_unsigned(743, 12), 1356 => to_unsigned(3937, 12), 1357 => to_unsigned(2828, 12), 1358 => to_unsigned(1121, 12), 1359 => to_unsigned(3099, 12), 1360 => to_unsigned(2972, 12), 1361 => to_unsigned(710, 12), 1362 => to_unsigned(750, 12), 1363 => to_unsigned(1548, 12), 1364 => to_unsigned(1911, 12), 1365 => to_unsigned(2239, 12), 1366 => to_unsigned(2848, 12), 1367 => to_unsigned(3057, 12), 1368 => to_unsigned(577, 12), 1369 => to_unsigned(2022, 12), 1370 => to_unsigned(827, 12), 1371 => to_unsigned(3473, 12), 1372 => to_unsigned(1749, 12), 1373 => to_unsigned(3954, 12), 1374 => to_unsigned(783, 12), 1375 => to_unsigned(630, 12), 1376 => to_unsigned(2724, 12), 1377 => to_unsigned(1011, 12), 1378 => to_unsigned(91, 12), 1379 => to_unsigned(405, 12), 1380 => to_unsigned(2868, 12), 1381 => to_unsigned(1133, 12), 1382 => to_unsigned(63, 12), 1383 => to_unsigned(1574, 12), 1384 => to_unsigned(226, 12), 1385 => to_unsigned(1894, 12), 1386 => to_unsigned(1493, 12), 1387 => to_unsigned(2479, 12), 1388 => to_unsigned(3515, 12), 1389 => to_unsigned(2247, 12), 1390 => to_unsigned(294, 12), 1391 => to_unsigned(2799, 12), 1392 => to_unsigned(3414, 12), 1393 => to_unsigned(3148, 12), 1394 => to_unsigned(3344, 12), 1395 => to_unsigned(2185, 12), 1396 => to_unsigned(1770, 12), 1397 => to_unsigned(281, 12), 1398 => to_unsigned(3165, 12), 1399 => to_unsigned(1112, 12), 1400 => to_unsigned(1183, 12), 1401 => to_unsigned(2692, 12), 1402 => to_unsigned(2056, 12), 1403 => to_unsigned(3001, 12), 1404 => to_unsigned(2930, 12), 1405 => to_unsigned(3040, 12), 1406 => to_unsigned(3788, 12), 1407 => to_unsigned(3096, 12), 1408 => to_unsigned(1563, 12), 1409 => to_unsigned(254, 12), 1410 => to_unsigned(1555, 12), 1411 => to_unsigned(2853, 12), 1412 => to_unsigned(201, 12), 1413 => to_unsigned(1730, 12), 1414 => to_unsigned(491, 12), 1415 => to_unsigned(1453, 12), 1416 => to_unsigned(1870, 12), 1417 => to_unsigned(1511, 12), 1418 => to_unsigned(2331, 12), 1419 => to_unsigned(3612, 12), 1420 => to_unsigned(2830, 12), 1421 => to_unsigned(3775, 12), 1422 => to_unsigned(369, 12), 1423 => to_unsigned(1832, 12), 1424 => to_unsigned(2623, 12), 1425 => to_unsigned(1104, 12), 1426 => to_unsigned(876, 12), 1427 => to_unsigned(672, 12), 1428 => to_unsigned(3055, 12), 1429 => to_unsigned(583, 12), 1430 => to_unsigned(1383, 12), 1431 => to_unsigned(3566, 12), 1432 => to_unsigned(2949, 12), 1433 => to_unsigned(991, 12), 1434 => to_unsigned(2705, 12), 1435 => to_unsigned(628, 12), 1436 => to_unsigned(3710, 12), 1437 => to_unsigned(2287, 12), 1438 => to_unsigned(3201, 12), 1439 => to_unsigned(1382, 12), 1440 => to_unsigned(2378, 12), 1441 => to_unsigned(1627, 12), 1442 => to_unsigned(1506, 12), 1443 => to_unsigned(929, 12), 1444 => to_unsigned(2114, 12), 1445 => to_unsigned(4087, 12), 1446 => to_unsigned(2590, 12), 1447 => to_unsigned(3953, 12), 1448 => to_unsigned(111, 12), 1449 => to_unsigned(906, 12), 1450 => to_unsigned(774, 12), 1451 => to_unsigned(3712, 12), 1452 => to_unsigned(3467, 12), 1453 => to_unsigned(2880, 12), 1454 => to_unsigned(2999, 12), 1455 => to_unsigned(3337, 12), 1456 => to_unsigned(2578, 12), 1457 => to_unsigned(1843, 12), 1458 => to_unsigned(76, 12), 1459 => to_unsigned(434, 12), 1460 => to_unsigned(562, 12), 1461 => to_unsigned(2638, 12), 1462 => to_unsigned(1769, 12), 1463 => to_unsigned(2828, 12), 1464 => to_unsigned(4065, 12), 1465 => to_unsigned(3360, 12), 1466 => to_unsigned(281, 12), 1467 => to_unsigned(1245, 12), 1468 => to_unsigned(3479, 12), 1469 => to_unsigned(791, 12), 1470 => to_unsigned(940, 12), 1471 => to_unsigned(1663, 12), 1472 => to_unsigned(602, 12), 1473 => to_unsigned(3947, 12), 1474 => to_unsigned(2789, 12), 1475 => to_unsigned(2389, 12), 1476 => to_unsigned(2739, 12), 1477 => to_unsigned(117, 12), 1478 => to_unsigned(3299, 12), 1479 => to_unsigned(3118, 12), 1480 => to_unsigned(141, 12), 1481 => to_unsigned(1963, 12), 1482 => to_unsigned(1934, 12), 1483 => to_unsigned(3477, 12), 1484 => to_unsigned(3324, 12), 1485 => to_unsigned(3876, 12), 1486 => to_unsigned(1775, 12), 1487 => to_unsigned(175, 12), 1488 => to_unsigned(3349, 12), 1489 => to_unsigned(2025, 12), 1490 => to_unsigned(2859, 12), 1491 => to_unsigned(1263, 12), 1492 => to_unsigned(1282, 12), 1493 => to_unsigned(2563, 12), 1494 => to_unsigned(1732, 12), 1495 => to_unsigned(1189, 12), 1496 => to_unsigned(1569, 12), 1497 => to_unsigned(2973, 12), 1498 => to_unsigned(2542, 12), 1499 => to_unsigned(3243, 12), 1500 => to_unsigned(340, 12), 1501 => to_unsigned(806, 12), 1502 => to_unsigned(2216, 12), 1503 => to_unsigned(3532, 12), 1504 => to_unsigned(2179, 12), 1505 => to_unsigned(2899, 12), 1506 => to_unsigned(4024, 12), 1507 => to_unsigned(1239, 12), 1508 => to_unsigned(2967, 12), 1509 => to_unsigned(2780, 12), 1510 => to_unsigned(3842, 12), 1511 => to_unsigned(3271, 12), 1512 => to_unsigned(3677, 12), 1513 => to_unsigned(1096, 12), 1514 => to_unsigned(1252, 12), 1515 => to_unsigned(2994, 12), 1516 => to_unsigned(96, 12), 1517 => to_unsigned(4055, 12), 1518 => to_unsigned(1354, 12), 1519 => to_unsigned(788, 12), 1520 => to_unsigned(1261, 12), 1521 => to_unsigned(83, 12), 1522 => to_unsigned(72, 12), 1523 => to_unsigned(1103, 12), 1524 => to_unsigned(1961, 12), 1525 => to_unsigned(1916, 12), 1526 => to_unsigned(694, 12), 1527 => to_unsigned(1704, 12), 1528 => to_unsigned(2027, 12), 1529 => to_unsigned(3557, 12), 1530 => to_unsigned(1344, 12), 1531 => to_unsigned(1747, 12), 1532 => to_unsigned(2263, 12), 1533 => to_unsigned(2118, 12), 1534 => to_unsigned(3156, 12), 1535 => to_unsigned(125, 12), 1536 => to_unsigned(1926, 12), 1537 => to_unsigned(3940, 12), 1538 => to_unsigned(495, 12), 1539 => to_unsigned(3522, 12), 1540 => to_unsigned(1298, 12), 1541 => to_unsigned(3031, 12), 1542 => to_unsigned(2847, 12), 1543 => to_unsigned(3020, 12), 1544 => to_unsigned(2099, 12), 1545 => to_unsigned(1590, 12), 1546 => to_unsigned(793, 12), 1547 => to_unsigned(3225, 12), 1548 => to_unsigned(3066, 12), 1549 => to_unsigned(2564, 12), 1550 => to_unsigned(2798, 12), 1551 => to_unsigned(3094, 12), 1552 => to_unsigned(438, 12), 1553 => to_unsigned(881, 12), 1554 => to_unsigned(1122, 12), 1555 => to_unsigned(3033, 12), 1556 => to_unsigned(423, 12), 1557 => to_unsigned(3498, 12), 1558 => to_unsigned(226, 12), 1559 => to_unsigned(2872, 12), 1560 => to_unsigned(2326, 12), 1561 => to_unsigned(3397, 12), 1562 => to_unsigned(1218, 12), 1563 => to_unsigned(4075, 12), 1564 => to_unsigned(2290, 12), 1565 => to_unsigned(3325, 12), 1566 => to_unsigned(4059, 12), 1567 => to_unsigned(521, 12), 1568 => to_unsigned(1106, 12), 1569 => to_unsigned(2330, 12), 1570 => to_unsigned(103, 12), 1571 => to_unsigned(262, 12), 1572 => to_unsigned(2317, 12), 1573 => to_unsigned(3024, 12), 1574 => to_unsigned(1376, 12), 1575 => to_unsigned(2746, 12), 1576 => to_unsigned(3929, 12), 1577 => to_unsigned(2715, 12), 1578 => to_unsigned(1304, 12), 1579 => to_unsigned(1464, 12), 1580 => to_unsigned(214, 12), 1581 => to_unsigned(1100, 12), 1582 => to_unsigned(2716, 12), 1583 => to_unsigned(908, 12), 1584 => to_unsigned(3652, 12), 1585 => to_unsigned(2185, 12), 1586 => to_unsigned(1096, 12), 1587 => to_unsigned(1465, 12), 1588 => to_unsigned(2534, 12), 1589 => to_unsigned(117, 12), 1590 => to_unsigned(3874, 12), 1591 => to_unsigned(41, 12), 1592 => to_unsigned(2112, 12), 1593 => to_unsigned(1808, 12), 1594 => to_unsigned(2393, 12), 1595 => to_unsigned(3759, 12), 1596 => to_unsigned(3923, 12), 1597 => to_unsigned(670, 12), 1598 => to_unsigned(1570, 12), 1599 => to_unsigned(570, 12), 1600 => to_unsigned(1767, 12), 1601 => to_unsigned(3173, 12), 1602 => to_unsigned(3733, 12), 1603 => to_unsigned(3896, 12), 1604 => to_unsigned(2632, 12), 1605 => to_unsigned(1732, 12), 1606 => to_unsigned(4042, 12), 1607 => to_unsigned(139, 12), 1608 => to_unsigned(763, 12), 1609 => to_unsigned(1029, 12), 1610 => to_unsigned(944, 12), 1611 => to_unsigned(1351, 12), 1612 => to_unsigned(3963, 12), 1613 => to_unsigned(359, 12), 1614 => to_unsigned(3264, 12), 1615 => to_unsigned(3876, 12), 1616 => to_unsigned(1310, 12), 1617 => to_unsigned(3908, 12), 1618 => to_unsigned(3457, 12), 1619 => to_unsigned(2386, 12), 1620 => to_unsigned(1086, 12), 1621 => to_unsigned(1394, 12), 1622 => to_unsigned(1692, 12), 1623 => to_unsigned(1585, 12), 1624 => to_unsigned(1987, 12), 1625 => to_unsigned(1916, 12), 1626 => to_unsigned(1310, 12), 1627 => to_unsigned(549, 12), 1628 => to_unsigned(790, 12), 1629 => to_unsigned(1015, 12), 1630 => to_unsigned(480, 12), 1631 => to_unsigned(3197, 12), 1632 => to_unsigned(2026, 12), 1633 => to_unsigned(2028, 12), 1634 => to_unsigned(2642, 12), 1635 => to_unsigned(508, 12), 1636 => to_unsigned(1579, 12), 1637 => to_unsigned(116, 12), 1638 => to_unsigned(1338, 12), 1639 => to_unsigned(907, 12), 1640 => to_unsigned(1594, 12), 1641 => to_unsigned(3316, 12), 1642 => to_unsigned(3674, 12), 1643 => to_unsigned(3589, 12), 1644 => to_unsigned(83, 12), 1645 => to_unsigned(3542, 12), 1646 => to_unsigned(2030, 12), 1647 => to_unsigned(1534, 12), 1648 => to_unsigned(1720, 12), 1649 => to_unsigned(634, 12), 1650 => to_unsigned(2884, 12), 1651 => to_unsigned(2267, 12), 1652 => to_unsigned(2861, 12), 1653 => to_unsigned(3405, 12), 1654 => to_unsigned(197, 12), 1655 => to_unsigned(3054, 12), 1656 => to_unsigned(3330, 12), 1657 => to_unsigned(1193, 12), 1658 => to_unsigned(562, 12), 1659 => to_unsigned(1853, 12), 1660 => to_unsigned(3416, 12), 1661 => to_unsigned(3245, 12), 1662 => to_unsigned(1979, 12), 1663 => to_unsigned(1453, 12), 1664 => to_unsigned(3037, 12), 1665 => to_unsigned(668, 12), 1666 => to_unsigned(2885, 12), 1667 => to_unsigned(737, 12), 1668 => to_unsigned(1945, 12), 1669 => to_unsigned(1760, 12), 1670 => to_unsigned(732, 12), 1671 => to_unsigned(2653, 12), 1672 => to_unsigned(3435, 12), 1673 => to_unsigned(3273, 12), 1674 => to_unsigned(2117, 12), 1675 => to_unsigned(4090, 12), 1676 => to_unsigned(916, 12), 1677 => to_unsigned(2392, 12), 1678 => to_unsigned(2814, 12), 1679 => to_unsigned(2524, 12), 1680 => to_unsigned(536, 12), 1681 => to_unsigned(1269, 12), 1682 => to_unsigned(1809, 12), 1683 => to_unsigned(1196, 12), 1684 => to_unsigned(2370, 12), 1685 => to_unsigned(3355, 12), 1686 => to_unsigned(25, 12), 1687 => to_unsigned(3770, 12), 1688 => to_unsigned(1168, 12), 1689 => to_unsigned(2080, 12), 1690 => to_unsigned(614, 12), 1691 => to_unsigned(2142, 12), 1692 => to_unsigned(1071, 12), 1693 => to_unsigned(3333, 12), 1694 => to_unsigned(40, 12), 1695 => to_unsigned(146, 12), 1696 => to_unsigned(2842, 12), 1697 => to_unsigned(1380, 12), 1698 => to_unsigned(3247, 12), 1699 => to_unsigned(1911, 12), 1700 => to_unsigned(498, 12), 1701 => to_unsigned(3867, 12), 1702 => to_unsigned(1838, 12), 1703 => to_unsigned(1266, 12), 1704 => to_unsigned(3747, 12), 1705 => to_unsigned(3735, 12), 1706 => to_unsigned(2360, 12), 1707 => to_unsigned(3210, 12), 1708 => to_unsigned(948, 12), 1709 => to_unsigned(1660, 12), 1710 => to_unsigned(1663, 12), 1711 => to_unsigned(442, 12), 1712 => to_unsigned(394, 12), 1713 => to_unsigned(3779, 12), 1714 => to_unsigned(3083, 12), 1715 => to_unsigned(3080, 12), 1716 => to_unsigned(4087, 12), 1717 => to_unsigned(3217, 12), 1718 => to_unsigned(3021, 12), 1719 => to_unsigned(2901, 12), 1720 => to_unsigned(936, 12), 1721 => to_unsigned(1033, 12), 1722 => to_unsigned(1674, 12), 1723 => to_unsigned(2710, 12), 1724 => to_unsigned(1501, 12), 1725 => to_unsigned(1494, 12), 1726 => to_unsigned(361, 12), 1727 => to_unsigned(1757, 12), 1728 => to_unsigned(126, 12), 1729 => to_unsigned(3681, 12), 1730 => to_unsigned(586, 12), 1731 => to_unsigned(199, 12), 1732 => to_unsigned(1742, 12), 1733 => to_unsigned(3178, 12), 1734 => to_unsigned(1718, 12), 1735 => to_unsigned(99, 12), 1736 => to_unsigned(2118, 12), 1737 => to_unsigned(408, 12), 1738 => to_unsigned(890, 12), 1739 => to_unsigned(1899, 12), 1740 => to_unsigned(1352, 12), 1741 => to_unsigned(3507, 12), 1742 => to_unsigned(2306, 12), 1743 => to_unsigned(2215, 12), 1744 => to_unsigned(3502, 12), 1745 => to_unsigned(2857, 12), 1746 => to_unsigned(909, 12), 1747 => to_unsigned(2836, 12), 1748 => to_unsigned(3137, 12), 1749 => to_unsigned(2898, 12), 1750 => to_unsigned(3404, 12), 1751 => to_unsigned(3457, 12), 1752 => to_unsigned(649, 12), 1753 => to_unsigned(3670, 12), 1754 => to_unsigned(1410, 12), 1755 => to_unsigned(572, 12), 1756 => to_unsigned(2489, 12), 1757 => to_unsigned(204, 12), 1758 => to_unsigned(2325, 12), 1759 => to_unsigned(1242, 12), 1760 => to_unsigned(2054, 12), 1761 => to_unsigned(3236, 12), 1762 => to_unsigned(1922, 12), 1763 => to_unsigned(316, 12), 1764 => to_unsigned(3770, 12), 1765 => to_unsigned(357, 12), 1766 => to_unsigned(1088, 12), 1767 => to_unsigned(2956, 12), 1768 => to_unsigned(48, 12), 1769 => to_unsigned(1965, 12), 1770 => to_unsigned(1810, 12), 1771 => to_unsigned(2340, 12), 1772 => to_unsigned(2042, 12), 1773 => to_unsigned(3577, 12), 1774 => to_unsigned(3184, 12), 1775 => to_unsigned(1888, 12), 1776 => to_unsigned(881, 12), 1777 => to_unsigned(3438, 12), 1778 => to_unsigned(2825, 12), 1779 => to_unsigned(2083, 12), 1780 => to_unsigned(3196, 12), 1781 => to_unsigned(1055, 12), 1782 => to_unsigned(251, 12), 1783 => to_unsigned(2678, 12), 1784 => to_unsigned(3994, 12), 1785 => to_unsigned(586, 12), 1786 => to_unsigned(402, 12), 1787 => to_unsigned(3005, 12), 1788 => to_unsigned(3839, 12), 1789 => to_unsigned(3337, 12), 1790 => to_unsigned(1810, 12), 1791 => to_unsigned(1941, 12), 1792 => to_unsigned(3248, 12), 1793 => to_unsigned(3089, 12), 1794 => to_unsigned(4077, 12), 1795 => to_unsigned(724, 12), 1796 => to_unsigned(882, 12), 1797 => to_unsigned(2637, 12), 1798 => to_unsigned(2203, 12), 1799 => to_unsigned(243, 12), 1800 => to_unsigned(1463, 12), 1801 => to_unsigned(1127, 12), 1802 => to_unsigned(2038, 12), 1803 => to_unsigned(2281, 12), 1804 => to_unsigned(1119, 12), 1805 => to_unsigned(2263, 12), 1806 => to_unsigned(3797, 12), 1807 => to_unsigned(78, 12), 1808 => to_unsigned(1122, 12), 1809 => to_unsigned(2196, 12), 1810 => to_unsigned(1310, 12), 1811 => to_unsigned(1620, 12), 1812 => to_unsigned(3526, 12), 1813 => to_unsigned(957, 12), 1814 => to_unsigned(1763, 12), 1815 => to_unsigned(686, 12), 1816 => to_unsigned(2997, 12), 1817 => to_unsigned(1029, 12), 1818 => to_unsigned(2454, 12), 1819 => to_unsigned(4013, 12), 1820 => to_unsigned(3892, 12), 1821 => to_unsigned(766, 12), 1822 => to_unsigned(1364, 12), 1823 => to_unsigned(3112, 12), 1824 => to_unsigned(1854, 12), 1825 => to_unsigned(1266, 12), 1826 => to_unsigned(1199, 12), 1827 => to_unsigned(2995, 12), 1828 => to_unsigned(3603, 12), 1829 => to_unsigned(301, 12), 1830 => to_unsigned(2965, 12), 1831 => to_unsigned(1701, 12), 1832 => to_unsigned(3796, 12), 1833 => to_unsigned(2035, 12), 1834 => to_unsigned(3511, 12), 1835 => to_unsigned(1175, 12), 1836 => to_unsigned(3289, 12), 1837 => to_unsigned(1433, 12), 1838 => to_unsigned(1614, 12), 1839 => to_unsigned(2168, 12), 1840 => to_unsigned(3151, 12), 1841 => to_unsigned(2359, 12), 1842 => to_unsigned(3373, 12), 1843 => to_unsigned(2704, 12), 1844 => to_unsigned(509, 12), 1845 => to_unsigned(2302, 12), 1846 => to_unsigned(2952, 12), 1847 => to_unsigned(4042, 12), 1848 => to_unsigned(618, 12), 1849 => to_unsigned(1429, 12), 1850 => to_unsigned(1808, 12), 1851 => to_unsigned(2398, 12), 1852 => to_unsigned(3004, 12), 1853 => to_unsigned(2454, 12), 1854 => to_unsigned(2668, 12), 1855 => to_unsigned(1625, 12), 1856 => to_unsigned(1819, 12), 1857 => to_unsigned(2985, 12), 1858 => to_unsigned(2515, 12), 1859 => to_unsigned(2078, 12), 1860 => to_unsigned(2043, 12), 1861 => to_unsigned(2218, 12), 1862 => to_unsigned(1594, 12), 1863 => to_unsigned(1895, 12), 1864 => to_unsigned(3489, 12), 1865 => to_unsigned(3477, 12), 1866 => to_unsigned(970, 12), 1867 => to_unsigned(2180, 12), 1868 => to_unsigned(2664, 12), 1869 => to_unsigned(2850, 12), 1870 => to_unsigned(3188, 12), 1871 => to_unsigned(151, 12), 1872 => to_unsigned(1600, 12), 1873 => to_unsigned(1360, 12), 1874 => to_unsigned(4074, 12), 1875 => to_unsigned(2894, 12), 1876 => to_unsigned(4033, 12), 1877 => to_unsigned(201, 12), 1878 => to_unsigned(485, 12), 1879 => to_unsigned(19, 12), 1880 => to_unsigned(320, 12), 1881 => to_unsigned(1155, 12), 1882 => to_unsigned(941, 12), 1883 => to_unsigned(425, 12), 1884 => to_unsigned(1835, 12), 1885 => to_unsigned(631, 12), 1886 => to_unsigned(793, 12), 1887 => to_unsigned(1729, 12), 1888 => to_unsigned(2096, 12), 1889 => to_unsigned(3352, 12), 1890 => to_unsigned(3457, 12), 1891 => to_unsigned(3979, 12), 1892 => to_unsigned(2991, 12), 1893 => to_unsigned(3407, 12), 1894 => to_unsigned(2711, 12), 1895 => to_unsigned(734, 12), 1896 => to_unsigned(2358, 12), 1897 => to_unsigned(660, 12), 1898 => to_unsigned(2020, 12), 1899 => to_unsigned(2562, 12), 1900 => to_unsigned(619, 12), 1901 => to_unsigned(3384, 12), 1902 => to_unsigned(1879, 12), 1903 => to_unsigned(1513, 12), 1904 => to_unsigned(605, 12), 1905 => to_unsigned(3505, 12), 1906 => to_unsigned(699, 12), 1907 => to_unsigned(3874, 12), 1908 => to_unsigned(2468, 12), 1909 => to_unsigned(1373, 12), 1910 => to_unsigned(1283, 12), 1911 => to_unsigned(1595, 12), 1912 => to_unsigned(3483, 12), 1913 => to_unsigned(2771, 12), 1914 => to_unsigned(2851, 12), 1915 => to_unsigned(3844, 12), 1916 => to_unsigned(2908, 12), 1917 => to_unsigned(3891, 12), 1918 => to_unsigned(139, 12), 1919 => to_unsigned(3950, 12), 1920 => to_unsigned(1289, 12), 1921 => to_unsigned(2252, 12), 1922 => to_unsigned(2965, 12), 1923 => to_unsigned(3357, 12), 1924 => to_unsigned(2481, 12), 1925 => to_unsigned(2289, 12), 1926 => to_unsigned(707, 12), 1927 => to_unsigned(2758, 12), 1928 => to_unsigned(851, 12), 1929 => to_unsigned(3096, 12), 1930 => to_unsigned(157, 12), 1931 => to_unsigned(2458, 12), 1932 => to_unsigned(3662, 12), 1933 => to_unsigned(4025, 12), 1934 => to_unsigned(1891, 12), 1935 => to_unsigned(741, 12), 1936 => to_unsigned(1201, 12), 1937 => to_unsigned(2413, 12), 1938 => to_unsigned(3403, 12), 1939 => to_unsigned(2945, 12), 1940 => to_unsigned(641, 12), 1941 => to_unsigned(546, 12), 1942 => to_unsigned(878, 12), 1943 => to_unsigned(3051, 12), 1944 => to_unsigned(2130, 12), 1945 => to_unsigned(1014, 12), 1946 => to_unsigned(3028, 12), 1947 => to_unsigned(3369, 12), 1948 => to_unsigned(3846, 12), 1949 => to_unsigned(808, 12), 1950 => to_unsigned(2391, 12), 1951 => to_unsigned(228, 12), 1952 => to_unsigned(2776, 12), 1953 => to_unsigned(3096, 12), 1954 => to_unsigned(626, 12), 1955 => to_unsigned(2670, 12), 1956 => to_unsigned(224, 12), 1957 => to_unsigned(726, 12), 1958 => to_unsigned(274, 12), 1959 => to_unsigned(3727, 12), 1960 => to_unsigned(2215, 12), 1961 => to_unsigned(1626, 12), 1962 => to_unsigned(2483, 12), 1963 => to_unsigned(3687, 12), 1964 => to_unsigned(329, 12), 1965 => to_unsigned(900, 12), 1966 => to_unsigned(2625, 12), 1967 => to_unsigned(2074, 12), 1968 => to_unsigned(2269, 12), 1969 => to_unsigned(1951, 12), 1970 => to_unsigned(3677, 12), 1971 => to_unsigned(549, 12), 1972 => to_unsigned(530, 12), 1973 => to_unsigned(3419, 12), 1974 => to_unsigned(2095, 12), 1975 => to_unsigned(3872, 12), 1976 => to_unsigned(2417, 12), 1977 => to_unsigned(2615, 12), 1978 => to_unsigned(1035, 12), 1979 => to_unsigned(699, 12), 1980 => to_unsigned(3482, 12), 1981 => to_unsigned(3260, 12), 1982 => to_unsigned(3009, 12), 1983 => to_unsigned(3301, 12), 1984 => to_unsigned(3521, 12), 1985 => to_unsigned(1191, 12), 1986 => to_unsigned(4087, 12), 1987 => to_unsigned(396, 12), 1988 => to_unsigned(348, 12), 1989 => to_unsigned(2965, 12), 1990 => to_unsigned(2011, 12), 1991 => to_unsigned(3974, 12), 1992 => to_unsigned(2672, 12), 1993 => to_unsigned(3413, 12), 1994 => to_unsigned(3222, 12), 1995 => to_unsigned(3927, 12), 1996 => to_unsigned(3616, 12), 1997 => to_unsigned(3032, 12), 1998 => to_unsigned(98, 12), 1999 => to_unsigned(1695, 12), 2000 => to_unsigned(2336, 12), 2001 => to_unsigned(1260, 12), 2002 => to_unsigned(1181, 12), 2003 => to_unsigned(1318, 12), 2004 => to_unsigned(3454, 12), 2005 => to_unsigned(568, 12), 2006 => to_unsigned(80, 12), 2007 => to_unsigned(3652, 12), 2008 => to_unsigned(3010, 12), 2009 => to_unsigned(3246, 12), 2010 => to_unsigned(2462, 12), 2011 => to_unsigned(221, 12), 2012 => to_unsigned(3111, 12), 2013 => to_unsigned(1002, 12), 2014 => to_unsigned(2697, 12), 2015 => to_unsigned(1591, 12), 2016 => to_unsigned(2650, 12), 2017 => to_unsigned(198, 12), 2018 => to_unsigned(3237, 12), 2019 => to_unsigned(1241, 12), 2020 => to_unsigned(1706, 12), 2021 => to_unsigned(1588, 12), 2022 => to_unsigned(3030, 12), 2023 => to_unsigned(2938, 12), 2024 => to_unsigned(1150, 12), 2025 => to_unsigned(1474, 12), 2026 => to_unsigned(2465, 12), 2027 => to_unsigned(435, 12), 2028 => to_unsigned(696, 12), 2029 => to_unsigned(1802, 12), 2030 => to_unsigned(818, 12), 2031 => to_unsigned(2403, 12), 2032 => to_unsigned(2339, 12), 2033 => to_unsigned(3841, 12), 2034 => to_unsigned(3286, 12), 2035 => to_unsigned(2638, 12), 2036 => to_unsigned(1465, 12), 2037 => to_unsigned(289, 12), 2038 => to_unsigned(2888, 12), 2039 => to_unsigned(3990, 12), 2040 => to_unsigned(3947, 12), 2041 => to_unsigned(3647, 12), 2042 => to_unsigned(449, 12), 2043 => to_unsigned(1203, 12), 2044 => to_unsigned(1312, 12), 2045 => to_unsigned(3562, 12), 2046 => to_unsigned(3235, 12), 2047 => to_unsigned(1856, 12)),
            5 => (0 => to_unsigned(84, 12), 1 => to_unsigned(3005, 12), 2 => to_unsigned(1561, 12), 3 => to_unsigned(2131, 12), 4 => to_unsigned(1, 12), 5 => to_unsigned(1078, 12), 6 => to_unsigned(2907, 12), 7 => to_unsigned(1124, 12), 8 => to_unsigned(2752, 12), 9 => to_unsigned(2634, 12), 10 => to_unsigned(2608, 12), 11 => to_unsigned(1986, 12), 12 => to_unsigned(1292, 12), 13 => to_unsigned(958, 12), 14 => to_unsigned(437, 12), 15 => to_unsigned(2636, 12), 16 => to_unsigned(3280, 12), 17 => to_unsigned(2551, 12), 18 => to_unsigned(323, 12), 19 => to_unsigned(3706, 12), 20 => to_unsigned(1833, 12), 21 => to_unsigned(2766, 12), 22 => to_unsigned(4081, 12), 23 => to_unsigned(1911, 12), 24 => to_unsigned(2676, 12), 25 => to_unsigned(255, 12), 26 => to_unsigned(3049, 12), 27 => to_unsigned(2773, 12), 28 => to_unsigned(3020, 12), 29 => to_unsigned(241, 12), 30 => to_unsigned(861, 12), 31 => to_unsigned(1400, 12), 32 => to_unsigned(2956, 12), 33 => to_unsigned(1082, 12), 34 => to_unsigned(3273, 12), 35 => to_unsigned(475, 12), 36 => to_unsigned(1249, 12), 37 => to_unsigned(293, 12), 38 => to_unsigned(2094, 12), 39 => to_unsigned(699, 12), 40 => to_unsigned(1359, 12), 41 => to_unsigned(722, 12), 42 => to_unsigned(123, 12), 43 => to_unsigned(1509, 12), 44 => to_unsigned(1641, 12), 45 => to_unsigned(2418, 12), 46 => to_unsigned(2031, 12), 47 => to_unsigned(2215, 12), 48 => to_unsigned(3852, 12), 49 => to_unsigned(3609, 12), 50 => to_unsigned(3878, 12), 51 => to_unsigned(2307, 12), 52 => to_unsigned(3076, 12), 53 => to_unsigned(1695, 12), 54 => to_unsigned(2919, 12), 55 => to_unsigned(1365, 12), 56 => to_unsigned(1985, 12), 57 => to_unsigned(439, 12), 58 => to_unsigned(2170, 12), 59 => to_unsigned(3783, 12), 60 => to_unsigned(3310, 12), 61 => to_unsigned(3583, 12), 62 => to_unsigned(2576, 12), 63 => to_unsigned(3143, 12), 64 => to_unsigned(1101, 12), 65 => to_unsigned(2554, 12), 66 => to_unsigned(1897, 12), 67 => to_unsigned(1241, 12), 68 => to_unsigned(1995, 12), 69 => to_unsigned(509, 12), 70 => to_unsigned(99, 12), 71 => to_unsigned(3513, 12), 72 => to_unsigned(2942, 12), 73 => to_unsigned(2557, 12), 74 => to_unsigned(1090, 12), 75 => to_unsigned(3149, 12), 76 => to_unsigned(2563, 12), 77 => to_unsigned(3019, 12), 78 => to_unsigned(3457, 12), 79 => to_unsigned(480, 12), 80 => to_unsigned(3395, 12), 81 => to_unsigned(3720, 12), 82 => to_unsigned(3249, 12), 83 => to_unsigned(2568, 12), 84 => to_unsigned(2853, 12), 85 => to_unsigned(106, 12), 86 => to_unsigned(817, 12), 87 => to_unsigned(769, 12), 88 => to_unsigned(3414, 12), 89 => to_unsigned(69, 12), 90 => to_unsigned(3755, 12), 91 => to_unsigned(1897, 12), 92 => to_unsigned(1323, 12), 93 => to_unsigned(1700, 12), 94 => to_unsigned(3945, 12), 95 => to_unsigned(3368, 12), 96 => to_unsigned(3748, 12), 97 => to_unsigned(3892, 12), 98 => to_unsigned(2546, 12), 99 => to_unsigned(845, 12), 100 => to_unsigned(37, 12), 101 => to_unsigned(3757, 12), 102 => to_unsigned(41, 12), 103 => to_unsigned(2873, 12), 104 => to_unsigned(2248, 12), 105 => to_unsigned(3161, 12), 106 => to_unsigned(1304, 12), 107 => to_unsigned(901, 12), 108 => to_unsigned(2053, 12), 109 => to_unsigned(1444, 12), 110 => to_unsigned(1381, 12), 111 => to_unsigned(260, 12), 112 => to_unsigned(3663, 12), 113 => to_unsigned(2490, 12), 114 => to_unsigned(711, 12), 115 => to_unsigned(2455, 12), 116 => to_unsigned(2722, 12), 117 => to_unsigned(1993, 12), 118 => to_unsigned(521, 12), 119 => to_unsigned(440, 12), 120 => to_unsigned(3246, 12), 121 => to_unsigned(3619, 12), 122 => to_unsigned(3935, 12), 123 => to_unsigned(959, 12), 124 => to_unsigned(3016, 12), 125 => to_unsigned(562, 12), 126 => to_unsigned(3527, 12), 127 => to_unsigned(3128, 12), 128 => to_unsigned(453, 12), 129 => to_unsigned(2399, 12), 130 => to_unsigned(3983, 12), 131 => to_unsigned(2008, 12), 132 => to_unsigned(3926, 12), 133 => to_unsigned(511, 12), 134 => to_unsigned(1030, 12), 135 => to_unsigned(2086, 12), 136 => to_unsigned(2416, 12), 137 => to_unsigned(2792, 12), 138 => to_unsigned(589, 12), 139 => to_unsigned(4089, 12), 140 => to_unsigned(3346, 12), 141 => to_unsigned(3524, 12), 142 => to_unsigned(1412, 12), 143 => to_unsigned(1534, 12), 144 => to_unsigned(2036, 12), 145 => to_unsigned(1270, 12), 146 => to_unsigned(1990, 12), 147 => to_unsigned(3177, 12), 148 => to_unsigned(894, 12), 149 => to_unsigned(3532, 12), 150 => to_unsigned(2116, 12), 151 => to_unsigned(939, 12), 152 => to_unsigned(1177, 12), 153 => to_unsigned(576, 12), 154 => to_unsigned(1109, 12), 155 => to_unsigned(2299, 12), 156 => to_unsigned(3716, 12), 157 => to_unsigned(190, 12), 158 => to_unsigned(4092, 12), 159 => to_unsigned(804, 12), 160 => to_unsigned(3364, 12), 161 => to_unsigned(626, 12), 162 => to_unsigned(1212, 12), 163 => to_unsigned(2074, 12), 164 => to_unsigned(1854, 12), 165 => to_unsigned(1214, 12), 166 => to_unsigned(3741, 12), 167 => to_unsigned(1896, 12), 168 => to_unsigned(2462, 12), 169 => to_unsigned(207, 12), 170 => to_unsigned(3267, 12), 171 => to_unsigned(340, 12), 172 => to_unsigned(2039, 12), 173 => to_unsigned(630, 12), 174 => to_unsigned(3794, 12), 175 => to_unsigned(2151, 12), 176 => to_unsigned(830, 12), 177 => to_unsigned(3768, 12), 178 => to_unsigned(653, 12), 179 => to_unsigned(1559, 12), 180 => to_unsigned(3484, 12), 181 => to_unsigned(508, 12), 182 => to_unsigned(91, 12), 183 => to_unsigned(2153, 12), 184 => to_unsigned(3664, 12), 185 => to_unsigned(2802, 12), 186 => to_unsigned(2047, 12), 187 => to_unsigned(2309, 12), 188 => to_unsigned(450, 12), 189 => to_unsigned(57, 12), 190 => to_unsigned(2828, 12), 191 => to_unsigned(3716, 12), 192 => to_unsigned(3093, 12), 193 => to_unsigned(1217, 12), 194 => to_unsigned(2555, 12), 195 => to_unsigned(2805, 12), 196 => to_unsigned(3995, 12), 197 => to_unsigned(3230, 12), 198 => to_unsigned(3173, 12), 199 => to_unsigned(2032, 12), 200 => to_unsigned(1347, 12), 201 => to_unsigned(384, 12), 202 => to_unsigned(3111, 12), 203 => to_unsigned(3272, 12), 204 => to_unsigned(478, 12), 205 => to_unsigned(2673, 12), 206 => to_unsigned(2220, 12), 207 => to_unsigned(1571, 12), 208 => to_unsigned(780, 12), 209 => to_unsigned(2500, 12), 210 => to_unsigned(1240, 12), 211 => to_unsigned(445, 12), 212 => to_unsigned(1369, 12), 213 => to_unsigned(548, 12), 214 => to_unsigned(3139, 12), 215 => to_unsigned(951, 12), 216 => to_unsigned(3588, 12), 217 => to_unsigned(109, 12), 218 => to_unsigned(3043, 12), 219 => to_unsigned(1404, 12), 220 => to_unsigned(1794, 12), 221 => to_unsigned(1620, 12), 222 => to_unsigned(2852, 12), 223 => to_unsigned(3540, 12), 224 => to_unsigned(3213, 12), 225 => to_unsigned(3616, 12), 226 => to_unsigned(1820, 12), 227 => to_unsigned(168, 12), 228 => to_unsigned(1319, 12), 229 => to_unsigned(3969, 12), 230 => to_unsigned(2529, 12), 231 => to_unsigned(579, 12), 232 => to_unsigned(3365, 12), 233 => to_unsigned(3265, 12), 234 => to_unsigned(351, 12), 235 => to_unsigned(3779, 12), 236 => to_unsigned(488, 12), 237 => to_unsigned(899, 12), 238 => to_unsigned(1827, 12), 239 => to_unsigned(1250, 12), 240 => to_unsigned(90, 12), 241 => to_unsigned(3750, 12), 242 => to_unsigned(3375, 12), 243 => to_unsigned(888, 12), 244 => to_unsigned(2266, 12), 245 => to_unsigned(2424, 12), 246 => to_unsigned(2726, 12), 247 => to_unsigned(3009, 12), 248 => to_unsigned(97, 12), 249 => to_unsigned(3635, 12), 250 => to_unsigned(3166, 12), 251 => to_unsigned(1910, 12), 252 => to_unsigned(3855, 12), 253 => to_unsigned(876, 12), 254 => to_unsigned(3062, 12), 255 => to_unsigned(1893, 12), 256 => to_unsigned(3262, 12), 257 => to_unsigned(2475, 12), 258 => to_unsigned(2405, 12), 259 => to_unsigned(2662, 12), 260 => to_unsigned(2426, 12), 261 => to_unsigned(3738, 12), 262 => to_unsigned(2996, 12), 263 => to_unsigned(175, 12), 264 => to_unsigned(1472, 12), 265 => to_unsigned(2046, 12), 266 => to_unsigned(3376, 12), 267 => to_unsigned(1666, 12), 268 => to_unsigned(2788, 12), 269 => to_unsigned(1207, 12), 270 => to_unsigned(170, 12), 271 => to_unsigned(2254, 12), 272 => to_unsigned(472, 12), 273 => to_unsigned(2943, 12), 274 => to_unsigned(1618, 12), 275 => to_unsigned(2152, 12), 276 => to_unsigned(3078, 12), 277 => to_unsigned(515, 12), 278 => to_unsigned(3934, 12), 279 => to_unsigned(622, 12), 280 => to_unsigned(2998, 12), 281 => to_unsigned(2126, 12), 282 => to_unsigned(3551, 12), 283 => to_unsigned(3862, 12), 284 => to_unsigned(1808, 12), 285 => to_unsigned(2577, 12), 286 => to_unsigned(2442, 12), 287 => to_unsigned(657, 12), 288 => to_unsigned(1725, 12), 289 => to_unsigned(3653, 12), 290 => to_unsigned(568, 12), 291 => to_unsigned(3735, 12), 292 => to_unsigned(3963, 12), 293 => to_unsigned(227, 12), 294 => to_unsigned(3385, 12), 295 => to_unsigned(2226, 12), 296 => to_unsigned(1667, 12), 297 => to_unsigned(941, 12), 298 => to_unsigned(2942, 12), 299 => to_unsigned(3355, 12), 300 => to_unsigned(702, 12), 301 => to_unsigned(3972, 12), 302 => to_unsigned(517, 12), 303 => to_unsigned(1652, 12), 304 => to_unsigned(498, 12), 305 => to_unsigned(3241, 12), 306 => to_unsigned(1526, 12), 307 => to_unsigned(3690, 12), 308 => to_unsigned(650, 12), 309 => to_unsigned(2239, 12), 310 => to_unsigned(2908, 12), 311 => to_unsigned(2615, 12), 312 => to_unsigned(3084, 12), 313 => to_unsigned(945, 12), 314 => to_unsigned(945, 12), 315 => to_unsigned(227, 12), 316 => to_unsigned(4003, 12), 317 => to_unsigned(3808, 12), 318 => to_unsigned(1612, 12), 319 => to_unsigned(2279, 12), 320 => to_unsigned(2992, 12), 321 => to_unsigned(1110, 12), 322 => to_unsigned(2515, 12), 323 => to_unsigned(3702, 12), 324 => to_unsigned(659, 12), 325 => to_unsigned(3009, 12), 326 => to_unsigned(2947, 12), 327 => to_unsigned(1217, 12), 328 => to_unsigned(1245, 12), 329 => to_unsigned(1122, 12), 330 => to_unsigned(2217, 12), 331 => to_unsigned(898, 12), 332 => to_unsigned(810, 12), 333 => to_unsigned(1096, 12), 334 => to_unsigned(1385, 12), 335 => to_unsigned(2052, 12), 336 => to_unsigned(1194, 12), 337 => to_unsigned(2878, 12), 338 => to_unsigned(2769, 12), 339 => to_unsigned(3002, 12), 340 => to_unsigned(915, 12), 341 => to_unsigned(53, 12), 342 => to_unsigned(3916, 12), 343 => to_unsigned(10, 12), 344 => to_unsigned(3833, 12), 345 => to_unsigned(1149, 12), 346 => to_unsigned(3704, 12), 347 => to_unsigned(708, 12), 348 => to_unsigned(891, 12), 349 => to_unsigned(3078, 12), 350 => to_unsigned(3333, 12), 351 => to_unsigned(284, 12), 352 => to_unsigned(1225, 12), 353 => to_unsigned(2272, 12), 354 => to_unsigned(3180, 12), 355 => to_unsigned(945, 12), 356 => to_unsigned(1850, 12), 357 => to_unsigned(3781, 12), 358 => to_unsigned(880, 12), 359 => to_unsigned(810, 12), 360 => to_unsigned(1853, 12), 361 => to_unsigned(3539, 12), 362 => to_unsigned(3568, 12), 363 => to_unsigned(288, 12), 364 => to_unsigned(1345, 12), 365 => to_unsigned(1328, 12), 366 => to_unsigned(19, 12), 367 => to_unsigned(1825, 12), 368 => to_unsigned(1805, 12), 369 => to_unsigned(1412, 12), 370 => to_unsigned(1878, 12), 371 => to_unsigned(2228, 12), 372 => to_unsigned(2018, 12), 373 => to_unsigned(2983, 12), 374 => to_unsigned(1537, 12), 375 => to_unsigned(654, 12), 376 => to_unsigned(923, 12), 377 => to_unsigned(1855, 12), 378 => to_unsigned(1480, 12), 379 => to_unsigned(3152, 12), 380 => to_unsigned(2637, 12), 381 => to_unsigned(1071, 12), 382 => to_unsigned(3730, 12), 383 => to_unsigned(559, 12), 384 => to_unsigned(2284, 12), 385 => to_unsigned(1325, 12), 386 => to_unsigned(666, 12), 387 => to_unsigned(3975, 12), 388 => to_unsigned(2202, 12), 389 => to_unsigned(1381, 12), 390 => to_unsigned(3897, 12), 391 => to_unsigned(2730, 12), 392 => to_unsigned(1701, 12), 393 => to_unsigned(48, 12), 394 => to_unsigned(318, 12), 395 => to_unsigned(1798, 12), 396 => to_unsigned(2786, 12), 397 => to_unsigned(2722, 12), 398 => to_unsigned(2656, 12), 399 => to_unsigned(1191, 12), 400 => to_unsigned(1975, 12), 401 => to_unsigned(3562, 12), 402 => to_unsigned(3022, 12), 403 => to_unsigned(2982, 12), 404 => to_unsigned(1978, 12), 405 => to_unsigned(176, 12), 406 => to_unsigned(3307, 12), 407 => to_unsigned(1841, 12), 408 => to_unsigned(3347, 12), 409 => to_unsigned(551, 12), 410 => to_unsigned(484, 12), 411 => to_unsigned(3139, 12), 412 => to_unsigned(65, 12), 413 => to_unsigned(2609, 12), 414 => to_unsigned(3746, 12), 415 => to_unsigned(1798, 12), 416 => to_unsigned(2790, 12), 417 => to_unsigned(1111, 12), 418 => to_unsigned(2525, 12), 419 => to_unsigned(44, 12), 420 => to_unsigned(3785, 12), 421 => to_unsigned(3226, 12), 422 => to_unsigned(1432, 12), 423 => to_unsigned(3381, 12), 424 => to_unsigned(1357, 12), 425 => to_unsigned(1757, 12), 426 => to_unsigned(12, 12), 427 => to_unsigned(3138, 12), 428 => to_unsigned(2727, 12), 429 => to_unsigned(15, 12), 430 => to_unsigned(3140, 12), 431 => to_unsigned(613, 12), 432 => to_unsigned(3625, 12), 433 => to_unsigned(2556, 12), 434 => to_unsigned(1267, 12), 435 => to_unsigned(2291, 12), 436 => to_unsigned(3392, 12), 437 => to_unsigned(3416, 12), 438 => to_unsigned(346, 12), 439 => to_unsigned(3348, 12), 440 => to_unsigned(1392, 12), 441 => to_unsigned(2284, 12), 442 => to_unsigned(3677, 12), 443 => to_unsigned(1844, 12), 444 => to_unsigned(3722, 12), 445 => to_unsigned(1626, 12), 446 => to_unsigned(1492, 12), 447 => to_unsigned(1312, 12), 448 => to_unsigned(1127, 12), 449 => to_unsigned(3878, 12), 450 => to_unsigned(1820, 12), 451 => to_unsigned(2135, 12), 452 => to_unsigned(2462, 12), 453 => to_unsigned(4012, 12), 454 => to_unsigned(2238, 12), 455 => to_unsigned(237, 12), 456 => to_unsigned(343, 12), 457 => to_unsigned(2314, 12), 458 => to_unsigned(2148, 12), 459 => to_unsigned(3543, 12), 460 => to_unsigned(1267, 12), 461 => to_unsigned(1757, 12), 462 => to_unsigned(3459, 12), 463 => to_unsigned(2700, 12), 464 => to_unsigned(1520, 12), 465 => to_unsigned(2385, 12), 466 => to_unsigned(246, 12), 467 => to_unsigned(2529, 12), 468 => to_unsigned(36, 12), 469 => to_unsigned(708, 12), 470 => to_unsigned(3393, 12), 471 => to_unsigned(3517, 12), 472 => to_unsigned(2825, 12), 473 => to_unsigned(3143, 12), 474 => to_unsigned(3485, 12), 475 => to_unsigned(4024, 12), 476 => to_unsigned(1109, 12), 477 => to_unsigned(1317, 12), 478 => to_unsigned(2731, 12), 479 => to_unsigned(2022, 12), 480 => to_unsigned(2717, 12), 481 => to_unsigned(1532, 12), 482 => to_unsigned(630, 12), 483 => to_unsigned(1999, 12), 484 => to_unsigned(2022, 12), 485 => to_unsigned(2603, 12), 486 => to_unsigned(51, 12), 487 => to_unsigned(3601, 12), 488 => to_unsigned(2647, 12), 489 => to_unsigned(3410, 12), 490 => to_unsigned(0, 12), 491 => to_unsigned(1249, 12), 492 => to_unsigned(4067, 12), 493 => to_unsigned(1950, 12), 494 => to_unsigned(2938, 12), 495 => to_unsigned(3874, 12), 496 => to_unsigned(1322, 12), 497 => to_unsigned(3637, 12), 498 => to_unsigned(3515, 12), 499 => to_unsigned(3782, 12), 500 => to_unsigned(2585, 12), 501 => to_unsigned(805, 12), 502 => to_unsigned(949, 12), 503 => to_unsigned(292, 12), 504 => to_unsigned(1747, 12), 505 => to_unsigned(2626, 12), 506 => to_unsigned(1735, 12), 507 => to_unsigned(3978, 12), 508 => to_unsigned(146, 12), 509 => to_unsigned(1660, 12), 510 => to_unsigned(1175, 12), 511 => to_unsigned(2103, 12), 512 => to_unsigned(812, 12), 513 => to_unsigned(917, 12), 514 => to_unsigned(1275, 12), 515 => to_unsigned(1100, 12), 516 => to_unsigned(1435, 12), 517 => to_unsigned(2086, 12), 518 => to_unsigned(1427, 12), 519 => to_unsigned(2917, 12), 520 => to_unsigned(2365, 12), 521 => to_unsigned(1647, 12), 522 => to_unsigned(3601, 12), 523 => to_unsigned(1312, 12), 524 => to_unsigned(635, 12), 525 => to_unsigned(3109, 12), 526 => to_unsigned(3781, 12), 527 => to_unsigned(1708, 12), 528 => to_unsigned(3924, 12), 529 => to_unsigned(1864, 12), 530 => to_unsigned(243, 12), 531 => to_unsigned(2049, 12), 532 => to_unsigned(3872, 12), 533 => to_unsigned(2462, 12), 534 => to_unsigned(2625, 12), 535 => to_unsigned(419, 12), 536 => to_unsigned(3193, 12), 537 => to_unsigned(3020, 12), 538 => to_unsigned(161, 12), 539 => to_unsigned(1061, 12), 540 => to_unsigned(907, 12), 541 => to_unsigned(2781, 12), 542 => to_unsigned(1116, 12), 543 => to_unsigned(803, 12), 544 => to_unsigned(2894, 12), 545 => to_unsigned(991, 12), 546 => to_unsigned(1905, 12), 547 => to_unsigned(944, 12), 548 => to_unsigned(4076, 12), 549 => to_unsigned(3170, 12), 550 => to_unsigned(2687, 12), 551 => to_unsigned(523, 12), 552 => to_unsigned(2182, 12), 553 => to_unsigned(322, 12), 554 => to_unsigned(3798, 12), 555 => to_unsigned(1182, 12), 556 => to_unsigned(2264, 12), 557 => to_unsigned(3694, 12), 558 => to_unsigned(2704, 12), 559 => to_unsigned(3154, 12), 560 => to_unsigned(1678, 12), 561 => to_unsigned(1315, 12), 562 => to_unsigned(2018, 12), 563 => to_unsigned(3202, 12), 564 => to_unsigned(2435, 12), 565 => to_unsigned(1582, 12), 566 => to_unsigned(4039, 12), 567 => to_unsigned(2305, 12), 568 => to_unsigned(83, 12), 569 => to_unsigned(67, 12), 570 => to_unsigned(1367, 12), 571 => to_unsigned(2051, 12), 572 => to_unsigned(2778, 12), 573 => to_unsigned(2403, 12), 574 => to_unsigned(3146, 12), 575 => to_unsigned(579, 12), 576 => to_unsigned(3606, 12), 577 => to_unsigned(1942, 12), 578 => to_unsigned(3265, 12), 579 => to_unsigned(3469, 12), 580 => to_unsigned(2494, 12), 581 => to_unsigned(2128, 12), 582 => to_unsigned(1165, 12), 583 => to_unsigned(2832, 12), 584 => to_unsigned(2210, 12), 585 => to_unsigned(1820, 12), 586 => to_unsigned(2649, 12), 587 => to_unsigned(2065, 12), 588 => to_unsigned(723, 12), 589 => to_unsigned(558, 12), 590 => to_unsigned(3516, 12), 591 => to_unsigned(3853, 12), 592 => to_unsigned(2125, 12), 593 => to_unsigned(416, 12), 594 => to_unsigned(1522, 12), 595 => to_unsigned(390, 12), 596 => to_unsigned(187, 12), 597 => to_unsigned(787, 12), 598 => to_unsigned(2710, 12), 599 => to_unsigned(1716, 12), 600 => to_unsigned(1539, 12), 601 => to_unsigned(1704, 12), 602 => to_unsigned(279, 12), 603 => to_unsigned(892, 12), 604 => to_unsigned(1376, 12), 605 => to_unsigned(1998, 12), 606 => to_unsigned(131, 12), 607 => to_unsigned(2986, 12), 608 => to_unsigned(914, 12), 609 => to_unsigned(3939, 12), 610 => to_unsigned(2956, 12), 611 => to_unsigned(2897, 12), 612 => to_unsigned(1387, 12), 613 => to_unsigned(4038, 12), 614 => to_unsigned(238, 12), 615 => to_unsigned(2254, 12), 616 => to_unsigned(1409, 12), 617 => to_unsigned(2206, 12), 618 => to_unsigned(1351, 12), 619 => to_unsigned(2552, 12), 620 => to_unsigned(3545, 12), 621 => to_unsigned(3261, 12), 622 => to_unsigned(98, 12), 623 => to_unsigned(608, 12), 624 => to_unsigned(1040, 12), 625 => to_unsigned(1657, 12), 626 => to_unsigned(1923, 12), 627 => to_unsigned(1202, 12), 628 => to_unsigned(2437, 12), 629 => to_unsigned(3892, 12), 630 => to_unsigned(2470, 12), 631 => to_unsigned(53, 12), 632 => to_unsigned(3183, 12), 633 => to_unsigned(2475, 12), 634 => to_unsigned(216, 12), 635 => to_unsigned(614, 12), 636 => to_unsigned(367, 12), 637 => to_unsigned(1621, 12), 638 => to_unsigned(1636, 12), 639 => to_unsigned(1001, 12), 640 => to_unsigned(855, 12), 641 => to_unsigned(2994, 12), 642 => to_unsigned(3326, 12), 643 => to_unsigned(1616, 12), 644 => to_unsigned(2880, 12), 645 => to_unsigned(1928, 12), 646 => to_unsigned(2706, 12), 647 => to_unsigned(3044, 12), 648 => to_unsigned(564, 12), 649 => to_unsigned(3492, 12), 650 => to_unsigned(934, 12), 651 => to_unsigned(725, 12), 652 => to_unsigned(3740, 12), 653 => to_unsigned(144, 12), 654 => to_unsigned(2204, 12), 655 => to_unsigned(2951, 12), 656 => to_unsigned(2175, 12), 657 => to_unsigned(863, 12), 658 => to_unsigned(190, 12), 659 => to_unsigned(89, 12), 660 => to_unsigned(1029, 12), 661 => to_unsigned(942, 12), 662 => to_unsigned(1078, 12), 663 => to_unsigned(3982, 12), 664 => to_unsigned(1498, 12), 665 => to_unsigned(2094, 12), 666 => to_unsigned(2183, 12), 667 => to_unsigned(2004, 12), 668 => to_unsigned(1489, 12), 669 => to_unsigned(780, 12), 670 => to_unsigned(3836, 12), 671 => to_unsigned(2830, 12), 672 => to_unsigned(1573, 12), 673 => to_unsigned(3629, 12), 674 => to_unsigned(1418, 12), 675 => to_unsigned(2789, 12), 676 => to_unsigned(3962, 12), 677 => to_unsigned(3376, 12), 678 => to_unsigned(1302, 12), 679 => to_unsigned(1325, 12), 680 => to_unsigned(3433, 12), 681 => to_unsigned(1001, 12), 682 => to_unsigned(1314, 12), 683 => to_unsigned(3876, 12), 684 => to_unsigned(491, 12), 685 => to_unsigned(3447, 12), 686 => to_unsigned(3839, 12), 687 => to_unsigned(2006, 12), 688 => to_unsigned(3797, 12), 689 => to_unsigned(1649, 12), 690 => to_unsigned(2410, 12), 691 => to_unsigned(844, 12), 692 => to_unsigned(2500, 12), 693 => to_unsigned(1964, 12), 694 => to_unsigned(1653, 12), 695 => to_unsigned(390, 12), 696 => to_unsigned(799, 12), 697 => to_unsigned(1528, 12), 698 => to_unsigned(1314, 12), 699 => to_unsigned(2467, 12), 700 => to_unsigned(381, 12), 701 => to_unsigned(0, 12), 702 => to_unsigned(2946, 12), 703 => to_unsigned(870, 12), 704 => to_unsigned(1386, 12), 705 => to_unsigned(2767, 12), 706 => to_unsigned(1946, 12), 707 => to_unsigned(2953, 12), 708 => to_unsigned(4035, 12), 709 => to_unsigned(3699, 12), 710 => to_unsigned(2949, 12), 711 => to_unsigned(1379, 12), 712 => to_unsigned(1578, 12), 713 => to_unsigned(3318, 12), 714 => to_unsigned(564, 12), 715 => to_unsigned(535, 12), 716 => to_unsigned(2483, 12), 717 => to_unsigned(2968, 12), 718 => to_unsigned(1662, 12), 719 => to_unsigned(3878, 12), 720 => to_unsigned(4045, 12), 721 => to_unsigned(4075, 12), 722 => to_unsigned(1184, 12), 723 => to_unsigned(3479, 12), 724 => to_unsigned(932, 12), 725 => to_unsigned(1132, 12), 726 => to_unsigned(80, 12), 727 => to_unsigned(611, 12), 728 => to_unsigned(1269, 12), 729 => to_unsigned(2281, 12), 730 => to_unsigned(1033, 12), 731 => to_unsigned(3830, 12), 732 => to_unsigned(1914, 12), 733 => to_unsigned(2983, 12), 734 => to_unsigned(1272, 12), 735 => to_unsigned(1853, 12), 736 => to_unsigned(617, 12), 737 => to_unsigned(3262, 12), 738 => to_unsigned(1181, 12), 739 => to_unsigned(3129, 12), 740 => to_unsigned(1175, 12), 741 => to_unsigned(3989, 12), 742 => to_unsigned(1407, 12), 743 => to_unsigned(1918, 12), 744 => to_unsigned(2970, 12), 745 => to_unsigned(108, 12), 746 => to_unsigned(1056, 12), 747 => to_unsigned(609, 12), 748 => to_unsigned(3826, 12), 749 => to_unsigned(1311, 12), 750 => to_unsigned(230, 12), 751 => to_unsigned(411, 12), 752 => to_unsigned(2305, 12), 753 => to_unsigned(3551, 12), 754 => to_unsigned(2266, 12), 755 => to_unsigned(447, 12), 756 => to_unsigned(1458, 12), 757 => to_unsigned(375, 12), 758 => to_unsigned(165, 12), 759 => to_unsigned(439, 12), 760 => to_unsigned(3495, 12), 761 => to_unsigned(645, 12), 762 => to_unsigned(3036, 12), 763 => to_unsigned(775, 12), 764 => to_unsigned(229, 12), 765 => to_unsigned(3671, 12), 766 => to_unsigned(1536, 12), 767 => to_unsigned(424, 12), 768 => to_unsigned(2436, 12), 769 => to_unsigned(3496, 12), 770 => to_unsigned(1081, 12), 771 => to_unsigned(2339, 12), 772 => to_unsigned(1597, 12), 773 => to_unsigned(2733, 12), 774 => to_unsigned(3644, 12), 775 => to_unsigned(2607, 12), 776 => to_unsigned(2637, 12), 777 => to_unsigned(443, 12), 778 => to_unsigned(1285, 12), 779 => to_unsigned(818, 12), 780 => to_unsigned(3272, 12), 781 => to_unsigned(3701, 12), 782 => to_unsigned(2924, 12), 783 => to_unsigned(3486, 12), 784 => to_unsigned(4012, 12), 785 => to_unsigned(1324, 12), 786 => to_unsigned(1773, 12), 787 => to_unsigned(2224, 12), 788 => to_unsigned(1366, 12), 789 => to_unsigned(1396, 12), 790 => to_unsigned(2000, 12), 791 => to_unsigned(1401, 12), 792 => to_unsigned(974, 12), 793 => to_unsigned(2565, 12), 794 => to_unsigned(3082, 12), 795 => to_unsigned(867, 12), 796 => to_unsigned(2900, 12), 797 => to_unsigned(1948, 12), 798 => to_unsigned(2438, 12), 799 => to_unsigned(948, 12), 800 => to_unsigned(828, 12), 801 => to_unsigned(3572, 12), 802 => to_unsigned(2339, 12), 803 => to_unsigned(84, 12), 804 => to_unsigned(605, 12), 805 => to_unsigned(2388, 12), 806 => to_unsigned(999, 12), 807 => to_unsigned(2075, 12), 808 => to_unsigned(3287, 12), 809 => to_unsigned(3182, 12), 810 => to_unsigned(1360, 12), 811 => to_unsigned(2590, 12), 812 => to_unsigned(1378, 12), 813 => to_unsigned(472, 12), 814 => to_unsigned(2604, 12), 815 => to_unsigned(3262, 12), 816 => to_unsigned(2148, 12), 817 => to_unsigned(174, 12), 818 => to_unsigned(4037, 12), 819 => to_unsigned(1291, 12), 820 => to_unsigned(2497, 12), 821 => to_unsigned(763, 12), 822 => to_unsigned(1050, 12), 823 => to_unsigned(510, 12), 824 => to_unsigned(2099, 12), 825 => to_unsigned(3188, 12), 826 => to_unsigned(3436, 12), 827 => to_unsigned(1299, 12), 828 => to_unsigned(3928, 12), 829 => to_unsigned(4003, 12), 830 => to_unsigned(436, 12), 831 => to_unsigned(1612, 12), 832 => to_unsigned(3423, 12), 833 => to_unsigned(1457, 12), 834 => to_unsigned(450, 12), 835 => to_unsigned(28, 12), 836 => to_unsigned(3572, 12), 837 => to_unsigned(24, 12), 838 => to_unsigned(3625, 12), 839 => to_unsigned(1192, 12), 840 => to_unsigned(1425, 12), 841 => to_unsigned(3222, 12), 842 => to_unsigned(876, 12), 843 => to_unsigned(1606, 12), 844 => to_unsigned(2549, 12), 845 => to_unsigned(2810, 12), 846 => to_unsigned(2387, 12), 847 => to_unsigned(717, 12), 848 => to_unsigned(257, 12), 849 => to_unsigned(1827, 12), 850 => to_unsigned(2267, 12), 851 => to_unsigned(67, 12), 852 => to_unsigned(4080, 12), 853 => to_unsigned(1467, 12), 854 => to_unsigned(2570, 12), 855 => to_unsigned(2836, 12), 856 => to_unsigned(1767, 12), 857 => to_unsigned(1024, 12), 858 => to_unsigned(1169, 12), 859 => to_unsigned(1215, 12), 860 => to_unsigned(3209, 12), 861 => to_unsigned(1755, 12), 862 => to_unsigned(2220, 12), 863 => to_unsigned(2144, 12), 864 => to_unsigned(1264, 12), 865 => to_unsigned(3597, 12), 866 => to_unsigned(2370, 12), 867 => to_unsigned(3311, 12), 868 => to_unsigned(365, 12), 869 => to_unsigned(3244, 12), 870 => to_unsigned(134, 12), 871 => to_unsigned(1305, 12), 872 => to_unsigned(35, 12), 873 => to_unsigned(3831, 12), 874 => to_unsigned(649, 12), 875 => to_unsigned(1824, 12), 876 => to_unsigned(2127, 12), 877 => to_unsigned(1273, 12), 878 => to_unsigned(618, 12), 879 => to_unsigned(2870, 12), 880 => to_unsigned(921, 12), 881 => to_unsigned(203, 12), 882 => to_unsigned(1316, 12), 883 => to_unsigned(1216, 12), 884 => to_unsigned(1247, 12), 885 => to_unsigned(2809, 12), 886 => to_unsigned(237, 12), 887 => to_unsigned(621, 12), 888 => to_unsigned(2807, 12), 889 => to_unsigned(2787, 12), 890 => to_unsigned(1982, 12), 891 => to_unsigned(3729, 12), 892 => to_unsigned(1354, 12), 893 => to_unsigned(2470, 12), 894 => to_unsigned(714, 12), 895 => to_unsigned(2294, 12), 896 => to_unsigned(3335, 12), 897 => to_unsigned(573, 12), 898 => to_unsigned(874, 12), 899 => to_unsigned(2346, 12), 900 => to_unsigned(1407, 12), 901 => to_unsigned(1766, 12), 902 => to_unsigned(26, 12), 903 => to_unsigned(1537, 12), 904 => to_unsigned(657, 12), 905 => to_unsigned(1393, 12), 906 => to_unsigned(1484, 12), 907 => to_unsigned(2138, 12), 908 => to_unsigned(3326, 12), 909 => to_unsigned(1503, 12), 910 => to_unsigned(3452, 12), 911 => to_unsigned(811, 12), 912 => to_unsigned(1630, 12), 913 => to_unsigned(3870, 12), 914 => to_unsigned(3574, 12), 915 => to_unsigned(3961, 12), 916 => to_unsigned(1229, 12), 917 => to_unsigned(2968, 12), 918 => to_unsigned(2012, 12), 919 => to_unsigned(3782, 12), 920 => to_unsigned(3135, 12), 921 => to_unsigned(212, 12), 922 => to_unsigned(3049, 12), 923 => to_unsigned(3044, 12), 924 => to_unsigned(3338, 12), 925 => to_unsigned(2279, 12), 926 => to_unsigned(3715, 12), 927 => to_unsigned(1988, 12), 928 => to_unsigned(1366, 12), 929 => to_unsigned(1563, 12), 930 => to_unsigned(592, 12), 931 => to_unsigned(540, 12), 932 => to_unsigned(3559, 12), 933 => to_unsigned(998, 12), 934 => to_unsigned(1874, 12), 935 => to_unsigned(1587, 12), 936 => to_unsigned(2700, 12), 937 => to_unsigned(216, 12), 938 => to_unsigned(1662, 12), 939 => to_unsigned(1957, 12), 940 => to_unsigned(391, 12), 941 => to_unsigned(51, 12), 942 => to_unsigned(1100, 12), 943 => to_unsigned(3905, 12), 944 => to_unsigned(3145, 12), 945 => to_unsigned(3633, 12), 946 => to_unsigned(1307, 12), 947 => to_unsigned(3308, 12), 948 => to_unsigned(1123, 12), 949 => to_unsigned(3176, 12), 950 => to_unsigned(3144, 12), 951 => to_unsigned(1714, 12), 952 => to_unsigned(2481, 12), 953 => to_unsigned(3015, 12), 954 => to_unsigned(3267, 12), 955 => to_unsigned(3194, 12), 956 => to_unsigned(1994, 12), 957 => to_unsigned(470, 12), 958 => to_unsigned(3045, 12), 959 => to_unsigned(1775, 12), 960 => to_unsigned(2702, 12), 961 => to_unsigned(3939, 12), 962 => to_unsigned(4050, 12), 963 => to_unsigned(3123, 12), 964 => to_unsigned(2549, 12), 965 => to_unsigned(3789, 12), 966 => to_unsigned(2434, 12), 967 => to_unsigned(1362, 12), 968 => to_unsigned(838, 12), 969 => to_unsigned(2536, 12), 970 => to_unsigned(2951, 12), 971 => to_unsigned(854, 12), 972 => to_unsigned(1832, 12), 973 => to_unsigned(2703, 12), 974 => to_unsigned(3051, 12), 975 => to_unsigned(1563, 12), 976 => to_unsigned(3829, 12), 977 => to_unsigned(2025, 12), 978 => to_unsigned(2950, 12), 979 => to_unsigned(3832, 12), 980 => to_unsigned(488, 12), 981 => to_unsigned(1731, 12), 982 => to_unsigned(508, 12), 983 => to_unsigned(1125, 12), 984 => to_unsigned(2894, 12), 985 => to_unsigned(3165, 12), 986 => to_unsigned(3360, 12), 987 => to_unsigned(2839, 12), 988 => to_unsigned(528, 12), 989 => to_unsigned(1328, 12), 990 => to_unsigned(857, 12), 991 => to_unsigned(2501, 12), 992 => to_unsigned(1704, 12), 993 => to_unsigned(167, 12), 994 => to_unsigned(2430, 12), 995 => to_unsigned(3874, 12), 996 => to_unsigned(845, 12), 997 => to_unsigned(1319, 12), 998 => to_unsigned(2515, 12), 999 => to_unsigned(2903, 12), 1000 => to_unsigned(1069, 12), 1001 => to_unsigned(2554, 12), 1002 => to_unsigned(564, 12), 1003 => to_unsigned(2447, 12), 1004 => to_unsigned(196, 12), 1005 => to_unsigned(2207, 12), 1006 => to_unsigned(1915, 12), 1007 => to_unsigned(578, 12), 1008 => to_unsigned(2082, 12), 1009 => to_unsigned(520, 12), 1010 => to_unsigned(1238, 12), 1011 => to_unsigned(2990, 12), 1012 => to_unsigned(993, 12), 1013 => to_unsigned(1903, 12), 1014 => to_unsigned(1779, 12), 1015 => to_unsigned(3400, 12), 1016 => to_unsigned(241, 12), 1017 => to_unsigned(181, 12), 1018 => to_unsigned(1619, 12), 1019 => to_unsigned(3449, 12), 1020 => to_unsigned(2973, 12), 1021 => to_unsigned(2303, 12), 1022 => to_unsigned(2312, 12), 1023 => to_unsigned(1934, 12), 1024 => to_unsigned(3557, 12), 1025 => to_unsigned(3285, 12), 1026 => to_unsigned(918, 12), 1027 => to_unsigned(2531, 12), 1028 => to_unsigned(3556, 12), 1029 => to_unsigned(3542, 12), 1030 => to_unsigned(197, 12), 1031 => to_unsigned(2605, 12), 1032 => to_unsigned(3610, 12), 1033 => to_unsigned(3747, 12), 1034 => to_unsigned(235, 12), 1035 => to_unsigned(1056, 12), 1036 => to_unsigned(1108, 12), 1037 => to_unsigned(2631, 12), 1038 => to_unsigned(3033, 12), 1039 => to_unsigned(2373, 12), 1040 => to_unsigned(2607, 12), 1041 => to_unsigned(502, 12), 1042 => to_unsigned(3801, 12), 1043 => to_unsigned(500, 12), 1044 => to_unsigned(652, 12), 1045 => to_unsigned(553, 12), 1046 => to_unsigned(1544, 12), 1047 => to_unsigned(3568, 12), 1048 => to_unsigned(3144, 12), 1049 => to_unsigned(2394, 12), 1050 => to_unsigned(3118, 12), 1051 => to_unsigned(1758, 12), 1052 => to_unsigned(3350, 12), 1053 => to_unsigned(4054, 12), 1054 => to_unsigned(513, 12), 1055 => to_unsigned(1652, 12), 1056 => to_unsigned(2036, 12), 1057 => to_unsigned(714, 12), 1058 => to_unsigned(2226, 12), 1059 => to_unsigned(840, 12), 1060 => to_unsigned(497, 12), 1061 => to_unsigned(3019, 12), 1062 => to_unsigned(1621, 12), 1063 => to_unsigned(259, 12), 1064 => to_unsigned(488, 12), 1065 => to_unsigned(1597, 12), 1066 => to_unsigned(2731, 12), 1067 => to_unsigned(1827, 12), 1068 => to_unsigned(3424, 12), 1069 => to_unsigned(3303, 12), 1070 => to_unsigned(3459, 12), 1071 => to_unsigned(1771, 12), 1072 => to_unsigned(2703, 12), 1073 => to_unsigned(2665, 12), 1074 => to_unsigned(260, 12), 1075 => to_unsigned(2437, 12), 1076 => to_unsigned(1838, 12), 1077 => to_unsigned(2061, 12), 1078 => to_unsigned(3289, 12), 1079 => to_unsigned(2682, 12), 1080 => to_unsigned(2002, 12), 1081 => to_unsigned(3623, 12), 1082 => to_unsigned(1221, 12), 1083 => to_unsigned(1550, 12), 1084 => to_unsigned(715, 12), 1085 => to_unsigned(826, 12), 1086 => to_unsigned(4012, 12), 1087 => to_unsigned(586, 12), 1088 => to_unsigned(555, 12), 1089 => to_unsigned(1359, 12), 1090 => to_unsigned(3727, 12), 1091 => to_unsigned(3095, 12), 1092 => to_unsigned(3300, 12), 1093 => to_unsigned(3519, 12), 1094 => to_unsigned(528, 12), 1095 => to_unsigned(3134, 12), 1096 => to_unsigned(3921, 12), 1097 => to_unsigned(3496, 12), 1098 => to_unsigned(865, 12), 1099 => to_unsigned(2997, 12), 1100 => to_unsigned(3833, 12), 1101 => to_unsigned(3248, 12), 1102 => to_unsigned(3578, 12), 1103 => to_unsigned(1645, 12), 1104 => to_unsigned(1647, 12), 1105 => to_unsigned(180, 12), 1106 => to_unsigned(3087, 12), 1107 => to_unsigned(1918, 12), 1108 => to_unsigned(23, 12), 1109 => to_unsigned(4046, 12), 1110 => to_unsigned(1329, 12), 1111 => to_unsigned(2568, 12), 1112 => to_unsigned(2336, 12), 1113 => to_unsigned(929, 12), 1114 => to_unsigned(2427, 12), 1115 => to_unsigned(657, 12), 1116 => to_unsigned(1923, 12), 1117 => to_unsigned(2453, 12), 1118 => to_unsigned(56, 12), 1119 => to_unsigned(3147, 12), 1120 => to_unsigned(2012, 12), 1121 => to_unsigned(3574, 12), 1122 => to_unsigned(2024, 12), 1123 => to_unsigned(2720, 12), 1124 => to_unsigned(1305, 12), 1125 => to_unsigned(2906, 12), 1126 => to_unsigned(3037, 12), 1127 => to_unsigned(308, 12), 1128 => to_unsigned(1798, 12), 1129 => to_unsigned(1247, 12), 1130 => to_unsigned(3919, 12), 1131 => to_unsigned(521, 12), 1132 => to_unsigned(2905, 12), 1133 => to_unsigned(1761, 12), 1134 => to_unsigned(3919, 12), 1135 => to_unsigned(2267, 12), 1136 => to_unsigned(2795, 12), 1137 => to_unsigned(246, 12), 1138 => to_unsigned(2718, 12), 1139 => to_unsigned(3832, 12), 1140 => to_unsigned(1918, 12), 1141 => to_unsigned(2786, 12), 1142 => to_unsigned(1896, 12), 1143 => to_unsigned(2931, 12), 1144 => to_unsigned(706, 12), 1145 => to_unsigned(270, 12), 1146 => to_unsigned(2528, 12), 1147 => to_unsigned(1131, 12), 1148 => to_unsigned(1936, 12), 1149 => to_unsigned(1423, 12), 1150 => to_unsigned(3279, 12), 1151 => to_unsigned(3502, 12), 1152 => to_unsigned(1550, 12), 1153 => to_unsigned(2174, 12), 1154 => to_unsigned(1511, 12), 1155 => to_unsigned(3037, 12), 1156 => to_unsigned(3508, 12), 1157 => to_unsigned(2453, 12), 1158 => to_unsigned(359, 12), 1159 => to_unsigned(25, 12), 1160 => to_unsigned(1612, 12), 1161 => to_unsigned(2507, 12), 1162 => to_unsigned(3617, 12), 1163 => to_unsigned(576, 12), 1164 => to_unsigned(231, 12), 1165 => to_unsigned(1454, 12), 1166 => to_unsigned(3371, 12), 1167 => to_unsigned(611, 12), 1168 => to_unsigned(2068, 12), 1169 => to_unsigned(2088, 12), 1170 => to_unsigned(2588, 12), 1171 => to_unsigned(661, 12), 1172 => to_unsigned(1038, 12), 1173 => to_unsigned(850, 12), 1174 => to_unsigned(795, 12), 1175 => to_unsigned(394, 12), 1176 => to_unsigned(1168, 12), 1177 => to_unsigned(3051, 12), 1178 => to_unsigned(3340, 12), 1179 => to_unsigned(3759, 12), 1180 => to_unsigned(1204, 12), 1181 => to_unsigned(2604, 12), 1182 => to_unsigned(1457, 12), 1183 => to_unsigned(3862, 12), 1184 => to_unsigned(627, 12), 1185 => to_unsigned(1344, 12), 1186 => to_unsigned(2826, 12), 1187 => to_unsigned(2969, 12), 1188 => to_unsigned(2187, 12), 1189 => to_unsigned(3455, 12), 1190 => to_unsigned(1999, 12), 1191 => to_unsigned(1695, 12), 1192 => to_unsigned(2243, 12), 1193 => to_unsigned(994, 12), 1194 => to_unsigned(998, 12), 1195 => to_unsigned(2382, 12), 1196 => to_unsigned(4081, 12), 1197 => to_unsigned(1886, 12), 1198 => to_unsigned(2884, 12), 1199 => to_unsigned(936, 12), 1200 => to_unsigned(281, 12), 1201 => to_unsigned(1439, 12), 1202 => to_unsigned(2982, 12), 1203 => to_unsigned(2182, 12), 1204 => to_unsigned(3865, 12), 1205 => to_unsigned(2603, 12), 1206 => to_unsigned(3859, 12), 1207 => to_unsigned(1314, 12), 1208 => to_unsigned(1079, 12), 1209 => to_unsigned(277, 12), 1210 => to_unsigned(487, 12), 1211 => to_unsigned(2126, 12), 1212 => to_unsigned(3823, 12), 1213 => to_unsigned(310, 12), 1214 => to_unsigned(1297, 12), 1215 => to_unsigned(3828, 12), 1216 => to_unsigned(1817, 12), 1217 => to_unsigned(670, 12), 1218 => to_unsigned(2841, 12), 1219 => to_unsigned(3055, 12), 1220 => to_unsigned(693, 12), 1221 => to_unsigned(3317, 12), 1222 => to_unsigned(3263, 12), 1223 => to_unsigned(1370, 12), 1224 => to_unsigned(2936, 12), 1225 => to_unsigned(3590, 12), 1226 => to_unsigned(2049, 12), 1227 => to_unsigned(2410, 12), 1228 => to_unsigned(2660, 12), 1229 => to_unsigned(3525, 12), 1230 => to_unsigned(3447, 12), 1231 => to_unsigned(1453, 12), 1232 => to_unsigned(3123, 12), 1233 => to_unsigned(1622, 12), 1234 => to_unsigned(1346, 12), 1235 => to_unsigned(1041, 12), 1236 => to_unsigned(3510, 12), 1237 => to_unsigned(3481, 12), 1238 => to_unsigned(1230, 12), 1239 => to_unsigned(2990, 12), 1240 => to_unsigned(1147, 12), 1241 => to_unsigned(1331, 12), 1242 => to_unsigned(95, 12), 1243 => to_unsigned(483, 12), 1244 => to_unsigned(3568, 12), 1245 => to_unsigned(2036, 12), 1246 => to_unsigned(3630, 12), 1247 => to_unsigned(1952, 12), 1248 => to_unsigned(355, 12), 1249 => to_unsigned(580, 12), 1250 => to_unsigned(1481, 12), 1251 => to_unsigned(1615, 12), 1252 => to_unsigned(3934, 12), 1253 => to_unsigned(1886, 12), 1254 => to_unsigned(1011, 12), 1255 => to_unsigned(927, 12), 1256 => to_unsigned(430, 12), 1257 => to_unsigned(3269, 12), 1258 => to_unsigned(877, 12), 1259 => to_unsigned(808, 12), 1260 => to_unsigned(839, 12), 1261 => to_unsigned(222, 12), 1262 => to_unsigned(67, 12), 1263 => to_unsigned(3408, 12), 1264 => to_unsigned(155, 12), 1265 => to_unsigned(3624, 12), 1266 => to_unsigned(1121, 12), 1267 => to_unsigned(2301, 12), 1268 => to_unsigned(2801, 12), 1269 => to_unsigned(1907, 12), 1270 => to_unsigned(1574, 12), 1271 => to_unsigned(1167, 12), 1272 => to_unsigned(2593, 12), 1273 => to_unsigned(461, 12), 1274 => to_unsigned(165, 12), 1275 => to_unsigned(1843, 12), 1276 => to_unsigned(3783, 12), 1277 => to_unsigned(1969, 12), 1278 => to_unsigned(1624, 12), 1279 => to_unsigned(132, 12), 1280 => to_unsigned(3264, 12), 1281 => to_unsigned(2892, 12), 1282 => to_unsigned(247, 12), 1283 => to_unsigned(2699, 12), 1284 => to_unsigned(1007, 12), 1285 => to_unsigned(392, 12), 1286 => to_unsigned(1375, 12), 1287 => to_unsigned(3435, 12), 1288 => to_unsigned(3951, 12), 1289 => to_unsigned(3431, 12), 1290 => to_unsigned(1632, 12), 1291 => to_unsigned(3624, 12), 1292 => to_unsigned(2085, 12), 1293 => to_unsigned(2027, 12), 1294 => to_unsigned(252, 12), 1295 => to_unsigned(613, 12), 1296 => to_unsigned(3469, 12), 1297 => to_unsigned(1039, 12), 1298 => to_unsigned(3321, 12), 1299 => to_unsigned(1262, 12), 1300 => to_unsigned(627, 12), 1301 => to_unsigned(442, 12), 1302 => to_unsigned(347, 12), 1303 => to_unsigned(246, 12), 1304 => to_unsigned(3111, 12), 1305 => to_unsigned(785, 12), 1306 => to_unsigned(1622, 12), 1307 => to_unsigned(3826, 12), 1308 => to_unsigned(139, 12), 1309 => to_unsigned(2415, 12), 1310 => to_unsigned(1498, 12), 1311 => to_unsigned(3003, 12), 1312 => to_unsigned(2067, 12), 1313 => to_unsigned(1452, 12), 1314 => to_unsigned(19, 12), 1315 => to_unsigned(2485, 12), 1316 => to_unsigned(460, 12), 1317 => to_unsigned(118, 12), 1318 => to_unsigned(851, 12), 1319 => to_unsigned(2151, 12), 1320 => to_unsigned(3958, 12), 1321 => to_unsigned(3241, 12), 1322 => to_unsigned(3122, 12), 1323 => to_unsigned(2924, 12), 1324 => to_unsigned(1074, 12), 1325 => to_unsigned(3748, 12), 1326 => to_unsigned(939, 12), 1327 => to_unsigned(4066, 12), 1328 => to_unsigned(2218, 12), 1329 => to_unsigned(2153, 12), 1330 => to_unsigned(1972, 12), 1331 => to_unsigned(130, 12), 1332 => to_unsigned(2301, 12), 1333 => to_unsigned(2564, 12), 1334 => to_unsigned(1815, 12), 1335 => to_unsigned(2597, 12), 1336 => to_unsigned(2926, 12), 1337 => to_unsigned(887, 12), 1338 => to_unsigned(205, 12), 1339 => to_unsigned(2166, 12), 1340 => to_unsigned(3741, 12), 1341 => to_unsigned(3731, 12), 1342 => to_unsigned(1061, 12), 1343 => to_unsigned(3678, 12), 1344 => to_unsigned(3502, 12), 1345 => to_unsigned(3111, 12), 1346 => to_unsigned(496, 12), 1347 => to_unsigned(2582, 12), 1348 => to_unsigned(2618, 12), 1349 => to_unsigned(2144, 12), 1350 => to_unsigned(2320, 12), 1351 => to_unsigned(2134, 12), 1352 => to_unsigned(1494, 12), 1353 => to_unsigned(361, 12), 1354 => to_unsigned(1419, 12), 1355 => to_unsigned(435, 12), 1356 => to_unsigned(2352, 12), 1357 => to_unsigned(2803, 12), 1358 => to_unsigned(1830, 12), 1359 => to_unsigned(1944, 12), 1360 => to_unsigned(1770, 12), 1361 => to_unsigned(1516, 12), 1362 => to_unsigned(3083, 12), 1363 => to_unsigned(2936, 12), 1364 => to_unsigned(2864, 12), 1365 => to_unsigned(3583, 12), 1366 => to_unsigned(1460, 12), 1367 => to_unsigned(510, 12), 1368 => to_unsigned(1395, 12), 1369 => to_unsigned(1324, 12), 1370 => to_unsigned(1573, 12), 1371 => to_unsigned(976, 12), 1372 => to_unsigned(2840, 12), 1373 => to_unsigned(1010, 12), 1374 => to_unsigned(704, 12), 1375 => to_unsigned(1670, 12), 1376 => to_unsigned(2766, 12), 1377 => to_unsigned(2022, 12), 1378 => to_unsigned(4073, 12), 1379 => to_unsigned(2220, 12), 1380 => to_unsigned(476, 12), 1381 => to_unsigned(3625, 12), 1382 => to_unsigned(88, 12), 1383 => to_unsigned(2233, 12), 1384 => to_unsigned(866, 12), 1385 => to_unsigned(1076, 12), 1386 => to_unsigned(2767, 12), 1387 => to_unsigned(1436, 12), 1388 => to_unsigned(3206, 12), 1389 => to_unsigned(2840, 12), 1390 => to_unsigned(790, 12), 1391 => to_unsigned(386, 12), 1392 => to_unsigned(2440, 12), 1393 => to_unsigned(2731, 12), 1394 => to_unsigned(1188, 12), 1395 => to_unsigned(1260, 12), 1396 => to_unsigned(692, 12), 1397 => to_unsigned(3463, 12), 1398 => to_unsigned(2916, 12), 1399 => to_unsigned(2351, 12), 1400 => to_unsigned(1219, 12), 1401 => to_unsigned(1058, 12), 1402 => to_unsigned(1608, 12), 1403 => to_unsigned(1732, 12), 1404 => to_unsigned(244, 12), 1405 => to_unsigned(2712, 12), 1406 => to_unsigned(3141, 12), 1407 => to_unsigned(2765, 12), 1408 => to_unsigned(805, 12), 1409 => to_unsigned(2084, 12), 1410 => to_unsigned(374, 12), 1411 => to_unsigned(3962, 12), 1412 => to_unsigned(2633, 12), 1413 => to_unsigned(2758, 12), 1414 => to_unsigned(2165, 12), 1415 => to_unsigned(2899, 12), 1416 => to_unsigned(1590, 12), 1417 => to_unsigned(3876, 12), 1418 => to_unsigned(3936, 12), 1419 => to_unsigned(3258, 12), 1420 => to_unsigned(2462, 12), 1421 => to_unsigned(2286, 12), 1422 => to_unsigned(775, 12), 1423 => to_unsigned(1479, 12), 1424 => to_unsigned(2797, 12), 1425 => to_unsigned(2290, 12), 1426 => to_unsigned(1168, 12), 1427 => to_unsigned(136, 12), 1428 => to_unsigned(1519, 12), 1429 => to_unsigned(3909, 12), 1430 => to_unsigned(699, 12), 1431 => to_unsigned(885, 12), 1432 => to_unsigned(1919, 12), 1433 => to_unsigned(2743, 12), 1434 => to_unsigned(2806, 12), 1435 => to_unsigned(1364, 12), 1436 => to_unsigned(996, 12), 1437 => to_unsigned(654, 12), 1438 => to_unsigned(3826, 12), 1439 => to_unsigned(643, 12), 1440 => to_unsigned(405, 12), 1441 => to_unsigned(391, 12), 1442 => to_unsigned(623, 12), 1443 => to_unsigned(1712, 12), 1444 => to_unsigned(258, 12), 1445 => to_unsigned(745, 12), 1446 => to_unsigned(165, 12), 1447 => to_unsigned(1268, 12), 1448 => to_unsigned(734, 12), 1449 => to_unsigned(3605, 12), 1450 => to_unsigned(628, 12), 1451 => to_unsigned(3267, 12), 1452 => to_unsigned(1380, 12), 1453 => to_unsigned(2639, 12), 1454 => to_unsigned(1469, 12), 1455 => to_unsigned(2971, 12), 1456 => to_unsigned(2030, 12), 1457 => to_unsigned(1720, 12), 1458 => to_unsigned(2311, 12), 1459 => to_unsigned(3173, 12), 1460 => to_unsigned(2743, 12), 1461 => to_unsigned(3276, 12), 1462 => to_unsigned(1318, 12), 1463 => to_unsigned(2001, 12), 1464 => to_unsigned(2820, 12), 1465 => to_unsigned(3662, 12), 1466 => to_unsigned(3374, 12), 1467 => to_unsigned(1799, 12), 1468 => to_unsigned(201, 12), 1469 => to_unsigned(513, 12), 1470 => to_unsigned(276, 12), 1471 => to_unsigned(630, 12), 1472 => to_unsigned(388, 12), 1473 => to_unsigned(3045, 12), 1474 => to_unsigned(1344, 12), 1475 => to_unsigned(2012, 12), 1476 => to_unsigned(1118, 12), 1477 => to_unsigned(3751, 12), 1478 => to_unsigned(670, 12), 1479 => to_unsigned(695, 12), 1480 => to_unsigned(2988, 12), 1481 => to_unsigned(3689, 12), 1482 => to_unsigned(2610, 12), 1483 => to_unsigned(2666, 12), 1484 => to_unsigned(2276, 12), 1485 => to_unsigned(3096, 12), 1486 => to_unsigned(2389, 12), 1487 => to_unsigned(1297, 12), 1488 => to_unsigned(1095, 12), 1489 => to_unsigned(2202, 12), 1490 => to_unsigned(3234, 12), 1491 => to_unsigned(1019, 12), 1492 => to_unsigned(3813, 12), 1493 => to_unsigned(2408, 12), 1494 => to_unsigned(1339, 12), 1495 => to_unsigned(4071, 12), 1496 => to_unsigned(948, 12), 1497 => to_unsigned(2755, 12), 1498 => to_unsigned(2800, 12), 1499 => to_unsigned(3095, 12), 1500 => to_unsigned(1529, 12), 1501 => to_unsigned(2121, 12), 1502 => to_unsigned(356, 12), 1503 => to_unsigned(1262, 12), 1504 => to_unsigned(4077, 12), 1505 => to_unsigned(101, 12), 1506 => to_unsigned(2782, 12), 1507 => to_unsigned(405, 12), 1508 => to_unsigned(1443, 12), 1509 => to_unsigned(1796, 12), 1510 => to_unsigned(3155, 12), 1511 => to_unsigned(3398, 12), 1512 => to_unsigned(2102, 12), 1513 => to_unsigned(890, 12), 1514 => to_unsigned(792, 12), 1515 => to_unsigned(3300, 12), 1516 => to_unsigned(457, 12), 1517 => to_unsigned(3431, 12), 1518 => to_unsigned(2661, 12), 1519 => to_unsigned(63, 12), 1520 => to_unsigned(1800, 12), 1521 => to_unsigned(1248, 12), 1522 => to_unsigned(1651, 12), 1523 => to_unsigned(4050, 12), 1524 => to_unsigned(1239, 12), 1525 => to_unsigned(1038, 12), 1526 => to_unsigned(3977, 12), 1527 => to_unsigned(3007, 12), 1528 => to_unsigned(168, 12), 1529 => to_unsigned(121, 12), 1530 => to_unsigned(1901, 12), 1531 => to_unsigned(482, 12), 1532 => to_unsigned(3843, 12), 1533 => to_unsigned(1896, 12), 1534 => to_unsigned(3076, 12), 1535 => to_unsigned(3832, 12), 1536 => to_unsigned(3664, 12), 1537 => to_unsigned(2252, 12), 1538 => to_unsigned(3972, 12), 1539 => to_unsigned(2809, 12), 1540 => to_unsigned(3167, 12), 1541 => to_unsigned(1056, 12), 1542 => to_unsigned(1231, 12), 1543 => to_unsigned(2332, 12), 1544 => to_unsigned(2261, 12), 1545 => to_unsigned(1973, 12), 1546 => to_unsigned(3444, 12), 1547 => to_unsigned(717, 12), 1548 => to_unsigned(552, 12), 1549 => to_unsigned(819, 12), 1550 => to_unsigned(4083, 12), 1551 => to_unsigned(2268, 12), 1552 => to_unsigned(4032, 12), 1553 => to_unsigned(3785, 12), 1554 => to_unsigned(13, 12), 1555 => to_unsigned(602, 12), 1556 => to_unsigned(3659, 12), 1557 => to_unsigned(3500, 12), 1558 => to_unsigned(3849, 12), 1559 => to_unsigned(634, 12), 1560 => to_unsigned(3222, 12), 1561 => to_unsigned(2329, 12), 1562 => to_unsigned(3392, 12), 1563 => to_unsigned(2486, 12), 1564 => to_unsigned(152, 12), 1565 => to_unsigned(1732, 12), 1566 => to_unsigned(3247, 12), 1567 => to_unsigned(3057, 12), 1568 => to_unsigned(1641, 12), 1569 => to_unsigned(3988, 12), 1570 => to_unsigned(140, 12), 1571 => to_unsigned(884, 12), 1572 => to_unsigned(276, 12), 1573 => to_unsigned(2909, 12), 1574 => to_unsigned(2250, 12), 1575 => to_unsigned(971, 12), 1576 => to_unsigned(2005, 12), 1577 => to_unsigned(3865, 12), 1578 => to_unsigned(2654, 12), 1579 => to_unsigned(1447, 12), 1580 => to_unsigned(280, 12), 1581 => to_unsigned(981, 12), 1582 => to_unsigned(1353, 12), 1583 => to_unsigned(2598, 12), 1584 => to_unsigned(2084, 12), 1585 => to_unsigned(989, 12), 1586 => to_unsigned(3064, 12), 1587 => to_unsigned(1681, 12), 1588 => to_unsigned(3825, 12), 1589 => to_unsigned(1983, 12), 1590 => to_unsigned(2473, 12), 1591 => to_unsigned(486, 12), 1592 => to_unsigned(866, 12), 1593 => to_unsigned(3398, 12), 1594 => to_unsigned(956, 12), 1595 => to_unsigned(3020, 12), 1596 => to_unsigned(2393, 12), 1597 => to_unsigned(206, 12), 1598 => to_unsigned(3084, 12), 1599 => to_unsigned(2323, 12), 1600 => to_unsigned(3398, 12), 1601 => to_unsigned(1589, 12), 1602 => to_unsigned(1801, 12), 1603 => to_unsigned(3957, 12), 1604 => to_unsigned(3881, 12), 1605 => to_unsigned(2527, 12), 1606 => to_unsigned(2996, 12), 1607 => to_unsigned(3539, 12), 1608 => to_unsigned(3645, 12), 1609 => to_unsigned(2163, 12), 1610 => to_unsigned(3051, 12), 1611 => to_unsigned(2189, 12), 1612 => to_unsigned(1060, 12), 1613 => to_unsigned(2878, 12), 1614 => to_unsigned(1686, 12), 1615 => to_unsigned(1676, 12), 1616 => to_unsigned(2627, 12), 1617 => to_unsigned(1999, 12), 1618 => to_unsigned(2795, 12), 1619 => to_unsigned(3459, 12), 1620 => to_unsigned(1467, 12), 1621 => to_unsigned(2978, 12), 1622 => to_unsigned(1126, 12), 1623 => to_unsigned(291, 12), 1624 => to_unsigned(2950, 12), 1625 => to_unsigned(2699, 12), 1626 => to_unsigned(2877, 12), 1627 => to_unsigned(3010, 12), 1628 => to_unsigned(1371, 12), 1629 => to_unsigned(3147, 12), 1630 => to_unsigned(1978, 12), 1631 => to_unsigned(1222, 12), 1632 => to_unsigned(2616, 12), 1633 => to_unsigned(2527, 12), 1634 => to_unsigned(1870, 12), 1635 => to_unsigned(408, 12), 1636 => to_unsigned(1052, 12), 1637 => to_unsigned(2922, 12), 1638 => to_unsigned(4009, 12), 1639 => to_unsigned(1550, 12), 1640 => to_unsigned(2340, 12), 1641 => to_unsigned(1875, 12), 1642 => to_unsigned(3761, 12), 1643 => to_unsigned(2345, 12), 1644 => to_unsigned(2962, 12), 1645 => to_unsigned(1464, 12), 1646 => to_unsigned(567, 12), 1647 => to_unsigned(1266, 12), 1648 => to_unsigned(2542, 12), 1649 => to_unsigned(692, 12), 1650 => to_unsigned(747, 12), 1651 => to_unsigned(2481, 12), 1652 => to_unsigned(2842, 12), 1653 => to_unsigned(1571, 12), 1654 => to_unsigned(881, 12), 1655 => to_unsigned(3699, 12), 1656 => to_unsigned(3701, 12), 1657 => to_unsigned(2257, 12), 1658 => to_unsigned(3064, 12), 1659 => to_unsigned(3974, 12), 1660 => to_unsigned(836, 12), 1661 => to_unsigned(756, 12), 1662 => to_unsigned(250, 12), 1663 => to_unsigned(2618, 12), 1664 => to_unsigned(3813, 12), 1665 => to_unsigned(2769, 12), 1666 => to_unsigned(38, 12), 1667 => to_unsigned(1566, 12), 1668 => to_unsigned(695, 12), 1669 => to_unsigned(3747, 12), 1670 => to_unsigned(3024, 12), 1671 => to_unsigned(1496, 12), 1672 => to_unsigned(1453, 12), 1673 => to_unsigned(5, 12), 1674 => to_unsigned(4050, 12), 1675 => to_unsigned(2018, 12), 1676 => to_unsigned(815, 12), 1677 => to_unsigned(2670, 12), 1678 => to_unsigned(1005, 12), 1679 => to_unsigned(2492, 12), 1680 => to_unsigned(1623, 12), 1681 => to_unsigned(987, 12), 1682 => to_unsigned(1728, 12), 1683 => to_unsigned(3060, 12), 1684 => to_unsigned(3912, 12), 1685 => to_unsigned(549, 12), 1686 => to_unsigned(1998, 12), 1687 => to_unsigned(2076, 12), 1688 => to_unsigned(658, 12), 1689 => to_unsigned(1862, 12), 1690 => to_unsigned(2312, 12), 1691 => to_unsigned(612, 12), 1692 => to_unsigned(3430, 12), 1693 => to_unsigned(2114, 12), 1694 => to_unsigned(1507, 12), 1695 => to_unsigned(462, 12), 1696 => to_unsigned(55, 12), 1697 => to_unsigned(1793, 12), 1698 => to_unsigned(2237, 12), 1699 => to_unsigned(2707, 12), 1700 => to_unsigned(3255, 12), 1701 => to_unsigned(754, 12), 1702 => to_unsigned(1393, 12), 1703 => to_unsigned(3770, 12), 1704 => to_unsigned(2279, 12), 1705 => to_unsigned(2912, 12), 1706 => to_unsigned(3530, 12), 1707 => to_unsigned(3599, 12), 1708 => to_unsigned(1040, 12), 1709 => to_unsigned(1437, 12), 1710 => to_unsigned(1181, 12), 1711 => to_unsigned(2091, 12), 1712 => to_unsigned(1812, 12), 1713 => to_unsigned(3513, 12), 1714 => to_unsigned(3933, 12), 1715 => to_unsigned(215, 12), 1716 => to_unsigned(54, 12), 1717 => to_unsigned(1197, 12), 1718 => to_unsigned(1062, 12), 1719 => to_unsigned(3187, 12), 1720 => to_unsigned(2342, 12), 1721 => to_unsigned(1886, 12), 1722 => to_unsigned(1068, 12), 1723 => to_unsigned(1302, 12), 1724 => to_unsigned(3526, 12), 1725 => to_unsigned(3059, 12), 1726 => to_unsigned(3854, 12), 1727 => to_unsigned(2133, 12), 1728 => to_unsigned(3141, 12), 1729 => to_unsigned(350, 12), 1730 => to_unsigned(2392, 12), 1731 => to_unsigned(498, 12), 1732 => to_unsigned(199, 12), 1733 => to_unsigned(1216, 12), 1734 => to_unsigned(1148, 12), 1735 => to_unsigned(2809, 12), 1736 => to_unsigned(1840, 12), 1737 => to_unsigned(571, 12), 1738 => to_unsigned(63, 12), 1739 => to_unsigned(2028, 12), 1740 => to_unsigned(2837, 12), 1741 => to_unsigned(2222, 12), 1742 => to_unsigned(2554, 12), 1743 => to_unsigned(3409, 12), 1744 => to_unsigned(1491, 12), 1745 => to_unsigned(2831, 12), 1746 => to_unsigned(2565, 12), 1747 => to_unsigned(3752, 12), 1748 => to_unsigned(286, 12), 1749 => to_unsigned(177, 12), 1750 => to_unsigned(358, 12), 1751 => to_unsigned(3629, 12), 1752 => to_unsigned(162, 12), 1753 => to_unsigned(709, 12), 1754 => to_unsigned(728, 12), 1755 => to_unsigned(4053, 12), 1756 => to_unsigned(2370, 12), 1757 => to_unsigned(3368, 12), 1758 => to_unsigned(3404, 12), 1759 => to_unsigned(3301, 12), 1760 => to_unsigned(2291, 12), 1761 => to_unsigned(1696, 12), 1762 => to_unsigned(3082, 12), 1763 => to_unsigned(847, 12), 1764 => to_unsigned(3288, 12), 1765 => to_unsigned(3451, 12), 1766 => to_unsigned(2600, 12), 1767 => to_unsigned(2027, 12), 1768 => to_unsigned(23, 12), 1769 => to_unsigned(1787, 12), 1770 => to_unsigned(3737, 12), 1771 => to_unsigned(2878, 12), 1772 => to_unsigned(2822, 12), 1773 => to_unsigned(2335, 12), 1774 => to_unsigned(619, 12), 1775 => to_unsigned(2552, 12), 1776 => to_unsigned(1631, 12), 1777 => to_unsigned(840, 12), 1778 => to_unsigned(135, 12), 1779 => to_unsigned(936, 12), 1780 => to_unsigned(3748, 12), 1781 => to_unsigned(3763, 12), 1782 => to_unsigned(529, 12), 1783 => to_unsigned(3785, 12), 1784 => to_unsigned(1854, 12), 1785 => to_unsigned(2903, 12), 1786 => to_unsigned(3438, 12), 1787 => to_unsigned(1720, 12), 1788 => to_unsigned(3053, 12), 1789 => to_unsigned(2073, 12), 1790 => to_unsigned(3888, 12), 1791 => to_unsigned(3355, 12), 1792 => to_unsigned(923, 12), 1793 => to_unsigned(2061, 12), 1794 => to_unsigned(1833, 12), 1795 => to_unsigned(489, 12), 1796 => to_unsigned(1224, 12), 1797 => to_unsigned(3741, 12), 1798 => to_unsigned(3767, 12), 1799 => to_unsigned(1833, 12), 1800 => to_unsigned(3246, 12), 1801 => to_unsigned(1339, 12), 1802 => to_unsigned(3490, 12), 1803 => to_unsigned(1054, 12), 1804 => to_unsigned(2334, 12), 1805 => to_unsigned(788, 12), 1806 => to_unsigned(1818, 12), 1807 => to_unsigned(1259, 12), 1808 => to_unsigned(1449, 12), 1809 => to_unsigned(1292, 12), 1810 => to_unsigned(3471, 12), 1811 => to_unsigned(1143, 12), 1812 => to_unsigned(2592, 12), 1813 => to_unsigned(3416, 12), 1814 => to_unsigned(3939, 12), 1815 => to_unsigned(2883, 12), 1816 => to_unsigned(2090, 12), 1817 => to_unsigned(3844, 12), 1818 => to_unsigned(943, 12), 1819 => to_unsigned(1639, 12), 1820 => to_unsigned(2621, 12), 1821 => to_unsigned(149, 12), 1822 => to_unsigned(945, 12), 1823 => to_unsigned(1579, 12), 1824 => to_unsigned(3172, 12), 1825 => to_unsigned(2655, 12), 1826 => to_unsigned(2756, 12), 1827 => to_unsigned(3410, 12), 1828 => to_unsigned(1438, 12), 1829 => to_unsigned(664, 12), 1830 => to_unsigned(397, 12), 1831 => to_unsigned(1949, 12), 1832 => to_unsigned(2170, 12), 1833 => to_unsigned(798, 12), 1834 => to_unsigned(484, 12), 1835 => to_unsigned(1689, 12), 1836 => to_unsigned(3518, 12), 1837 => to_unsigned(1714, 12), 1838 => to_unsigned(3039, 12), 1839 => to_unsigned(2881, 12), 1840 => to_unsigned(3925, 12), 1841 => to_unsigned(2182, 12), 1842 => to_unsigned(1889, 12), 1843 => to_unsigned(1061, 12), 1844 => to_unsigned(3986, 12), 1845 => to_unsigned(281, 12), 1846 => to_unsigned(3466, 12), 1847 => to_unsigned(71, 12), 1848 => to_unsigned(205, 12), 1849 => to_unsigned(2277, 12), 1850 => to_unsigned(3710, 12), 1851 => to_unsigned(2769, 12), 1852 => to_unsigned(3328, 12), 1853 => to_unsigned(1425, 12), 1854 => to_unsigned(735, 12), 1855 => to_unsigned(3247, 12), 1856 => to_unsigned(3289, 12), 1857 => to_unsigned(1351, 12), 1858 => to_unsigned(3117, 12), 1859 => to_unsigned(51, 12), 1860 => to_unsigned(3755, 12), 1861 => to_unsigned(3984, 12), 1862 => to_unsigned(1623, 12), 1863 => to_unsigned(1895, 12), 1864 => to_unsigned(3556, 12), 1865 => to_unsigned(902, 12), 1866 => to_unsigned(4093, 12), 1867 => to_unsigned(3094, 12), 1868 => to_unsigned(2635, 12), 1869 => to_unsigned(1143, 12), 1870 => to_unsigned(3410, 12), 1871 => to_unsigned(1973, 12), 1872 => to_unsigned(2666, 12), 1873 => to_unsigned(2933, 12), 1874 => to_unsigned(1855, 12), 1875 => to_unsigned(1250, 12), 1876 => to_unsigned(1462, 12), 1877 => to_unsigned(1180, 12), 1878 => to_unsigned(3357, 12), 1879 => to_unsigned(2811, 12), 1880 => to_unsigned(3805, 12), 1881 => to_unsigned(2507, 12), 1882 => to_unsigned(44, 12), 1883 => to_unsigned(2513, 12), 1884 => to_unsigned(3509, 12), 1885 => to_unsigned(2966, 12), 1886 => to_unsigned(3234, 12), 1887 => to_unsigned(649, 12), 1888 => to_unsigned(513, 12), 1889 => to_unsigned(811, 12), 1890 => to_unsigned(3164, 12), 1891 => to_unsigned(645, 12), 1892 => to_unsigned(1288, 12), 1893 => to_unsigned(3098, 12), 1894 => to_unsigned(1030, 12), 1895 => to_unsigned(4020, 12), 1896 => to_unsigned(2121, 12), 1897 => to_unsigned(2111, 12), 1898 => to_unsigned(477, 12), 1899 => to_unsigned(1763, 12), 1900 => to_unsigned(1772, 12), 1901 => to_unsigned(1790, 12), 1902 => to_unsigned(285, 12), 1903 => to_unsigned(1178, 12), 1904 => to_unsigned(3521, 12), 1905 => to_unsigned(2039, 12), 1906 => to_unsigned(1125, 12), 1907 => to_unsigned(3474, 12), 1908 => to_unsigned(3994, 12), 1909 => to_unsigned(3555, 12), 1910 => to_unsigned(2275, 12), 1911 => to_unsigned(855, 12), 1912 => to_unsigned(3884, 12), 1913 => to_unsigned(3739, 12), 1914 => to_unsigned(575, 12), 1915 => to_unsigned(2731, 12), 1916 => to_unsigned(2756, 12), 1917 => to_unsigned(2114, 12), 1918 => to_unsigned(1823, 12), 1919 => to_unsigned(4025, 12), 1920 => to_unsigned(2888, 12), 1921 => to_unsigned(521, 12), 1922 => to_unsigned(2986, 12), 1923 => to_unsigned(916, 12), 1924 => to_unsigned(1335, 12), 1925 => to_unsigned(3232, 12), 1926 => to_unsigned(2120, 12), 1927 => to_unsigned(892, 12), 1928 => to_unsigned(2982, 12), 1929 => to_unsigned(2808, 12), 1930 => to_unsigned(492, 12), 1931 => to_unsigned(985, 12), 1932 => to_unsigned(404, 12), 1933 => to_unsigned(1426, 12), 1934 => to_unsigned(1492, 12), 1935 => to_unsigned(174, 12), 1936 => to_unsigned(1459, 12), 1937 => to_unsigned(1947, 12), 1938 => to_unsigned(1522, 12), 1939 => to_unsigned(2353, 12), 1940 => to_unsigned(3665, 12), 1941 => to_unsigned(153, 12), 1942 => to_unsigned(1585, 12), 1943 => to_unsigned(2950, 12), 1944 => to_unsigned(3161, 12), 1945 => to_unsigned(1573, 12), 1946 => to_unsigned(2473, 12), 1947 => to_unsigned(3654, 12), 1948 => to_unsigned(4075, 12), 1949 => to_unsigned(1305, 12), 1950 => to_unsigned(3068, 12), 1951 => to_unsigned(464, 12), 1952 => to_unsigned(1938, 12), 1953 => to_unsigned(314, 12), 1954 => to_unsigned(3183, 12), 1955 => to_unsigned(2666, 12), 1956 => to_unsigned(575, 12), 1957 => to_unsigned(1358, 12), 1958 => to_unsigned(3216, 12), 1959 => to_unsigned(3347, 12), 1960 => to_unsigned(932, 12), 1961 => to_unsigned(453, 12), 1962 => to_unsigned(531, 12), 1963 => to_unsigned(1706, 12), 1964 => to_unsigned(980, 12), 1965 => to_unsigned(3917, 12), 1966 => to_unsigned(2847, 12), 1967 => to_unsigned(525, 12), 1968 => to_unsigned(1038, 12), 1969 => to_unsigned(1932, 12), 1970 => to_unsigned(1973, 12), 1971 => to_unsigned(3126, 12), 1972 => to_unsigned(1710, 12), 1973 => to_unsigned(79, 12), 1974 => to_unsigned(3271, 12), 1975 => to_unsigned(1047, 12), 1976 => to_unsigned(1135, 12), 1977 => to_unsigned(2290, 12), 1978 => to_unsigned(2406, 12), 1979 => to_unsigned(2377, 12), 1980 => to_unsigned(1156, 12), 1981 => to_unsigned(1638, 12), 1982 => to_unsigned(1299, 12), 1983 => to_unsigned(231, 12), 1984 => to_unsigned(3225, 12), 1985 => to_unsigned(3600, 12), 1986 => to_unsigned(1960, 12), 1987 => to_unsigned(2732, 12), 1988 => to_unsigned(4089, 12), 1989 => to_unsigned(2534, 12), 1990 => to_unsigned(2504, 12), 1991 => to_unsigned(3093, 12), 1992 => to_unsigned(3951, 12), 1993 => to_unsigned(3269, 12), 1994 => to_unsigned(427, 12), 1995 => to_unsigned(1821, 12), 1996 => to_unsigned(2923, 12), 1997 => to_unsigned(1552, 12), 1998 => to_unsigned(1820, 12), 1999 => to_unsigned(1585, 12), 2000 => to_unsigned(1948, 12), 2001 => to_unsigned(1893, 12), 2002 => to_unsigned(263, 12), 2003 => to_unsigned(68, 12), 2004 => to_unsigned(1835, 12), 2005 => to_unsigned(461, 12), 2006 => to_unsigned(379, 12), 2007 => to_unsigned(3705, 12), 2008 => to_unsigned(1066, 12), 2009 => to_unsigned(1534, 12), 2010 => to_unsigned(1944, 12), 2011 => to_unsigned(3837, 12), 2012 => to_unsigned(1213, 12), 2013 => to_unsigned(955, 12), 2014 => to_unsigned(3201, 12), 2015 => to_unsigned(3704, 12), 2016 => to_unsigned(96, 12), 2017 => to_unsigned(3942, 12), 2018 => to_unsigned(1403, 12), 2019 => to_unsigned(1469, 12), 2020 => to_unsigned(1456, 12), 2021 => to_unsigned(2283, 12), 2022 => to_unsigned(3982, 12), 2023 => to_unsigned(482, 12), 2024 => to_unsigned(479, 12), 2025 => to_unsigned(3844, 12), 2026 => to_unsigned(473, 12), 2027 => to_unsigned(1945, 12), 2028 => to_unsigned(2215, 12), 2029 => to_unsigned(2940, 12), 2030 => to_unsigned(3078, 12), 2031 => to_unsigned(3963, 12), 2032 => to_unsigned(1081, 12), 2033 => to_unsigned(1782, 12), 2034 => to_unsigned(1258, 12), 2035 => to_unsigned(306, 12), 2036 => to_unsigned(735, 12), 2037 => to_unsigned(3265, 12), 2038 => to_unsigned(514, 12), 2039 => to_unsigned(856, 12), 2040 => to_unsigned(2999, 12), 2041 => to_unsigned(553, 12), 2042 => to_unsigned(2927, 12), 2043 => to_unsigned(518, 12), 2044 => to_unsigned(237, 12), 2045 => to_unsigned(2610, 12), 2046 => to_unsigned(2619, 12), 2047 => to_unsigned(2982, 12)),
            6 => (0 => to_unsigned(3656, 12), 1 => to_unsigned(3788, 12), 2 => to_unsigned(3139, 12), 3 => to_unsigned(2370, 12), 4 => to_unsigned(3484, 12), 5 => to_unsigned(1904, 12), 6 => to_unsigned(3531, 12), 7 => to_unsigned(1030, 12), 8 => to_unsigned(3754, 12), 9 => to_unsigned(3608, 12), 10 => to_unsigned(436, 12), 11 => to_unsigned(3600, 12), 12 => to_unsigned(1625, 12), 13 => to_unsigned(3269, 12), 14 => to_unsigned(3508, 12), 15 => to_unsigned(3854, 12), 16 => to_unsigned(379, 12), 17 => to_unsigned(1245, 12), 18 => to_unsigned(291, 12), 19 => to_unsigned(3115, 12), 20 => to_unsigned(1307, 12), 21 => to_unsigned(1021, 12), 22 => to_unsigned(620, 12), 23 => to_unsigned(311, 12), 24 => to_unsigned(3709, 12), 25 => to_unsigned(496, 12), 26 => to_unsigned(1350, 12), 27 => to_unsigned(1465, 12), 28 => to_unsigned(936, 12), 29 => to_unsigned(2749, 12), 30 => to_unsigned(1191, 12), 31 => to_unsigned(2864, 12), 32 => to_unsigned(3459, 12), 33 => to_unsigned(182, 12), 34 => to_unsigned(3979, 12), 35 => to_unsigned(1058, 12), 36 => to_unsigned(1734, 12), 37 => to_unsigned(1510, 12), 38 => to_unsigned(704, 12), 39 => to_unsigned(2530, 12), 40 => to_unsigned(1637, 12), 41 => to_unsigned(2846, 12), 42 => to_unsigned(17, 12), 43 => to_unsigned(75, 12), 44 => to_unsigned(1098, 12), 45 => to_unsigned(4076, 12), 46 => to_unsigned(3284, 12), 47 => to_unsigned(1342, 12), 48 => to_unsigned(2724, 12), 49 => to_unsigned(582, 12), 50 => to_unsigned(3837, 12), 51 => to_unsigned(3644, 12), 52 => to_unsigned(2439, 12), 53 => to_unsigned(1536, 12), 54 => to_unsigned(2881, 12), 55 => to_unsigned(1169, 12), 56 => to_unsigned(2092, 12), 57 => to_unsigned(3727, 12), 58 => to_unsigned(2491, 12), 59 => to_unsigned(302, 12), 60 => to_unsigned(1662, 12), 61 => to_unsigned(3692, 12), 62 => to_unsigned(3695, 12), 63 => to_unsigned(1640, 12), 64 => to_unsigned(2678, 12), 65 => to_unsigned(3541, 12), 66 => to_unsigned(184, 12), 67 => to_unsigned(1810, 12), 68 => to_unsigned(3062, 12), 69 => to_unsigned(166, 12), 70 => to_unsigned(2758, 12), 71 => to_unsigned(662, 12), 72 => to_unsigned(2070, 12), 73 => to_unsigned(3122, 12), 74 => to_unsigned(1220, 12), 75 => to_unsigned(3287, 12), 76 => to_unsigned(848, 12), 77 => to_unsigned(2132, 12), 78 => to_unsigned(1343, 12), 79 => to_unsigned(898, 12), 80 => to_unsigned(2374, 12), 81 => to_unsigned(1462, 12), 82 => to_unsigned(1057, 12), 83 => to_unsigned(1922, 12), 84 => to_unsigned(981, 12), 85 => to_unsigned(3455, 12), 86 => to_unsigned(3914, 12), 87 => to_unsigned(1387, 12), 88 => to_unsigned(3517, 12), 89 => to_unsigned(2601, 12), 90 => to_unsigned(1318, 12), 91 => to_unsigned(3316, 12), 92 => to_unsigned(3039, 12), 93 => to_unsigned(1765, 12), 94 => to_unsigned(2162, 12), 95 => to_unsigned(66, 12), 96 => to_unsigned(3179, 12), 97 => to_unsigned(1962, 12), 98 => to_unsigned(1977, 12), 99 => to_unsigned(3620, 12), 100 => to_unsigned(3013, 12), 101 => to_unsigned(3524, 12), 102 => to_unsigned(2237, 12), 103 => to_unsigned(2285, 12), 104 => to_unsigned(4025, 12), 105 => to_unsigned(3966, 12), 106 => to_unsigned(1025, 12), 107 => to_unsigned(1038, 12), 108 => to_unsigned(2079, 12), 109 => to_unsigned(2173, 12), 110 => to_unsigned(3897, 12), 111 => to_unsigned(1218, 12), 112 => to_unsigned(2609, 12), 113 => to_unsigned(952, 12), 114 => to_unsigned(2427, 12), 115 => to_unsigned(3893, 12), 116 => to_unsigned(2317, 12), 117 => to_unsigned(2841, 12), 118 => to_unsigned(3076, 12), 119 => to_unsigned(823, 12), 120 => to_unsigned(666, 12), 121 => to_unsigned(2088, 12), 122 => to_unsigned(782, 12), 123 => to_unsigned(3846, 12), 124 => to_unsigned(1838, 12), 125 => to_unsigned(3813, 12), 126 => to_unsigned(3683, 12), 127 => to_unsigned(1499, 12), 128 => to_unsigned(2300, 12), 129 => to_unsigned(1851, 12), 130 => to_unsigned(3959, 12), 131 => to_unsigned(374, 12), 132 => to_unsigned(2662, 12), 133 => to_unsigned(1921, 12), 134 => to_unsigned(91, 12), 135 => to_unsigned(809, 12), 136 => to_unsigned(507, 12), 137 => to_unsigned(3799, 12), 138 => to_unsigned(953, 12), 139 => to_unsigned(2275, 12), 140 => to_unsigned(2301, 12), 141 => to_unsigned(798, 12), 142 => to_unsigned(2612, 12), 143 => to_unsigned(2400, 12), 144 => to_unsigned(117, 12), 145 => to_unsigned(3745, 12), 146 => to_unsigned(2208, 12), 147 => to_unsigned(2638, 12), 148 => to_unsigned(1220, 12), 149 => to_unsigned(1822, 12), 150 => to_unsigned(53, 12), 151 => to_unsigned(1052, 12), 152 => to_unsigned(3890, 12), 153 => to_unsigned(885, 12), 154 => to_unsigned(2076, 12), 155 => to_unsigned(1550, 12), 156 => to_unsigned(1925, 12), 157 => to_unsigned(3361, 12), 158 => to_unsigned(332, 12), 159 => to_unsigned(2222, 12), 160 => to_unsigned(1886, 12), 161 => to_unsigned(245, 12), 162 => to_unsigned(1471, 12), 163 => to_unsigned(3985, 12), 164 => to_unsigned(3878, 12), 165 => to_unsigned(2125, 12), 166 => to_unsigned(3171, 12), 167 => to_unsigned(27, 12), 168 => to_unsigned(2979, 12), 169 => to_unsigned(3726, 12), 170 => to_unsigned(98, 12), 171 => to_unsigned(2333, 12), 172 => to_unsigned(2306, 12), 173 => to_unsigned(3350, 12), 174 => to_unsigned(1797, 12), 175 => to_unsigned(849, 12), 176 => to_unsigned(684, 12), 177 => to_unsigned(335, 12), 178 => to_unsigned(2233, 12), 179 => to_unsigned(3413, 12), 180 => to_unsigned(784, 12), 181 => to_unsigned(847, 12), 182 => to_unsigned(859, 12), 183 => to_unsigned(4045, 12), 184 => to_unsigned(3654, 12), 185 => to_unsigned(3139, 12), 186 => to_unsigned(1033, 12), 187 => to_unsigned(1843, 12), 188 => to_unsigned(571, 12), 189 => to_unsigned(2908, 12), 190 => to_unsigned(589, 12), 191 => to_unsigned(4068, 12), 192 => to_unsigned(1290, 12), 193 => to_unsigned(2911, 12), 194 => to_unsigned(2749, 12), 195 => to_unsigned(2932, 12), 196 => to_unsigned(3980, 12), 197 => to_unsigned(1447, 12), 198 => to_unsigned(116, 12), 199 => to_unsigned(1726, 12), 200 => to_unsigned(1666, 12), 201 => to_unsigned(28, 12), 202 => to_unsigned(2265, 12), 203 => to_unsigned(404, 12), 204 => to_unsigned(3248, 12), 205 => to_unsigned(1584, 12), 206 => to_unsigned(2607, 12), 207 => to_unsigned(1226, 12), 208 => to_unsigned(3852, 12), 209 => to_unsigned(3935, 12), 210 => to_unsigned(1095, 12), 211 => to_unsigned(2122, 12), 212 => to_unsigned(833, 12), 213 => to_unsigned(341, 12), 214 => to_unsigned(2012, 12), 215 => to_unsigned(2558, 12), 216 => to_unsigned(832, 12), 217 => to_unsigned(2507, 12), 218 => to_unsigned(1507, 12), 219 => to_unsigned(1078, 12), 220 => to_unsigned(3973, 12), 221 => to_unsigned(230, 12), 222 => to_unsigned(1794, 12), 223 => to_unsigned(1002, 12), 224 => to_unsigned(1088, 12), 225 => to_unsigned(570, 12), 226 => to_unsigned(3851, 12), 227 => to_unsigned(2878, 12), 228 => to_unsigned(2191, 12), 229 => to_unsigned(1185, 12), 230 => to_unsigned(3861, 12), 231 => to_unsigned(3939, 12), 232 => to_unsigned(1370, 12), 233 => to_unsigned(1387, 12), 234 => to_unsigned(1875, 12), 235 => to_unsigned(4095, 12), 236 => to_unsigned(574, 12), 237 => to_unsigned(3525, 12), 238 => to_unsigned(3954, 12), 239 => to_unsigned(1925, 12), 240 => to_unsigned(1685, 12), 241 => to_unsigned(2019, 12), 242 => to_unsigned(856, 12), 243 => to_unsigned(1619, 12), 244 => to_unsigned(1837, 12), 245 => to_unsigned(1564, 12), 246 => to_unsigned(1587, 12), 247 => to_unsigned(1983, 12), 248 => to_unsigned(2144, 12), 249 => to_unsigned(2776, 12), 250 => to_unsigned(3200, 12), 251 => to_unsigned(730, 12), 252 => to_unsigned(2813, 12), 253 => to_unsigned(108, 12), 254 => to_unsigned(1978, 12), 255 => to_unsigned(413, 12), 256 => to_unsigned(3594, 12), 257 => to_unsigned(2875, 12), 258 => to_unsigned(2702, 12), 259 => to_unsigned(1439, 12), 260 => to_unsigned(1662, 12), 261 => to_unsigned(2327, 12), 262 => to_unsigned(2759, 12), 263 => to_unsigned(3356, 12), 264 => to_unsigned(1662, 12), 265 => to_unsigned(2996, 12), 266 => to_unsigned(620, 12), 267 => to_unsigned(1733, 12), 268 => to_unsigned(3156, 12), 269 => to_unsigned(3927, 12), 270 => to_unsigned(758, 12), 271 => to_unsigned(2010, 12), 272 => to_unsigned(24, 12), 273 => to_unsigned(3488, 12), 274 => to_unsigned(522, 12), 275 => to_unsigned(1153, 12), 276 => to_unsigned(2373, 12), 277 => to_unsigned(3890, 12), 278 => to_unsigned(3197, 12), 279 => to_unsigned(471, 12), 280 => to_unsigned(1491, 12), 281 => to_unsigned(1489, 12), 282 => to_unsigned(1132, 12), 283 => to_unsigned(3493, 12), 284 => to_unsigned(2751, 12), 285 => to_unsigned(404, 12), 286 => to_unsigned(1056, 12), 287 => to_unsigned(1893, 12), 288 => to_unsigned(622, 12), 289 => to_unsigned(931, 12), 290 => to_unsigned(321, 12), 291 => to_unsigned(3713, 12), 292 => to_unsigned(1020, 12), 293 => to_unsigned(854, 12), 294 => to_unsigned(2065, 12), 295 => to_unsigned(1543, 12), 296 => to_unsigned(522, 12), 297 => to_unsigned(252, 12), 298 => to_unsigned(3971, 12), 299 => to_unsigned(3133, 12), 300 => to_unsigned(3815, 12), 301 => to_unsigned(32, 12), 302 => to_unsigned(2113, 12), 303 => to_unsigned(3851, 12), 304 => to_unsigned(1687, 12), 305 => to_unsigned(2680, 12), 306 => to_unsigned(1451, 12), 307 => to_unsigned(1453, 12), 308 => to_unsigned(2351, 12), 309 => to_unsigned(944, 12), 310 => to_unsigned(2119, 12), 311 => to_unsigned(3395, 12), 312 => to_unsigned(2764, 12), 313 => to_unsigned(82, 12), 314 => to_unsigned(3897, 12), 315 => to_unsigned(2962, 12), 316 => to_unsigned(2144, 12), 317 => to_unsigned(3584, 12), 318 => to_unsigned(964, 12), 319 => to_unsigned(1620, 12), 320 => to_unsigned(1900, 12), 321 => to_unsigned(1336, 12), 322 => to_unsigned(2678, 12), 323 => to_unsigned(3913, 12), 324 => to_unsigned(100, 12), 325 => to_unsigned(3351, 12), 326 => to_unsigned(3357, 12), 327 => to_unsigned(1453, 12), 328 => to_unsigned(1884, 12), 329 => to_unsigned(1256, 12), 330 => to_unsigned(2362, 12), 331 => to_unsigned(4012, 12), 332 => to_unsigned(3356, 12), 333 => to_unsigned(1537, 12), 334 => to_unsigned(1229, 12), 335 => to_unsigned(3173, 12), 336 => to_unsigned(2900, 12), 337 => to_unsigned(3974, 12), 338 => to_unsigned(4011, 12), 339 => to_unsigned(3627, 12), 340 => to_unsigned(1327, 12), 341 => to_unsigned(932, 12), 342 => to_unsigned(1259, 12), 343 => to_unsigned(3535, 12), 344 => to_unsigned(1688, 12), 345 => to_unsigned(2908, 12), 346 => to_unsigned(571, 12), 347 => to_unsigned(2780, 12), 348 => to_unsigned(695, 12), 349 => to_unsigned(3495, 12), 350 => to_unsigned(4038, 12), 351 => to_unsigned(2768, 12), 352 => to_unsigned(1337, 12), 353 => to_unsigned(87, 12), 354 => to_unsigned(1465, 12), 355 => to_unsigned(2270, 12), 356 => to_unsigned(1152, 12), 357 => to_unsigned(2282, 12), 358 => to_unsigned(816, 12), 359 => to_unsigned(1994, 12), 360 => to_unsigned(2209, 12), 361 => to_unsigned(85, 12), 362 => to_unsigned(3982, 12), 363 => to_unsigned(2487, 12), 364 => to_unsigned(1576, 12), 365 => to_unsigned(2869, 12), 366 => to_unsigned(3665, 12), 367 => to_unsigned(1004, 12), 368 => to_unsigned(1718, 12), 369 => to_unsigned(3058, 12), 370 => to_unsigned(2091, 12), 371 => to_unsigned(115, 12), 372 => to_unsigned(3732, 12), 373 => to_unsigned(3988, 12), 374 => to_unsigned(3929, 12), 375 => to_unsigned(1431, 12), 376 => to_unsigned(3987, 12), 377 => to_unsigned(3569, 12), 378 => to_unsigned(2376, 12), 379 => to_unsigned(3529, 12), 380 => to_unsigned(1626, 12), 381 => to_unsigned(345, 12), 382 => to_unsigned(904, 12), 383 => to_unsigned(1411, 12), 384 => to_unsigned(4061, 12), 385 => to_unsigned(2002, 12), 386 => to_unsigned(98, 12), 387 => to_unsigned(928, 12), 388 => to_unsigned(3218, 12), 389 => to_unsigned(3221, 12), 390 => to_unsigned(2705, 12), 391 => to_unsigned(2157, 12), 392 => to_unsigned(213, 12), 393 => to_unsigned(1739, 12), 394 => to_unsigned(4007, 12), 395 => to_unsigned(4074, 12), 396 => to_unsigned(3349, 12), 397 => to_unsigned(3142, 12), 398 => to_unsigned(4092, 12), 399 => to_unsigned(2463, 12), 400 => to_unsigned(755, 12), 401 => to_unsigned(3263, 12), 402 => to_unsigned(1700, 12), 403 => to_unsigned(998, 12), 404 => to_unsigned(3319, 12), 405 => to_unsigned(316, 12), 406 => to_unsigned(2410, 12), 407 => to_unsigned(684, 12), 408 => to_unsigned(3971, 12), 409 => to_unsigned(1185, 12), 410 => to_unsigned(1161, 12), 411 => to_unsigned(931, 12), 412 => to_unsigned(3861, 12), 413 => to_unsigned(2130, 12), 414 => to_unsigned(2297, 12), 415 => to_unsigned(2471, 12), 416 => to_unsigned(3361, 12), 417 => to_unsigned(651, 12), 418 => to_unsigned(148, 12), 419 => to_unsigned(653, 12), 420 => to_unsigned(3477, 12), 421 => to_unsigned(571, 12), 422 => to_unsigned(778, 12), 423 => to_unsigned(1971, 12), 424 => to_unsigned(3447, 12), 425 => to_unsigned(2241, 12), 426 => to_unsigned(1358, 12), 427 => to_unsigned(1303, 12), 428 => to_unsigned(2803, 12), 429 => to_unsigned(2781, 12), 430 => to_unsigned(2623, 12), 431 => to_unsigned(572, 12), 432 => to_unsigned(3408, 12), 433 => to_unsigned(3715, 12), 434 => to_unsigned(2224, 12), 435 => to_unsigned(3564, 12), 436 => to_unsigned(412, 12), 437 => to_unsigned(2233, 12), 438 => to_unsigned(2441, 12), 439 => to_unsigned(1296, 12), 440 => to_unsigned(2553, 12), 441 => to_unsigned(353, 12), 442 => to_unsigned(1938, 12), 443 => to_unsigned(926, 12), 444 => to_unsigned(1403, 12), 445 => to_unsigned(3738, 12), 446 => to_unsigned(1695, 12), 447 => to_unsigned(2617, 12), 448 => to_unsigned(910, 12), 449 => to_unsigned(2235, 12), 450 => to_unsigned(66, 12), 451 => to_unsigned(4059, 12), 452 => to_unsigned(2746, 12), 453 => to_unsigned(3876, 12), 454 => to_unsigned(3582, 12), 455 => to_unsigned(3390, 12), 456 => to_unsigned(550, 12), 457 => to_unsigned(3910, 12), 458 => to_unsigned(335, 12), 459 => to_unsigned(3779, 12), 460 => to_unsigned(2036, 12), 461 => to_unsigned(2529, 12), 462 => to_unsigned(673, 12), 463 => to_unsigned(3571, 12), 464 => to_unsigned(611, 12), 465 => to_unsigned(1243, 12), 466 => to_unsigned(3233, 12), 467 => to_unsigned(3247, 12), 468 => to_unsigned(2367, 12), 469 => to_unsigned(1251, 12), 470 => to_unsigned(3602, 12), 471 => to_unsigned(2833, 12), 472 => to_unsigned(1249, 12), 473 => to_unsigned(3313, 12), 474 => to_unsigned(1832, 12), 475 => to_unsigned(1169, 12), 476 => to_unsigned(3780, 12), 477 => to_unsigned(3945, 12), 478 => to_unsigned(1563, 12), 479 => to_unsigned(1236, 12), 480 => to_unsigned(2125, 12), 481 => to_unsigned(2190, 12), 482 => to_unsigned(415, 12), 483 => to_unsigned(3386, 12), 484 => to_unsigned(843, 12), 485 => to_unsigned(892, 12), 486 => to_unsigned(880, 12), 487 => to_unsigned(3538, 12), 488 => to_unsigned(405, 12), 489 => to_unsigned(3159, 12), 490 => to_unsigned(276, 12), 491 => to_unsigned(976, 12), 492 => to_unsigned(875, 12), 493 => to_unsigned(3379, 12), 494 => to_unsigned(452, 12), 495 => to_unsigned(1861, 12), 496 => to_unsigned(2819, 12), 497 => to_unsigned(3385, 12), 498 => to_unsigned(636, 12), 499 => to_unsigned(456, 12), 500 => to_unsigned(1309, 12), 501 => to_unsigned(1905, 12), 502 => to_unsigned(609, 12), 503 => to_unsigned(949, 12), 504 => to_unsigned(2878, 12), 505 => to_unsigned(3484, 12), 506 => to_unsigned(1683, 12), 507 => to_unsigned(3136, 12), 508 => to_unsigned(428, 12), 509 => to_unsigned(2898, 12), 510 => to_unsigned(3957, 12), 511 => to_unsigned(924, 12), 512 => to_unsigned(2146, 12), 513 => to_unsigned(807, 12), 514 => to_unsigned(1258, 12), 515 => to_unsigned(1113, 12), 516 => to_unsigned(3590, 12), 517 => to_unsigned(2685, 12), 518 => to_unsigned(3019, 12), 519 => to_unsigned(2820, 12), 520 => to_unsigned(500, 12), 521 => to_unsigned(711, 12), 522 => to_unsigned(1466, 12), 523 => to_unsigned(1120, 12), 524 => to_unsigned(3780, 12), 525 => to_unsigned(3181, 12), 526 => to_unsigned(1482, 12), 527 => to_unsigned(1484, 12), 528 => to_unsigned(1526, 12), 529 => to_unsigned(1180, 12), 530 => to_unsigned(273, 12), 531 => to_unsigned(3892, 12), 532 => to_unsigned(3181, 12), 533 => to_unsigned(2314, 12), 534 => to_unsigned(557, 12), 535 => to_unsigned(2541, 12), 536 => to_unsigned(4053, 12), 537 => to_unsigned(450, 12), 538 => to_unsigned(3327, 12), 539 => to_unsigned(355, 12), 540 => to_unsigned(1568, 12), 541 => to_unsigned(1263, 12), 542 => to_unsigned(1331, 12), 543 => to_unsigned(1473, 12), 544 => to_unsigned(245, 12), 545 => to_unsigned(1515, 12), 546 => to_unsigned(747, 12), 547 => to_unsigned(3334, 12), 548 => to_unsigned(4059, 12), 549 => to_unsigned(2519, 12), 550 => to_unsigned(2743, 12), 551 => to_unsigned(3035, 12), 552 => to_unsigned(3960, 12), 553 => to_unsigned(1296, 12), 554 => to_unsigned(1848, 12), 555 => to_unsigned(3709, 12), 556 => to_unsigned(2326, 12), 557 => to_unsigned(3610, 12), 558 => to_unsigned(1196, 12), 559 => to_unsigned(1783, 12), 560 => to_unsigned(1460, 12), 561 => to_unsigned(3662, 12), 562 => to_unsigned(1490, 12), 563 => to_unsigned(144, 12), 564 => to_unsigned(1736, 12), 565 => to_unsigned(1425, 12), 566 => to_unsigned(156, 12), 567 => to_unsigned(2595, 12), 568 => to_unsigned(2458, 12), 569 => to_unsigned(3884, 12), 570 => to_unsigned(3144, 12), 571 => to_unsigned(2018, 12), 572 => to_unsigned(1405, 12), 573 => to_unsigned(1838, 12), 574 => to_unsigned(1250, 12), 575 => to_unsigned(2146, 12), 576 => to_unsigned(3744, 12), 577 => to_unsigned(851, 12), 578 => to_unsigned(1727, 12), 579 => to_unsigned(2665, 12), 580 => to_unsigned(1132, 12), 581 => to_unsigned(2737, 12), 582 => to_unsigned(3116, 12), 583 => to_unsigned(1560, 12), 584 => to_unsigned(1601, 12), 585 => to_unsigned(3572, 12), 586 => to_unsigned(3042, 12), 587 => to_unsigned(3743, 12), 588 => to_unsigned(3491, 12), 589 => to_unsigned(1745, 12), 590 => to_unsigned(198, 12), 591 => to_unsigned(2238, 12), 592 => to_unsigned(2471, 12), 593 => to_unsigned(3329, 12), 594 => to_unsigned(3017, 12), 595 => to_unsigned(399, 12), 596 => to_unsigned(2018, 12), 597 => to_unsigned(431, 12), 598 => to_unsigned(3922, 12), 599 => to_unsigned(800, 12), 600 => to_unsigned(1654, 12), 601 => to_unsigned(98, 12), 602 => to_unsigned(2551, 12), 603 => to_unsigned(3705, 12), 604 => to_unsigned(2845, 12), 605 => to_unsigned(224, 12), 606 => to_unsigned(2332, 12), 607 => to_unsigned(2570, 12), 608 => to_unsigned(1239, 12), 609 => to_unsigned(3001, 12), 610 => to_unsigned(3199, 12), 611 => to_unsigned(3359, 12), 612 => to_unsigned(2759, 12), 613 => to_unsigned(3631, 12), 614 => to_unsigned(1879, 12), 615 => to_unsigned(1440, 12), 616 => to_unsigned(3352, 12), 617 => to_unsigned(1145, 12), 618 => to_unsigned(2468, 12), 619 => to_unsigned(297, 12), 620 => to_unsigned(1773, 12), 621 => to_unsigned(2871, 12), 622 => to_unsigned(3895, 12), 623 => to_unsigned(2501, 12), 624 => to_unsigned(733, 12), 625 => to_unsigned(4083, 12), 626 => to_unsigned(3434, 12), 627 => to_unsigned(2812, 12), 628 => to_unsigned(1363, 12), 629 => to_unsigned(1046, 12), 630 => to_unsigned(3097, 12), 631 => to_unsigned(894, 12), 632 => to_unsigned(1675, 12), 633 => to_unsigned(1850, 12), 634 => to_unsigned(4034, 12), 635 => to_unsigned(1743, 12), 636 => to_unsigned(416, 12), 637 => to_unsigned(3983, 12), 638 => to_unsigned(4020, 12), 639 => to_unsigned(2926, 12), 640 => to_unsigned(1023, 12), 641 => to_unsigned(3699, 12), 642 => to_unsigned(3040, 12), 643 => to_unsigned(2114, 12), 644 => to_unsigned(2959, 12), 645 => to_unsigned(2006, 12), 646 => to_unsigned(527, 12), 647 => to_unsigned(492, 12), 648 => to_unsigned(1766, 12), 649 => to_unsigned(3326, 12), 650 => to_unsigned(3046, 12), 651 => to_unsigned(3668, 12), 652 => to_unsigned(284, 12), 653 => to_unsigned(2412, 12), 654 => to_unsigned(3335, 12), 655 => to_unsigned(1602, 12), 656 => to_unsigned(3215, 12), 657 => to_unsigned(1574, 12), 658 => to_unsigned(69, 12), 659 => to_unsigned(1702, 12), 660 => to_unsigned(370, 12), 661 => to_unsigned(2903, 12), 662 => to_unsigned(1577, 12), 663 => to_unsigned(2453, 12), 664 => to_unsigned(3210, 12), 665 => to_unsigned(2418, 12), 666 => to_unsigned(2198, 12), 667 => to_unsigned(1351, 12), 668 => to_unsigned(3481, 12), 669 => to_unsigned(2810, 12), 670 => to_unsigned(103, 12), 671 => to_unsigned(1342, 12), 672 => to_unsigned(3576, 12), 673 => to_unsigned(649, 12), 674 => to_unsigned(3044, 12), 675 => to_unsigned(2481, 12), 676 => to_unsigned(744, 12), 677 => to_unsigned(2856, 12), 678 => to_unsigned(1577, 12), 679 => to_unsigned(917, 12), 680 => to_unsigned(3256, 12), 681 => to_unsigned(2745, 12), 682 => to_unsigned(821, 12), 683 => to_unsigned(3601, 12), 684 => to_unsigned(1785, 12), 685 => to_unsigned(651, 12), 686 => to_unsigned(3063, 12), 687 => to_unsigned(1245, 12), 688 => to_unsigned(506, 12), 689 => to_unsigned(2281, 12), 690 => to_unsigned(1786, 12), 691 => to_unsigned(289, 12), 692 => to_unsigned(1173, 12), 693 => to_unsigned(2463, 12), 694 => to_unsigned(909, 12), 695 => to_unsigned(1139, 12), 696 => to_unsigned(701, 12), 697 => to_unsigned(2499, 12), 698 => to_unsigned(2553, 12), 699 => to_unsigned(3438, 12), 700 => to_unsigned(1874, 12), 701 => to_unsigned(2749, 12), 702 => to_unsigned(674, 12), 703 => to_unsigned(189, 12), 704 => to_unsigned(1617, 12), 705 => to_unsigned(3167, 12), 706 => to_unsigned(2467, 12), 707 => to_unsigned(1038, 12), 708 => to_unsigned(3480, 12), 709 => to_unsigned(3426, 12), 710 => to_unsigned(2426, 12), 711 => to_unsigned(2220, 12), 712 => to_unsigned(2122, 12), 713 => to_unsigned(726, 12), 714 => to_unsigned(2257, 12), 715 => to_unsigned(1082, 12), 716 => to_unsigned(697, 12), 717 => to_unsigned(3319, 12), 718 => to_unsigned(2355, 12), 719 => to_unsigned(4086, 12), 720 => to_unsigned(1450, 12), 721 => to_unsigned(2157, 12), 722 => to_unsigned(1817, 12), 723 => to_unsigned(3596, 12), 724 => to_unsigned(1881, 12), 725 => to_unsigned(1433, 12), 726 => to_unsigned(1725, 12), 727 => to_unsigned(1504, 12), 728 => to_unsigned(1524, 12), 729 => to_unsigned(1654, 12), 730 => to_unsigned(3975, 12), 731 => to_unsigned(1308, 12), 732 => to_unsigned(1740, 12), 733 => to_unsigned(3392, 12), 734 => to_unsigned(2859, 12), 735 => to_unsigned(3034, 12), 736 => to_unsigned(243, 12), 737 => to_unsigned(1371, 12), 738 => to_unsigned(1142, 12), 739 => to_unsigned(2453, 12), 740 => to_unsigned(1203, 12), 741 => to_unsigned(2287, 12), 742 => to_unsigned(3816, 12), 743 => to_unsigned(3405, 12), 744 => to_unsigned(2889, 12), 745 => to_unsigned(3149, 12), 746 => to_unsigned(4095, 12), 747 => to_unsigned(2363, 12), 748 => to_unsigned(2739, 12), 749 => to_unsigned(976, 12), 750 => to_unsigned(2283, 12), 751 => to_unsigned(1145, 12), 752 => to_unsigned(3752, 12), 753 => to_unsigned(423, 12), 754 => to_unsigned(1396, 12), 755 => to_unsigned(2173, 12), 756 => to_unsigned(127, 12), 757 => to_unsigned(1301, 12), 758 => to_unsigned(1537, 12), 759 => to_unsigned(3154, 12), 760 => to_unsigned(1961, 12), 761 => to_unsigned(505, 12), 762 => to_unsigned(452, 12), 763 => to_unsigned(303, 12), 764 => to_unsigned(902, 12), 765 => to_unsigned(2609, 12), 766 => to_unsigned(2790, 12), 767 => to_unsigned(866, 12), 768 => to_unsigned(1253, 12), 769 => to_unsigned(229, 12), 770 => to_unsigned(435, 12), 771 => to_unsigned(65, 12), 772 => to_unsigned(2431, 12), 773 => to_unsigned(700, 12), 774 => to_unsigned(2020, 12), 775 => to_unsigned(61, 12), 776 => to_unsigned(3001, 12), 777 => to_unsigned(2268, 12), 778 => to_unsigned(2423, 12), 779 => to_unsigned(2754, 12), 780 => to_unsigned(3043, 12), 781 => to_unsigned(1354, 12), 782 => to_unsigned(317, 12), 783 => to_unsigned(2589, 12), 784 => to_unsigned(3119, 12), 785 => to_unsigned(1032, 12), 786 => to_unsigned(2685, 12), 787 => to_unsigned(3126, 12), 788 => to_unsigned(1507, 12), 789 => to_unsigned(190, 12), 790 => to_unsigned(3563, 12), 791 => to_unsigned(2367, 12), 792 => to_unsigned(824, 12), 793 => to_unsigned(990, 12), 794 => to_unsigned(1528, 12), 795 => to_unsigned(136, 12), 796 => to_unsigned(455, 12), 797 => to_unsigned(964, 12), 798 => to_unsigned(3636, 12), 799 => to_unsigned(783, 12), 800 => to_unsigned(3287, 12), 801 => to_unsigned(390, 12), 802 => to_unsigned(3850, 12), 803 => to_unsigned(1122, 12), 804 => to_unsigned(269, 12), 805 => to_unsigned(234, 12), 806 => to_unsigned(3762, 12), 807 => to_unsigned(846, 12), 808 => to_unsigned(3721, 12), 809 => to_unsigned(2015, 12), 810 => to_unsigned(200, 12), 811 => to_unsigned(62, 12), 812 => to_unsigned(3429, 12), 813 => to_unsigned(3087, 12), 814 => to_unsigned(3707, 12), 815 => to_unsigned(1399, 12), 816 => to_unsigned(696, 12), 817 => to_unsigned(3061, 12), 818 => to_unsigned(994, 12), 819 => to_unsigned(1532, 12), 820 => to_unsigned(3196, 12), 821 => to_unsigned(1304, 12), 822 => to_unsigned(3762, 12), 823 => to_unsigned(3885, 12), 824 => to_unsigned(1930, 12), 825 => to_unsigned(1682, 12), 826 => to_unsigned(989, 12), 827 => to_unsigned(255, 12), 828 => to_unsigned(3632, 12), 829 => to_unsigned(1003, 12), 830 => to_unsigned(3307, 12), 831 => to_unsigned(904, 12), 832 => to_unsigned(2806, 12), 833 => to_unsigned(2392, 12), 834 => to_unsigned(2412, 12), 835 => to_unsigned(1134, 12), 836 => to_unsigned(1242, 12), 837 => to_unsigned(3844, 12), 838 => to_unsigned(3970, 12), 839 => to_unsigned(223, 12), 840 => to_unsigned(3707, 12), 841 => to_unsigned(1781, 12), 842 => to_unsigned(3680, 12), 843 => to_unsigned(2477, 12), 844 => to_unsigned(2158, 12), 845 => to_unsigned(1286, 12), 846 => to_unsigned(1670, 12), 847 => to_unsigned(3471, 12), 848 => to_unsigned(1797, 12), 849 => to_unsigned(2887, 12), 850 => to_unsigned(2750, 12), 851 => to_unsigned(3572, 12), 852 => to_unsigned(1107, 12), 853 => to_unsigned(339, 12), 854 => to_unsigned(524, 12), 855 => to_unsigned(1329, 12), 856 => to_unsigned(3310, 12), 857 => to_unsigned(1502, 12), 858 => to_unsigned(3714, 12), 859 => to_unsigned(1396, 12), 860 => to_unsigned(2628, 12), 861 => to_unsigned(1800, 12), 862 => to_unsigned(211, 12), 863 => to_unsigned(1552, 12), 864 => to_unsigned(226, 12), 865 => to_unsigned(697, 12), 866 => to_unsigned(1369, 12), 867 => to_unsigned(492, 12), 868 => to_unsigned(2454, 12), 869 => to_unsigned(1103, 12), 870 => to_unsigned(1948, 12), 871 => to_unsigned(428, 12), 872 => to_unsigned(1073, 12), 873 => to_unsigned(2267, 12), 874 => to_unsigned(3848, 12), 875 => to_unsigned(3489, 12), 876 => to_unsigned(2945, 12), 877 => to_unsigned(3646, 12), 878 => to_unsigned(2430, 12), 879 => to_unsigned(1564, 12), 880 => to_unsigned(2454, 12), 881 => to_unsigned(3163, 12), 882 => to_unsigned(959, 12), 883 => to_unsigned(2138, 12), 884 => to_unsigned(959, 12), 885 => to_unsigned(2341, 12), 886 => to_unsigned(725, 12), 887 => to_unsigned(1785, 12), 888 => to_unsigned(3643, 12), 889 => to_unsigned(914, 12), 890 => to_unsigned(3652, 12), 891 => to_unsigned(2374, 12), 892 => to_unsigned(1424, 12), 893 => to_unsigned(2353, 12), 894 => to_unsigned(1475, 12), 895 => to_unsigned(394, 12), 896 => to_unsigned(3663, 12), 897 => to_unsigned(3833, 12), 898 => to_unsigned(3367, 12), 899 => to_unsigned(2358, 12), 900 => to_unsigned(542, 12), 901 => to_unsigned(3320, 12), 902 => to_unsigned(1228, 12), 903 => to_unsigned(1961, 12), 904 => to_unsigned(2237, 12), 905 => to_unsigned(3426, 12), 906 => to_unsigned(3492, 12), 907 => to_unsigned(1870, 12), 908 => to_unsigned(485, 12), 909 => to_unsigned(1909, 12), 910 => to_unsigned(3743, 12), 911 => to_unsigned(1736, 12), 912 => to_unsigned(112, 12), 913 => to_unsigned(3915, 12), 914 => to_unsigned(2211, 12), 915 => to_unsigned(3919, 12), 916 => to_unsigned(528, 12), 917 => to_unsigned(904, 12), 918 => to_unsigned(911, 12), 919 => to_unsigned(1623, 12), 920 => to_unsigned(2743, 12), 921 => to_unsigned(3124, 12), 922 => to_unsigned(315, 12), 923 => to_unsigned(1904, 12), 924 => to_unsigned(3481, 12), 925 => to_unsigned(684, 12), 926 => to_unsigned(595, 12), 927 => to_unsigned(3538, 12), 928 => to_unsigned(1687, 12), 929 => to_unsigned(541, 12), 930 => to_unsigned(1467, 12), 931 => to_unsigned(1784, 12), 932 => to_unsigned(3143, 12), 933 => to_unsigned(275, 12), 934 => to_unsigned(1093, 12), 935 => to_unsigned(2053, 12), 936 => to_unsigned(1834, 12), 937 => to_unsigned(1580, 12), 938 => to_unsigned(2, 12), 939 => to_unsigned(2731, 12), 940 => to_unsigned(1647, 12), 941 => to_unsigned(1423, 12), 942 => to_unsigned(101, 12), 943 => to_unsigned(2613, 12), 944 => to_unsigned(2685, 12), 945 => to_unsigned(1416, 12), 946 => to_unsigned(2744, 12), 947 => to_unsigned(1748, 12), 948 => to_unsigned(332, 12), 949 => to_unsigned(2752, 12), 950 => to_unsigned(3541, 12), 951 => to_unsigned(1395, 12), 952 => to_unsigned(2144, 12), 953 => to_unsigned(502, 12), 954 => to_unsigned(2178, 12), 955 => to_unsigned(2949, 12), 956 => to_unsigned(1653, 12), 957 => to_unsigned(159, 12), 958 => to_unsigned(1778, 12), 959 => to_unsigned(204, 12), 960 => to_unsigned(3671, 12), 961 => to_unsigned(1549, 12), 962 => to_unsigned(1496, 12), 963 => to_unsigned(1481, 12), 964 => to_unsigned(181, 12), 965 => to_unsigned(1711, 12), 966 => to_unsigned(395, 12), 967 => to_unsigned(3128, 12), 968 => to_unsigned(761, 12), 969 => to_unsigned(86, 12), 970 => to_unsigned(414, 12), 971 => to_unsigned(3658, 12), 972 => to_unsigned(547, 12), 973 => to_unsigned(342, 12), 974 => to_unsigned(2284, 12), 975 => to_unsigned(3434, 12), 976 => to_unsigned(788, 12), 977 => to_unsigned(1331, 12), 978 => to_unsigned(2239, 12), 979 => to_unsigned(2942, 12), 980 => to_unsigned(1440, 12), 981 => to_unsigned(3772, 12), 982 => to_unsigned(986, 12), 983 => to_unsigned(2458, 12), 984 => to_unsigned(173, 12), 985 => to_unsigned(3400, 12), 986 => to_unsigned(3708, 12), 987 => to_unsigned(1744, 12), 988 => to_unsigned(1166, 12), 989 => to_unsigned(3781, 12), 990 => to_unsigned(2989, 12), 991 => to_unsigned(841, 12), 992 => to_unsigned(1038, 12), 993 => to_unsigned(2523, 12), 994 => to_unsigned(4051, 12), 995 => to_unsigned(3886, 12), 996 => to_unsigned(1842, 12), 997 => to_unsigned(606, 12), 998 => to_unsigned(1097, 12), 999 => to_unsigned(3363, 12), 1000 => to_unsigned(2185, 12), 1001 => to_unsigned(2891, 12), 1002 => to_unsigned(1638, 12), 1003 => to_unsigned(4081, 12), 1004 => to_unsigned(4047, 12), 1005 => to_unsigned(2873, 12), 1006 => to_unsigned(1452, 12), 1007 => to_unsigned(1322, 12), 1008 => to_unsigned(3022, 12), 1009 => to_unsigned(2573, 12), 1010 => to_unsigned(3195, 12), 1011 => to_unsigned(3775, 12), 1012 => to_unsigned(2521, 12), 1013 => to_unsigned(2518, 12), 1014 => to_unsigned(596, 12), 1015 => to_unsigned(986, 12), 1016 => to_unsigned(734, 12), 1017 => to_unsigned(799, 12), 1018 => to_unsigned(4021, 12), 1019 => to_unsigned(815, 12), 1020 => to_unsigned(992, 12), 1021 => to_unsigned(882, 12), 1022 => to_unsigned(2055, 12), 1023 => to_unsigned(555, 12), 1024 => to_unsigned(1883, 12), 1025 => to_unsigned(418, 12), 1026 => to_unsigned(1609, 12), 1027 => to_unsigned(4061, 12), 1028 => to_unsigned(403, 12), 1029 => to_unsigned(830, 12), 1030 => to_unsigned(2329, 12), 1031 => to_unsigned(3357, 12), 1032 => to_unsigned(1972, 12), 1033 => to_unsigned(2476, 12), 1034 => to_unsigned(565, 12), 1035 => to_unsigned(811, 12), 1036 => to_unsigned(3090, 12), 1037 => to_unsigned(25, 12), 1038 => to_unsigned(3069, 12), 1039 => to_unsigned(2783, 12), 1040 => to_unsigned(359, 12), 1041 => to_unsigned(3733, 12), 1042 => to_unsigned(2754, 12), 1043 => to_unsigned(2713, 12), 1044 => to_unsigned(193, 12), 1045 => to_unsigned(3682, 12), 1046 => to_unsigned(1236, 12), 1047 => to_unsigned(1771, 12), 1048 => to_unsigned(3949, 12), 1049 => to_unsigned(1862, 12), 1050 => to_unsigned(3410, 12), 1051 => to_unsigned(2302, 12), 1052 => to_unsigned(1295, 12), 1053 => to_unsigned(88, 12), 1054 => to_unsigned(633, 12), 1055 => to_unsigned(3514, 12), 1056 => to_unsigned(2362, 12), 1057 => to_unsigned(1204, 12), 1058 => to_unsigned(2043, 12), 1059 => to_unsigned(478, 12), 1060 => to_unsigned(897, 12), 1061 => to_unsigned(1610, 12), 1062 => to_unsigned(3687, 12), 1063 => to_unsigned(2303, 12), 1064 => to_unsigned(1549, 12), 1065 => to_unsigned(2717, 12), 1066 => to_unsigned(1068, 12), 1067 => to_unsigned(3991, 12), 1068 => to_unsigned(2164, 12), 1069 => to_unsigned(1733, 12), 1070 => to_unsigned(2626, 12), 1071 => to_unsigned(2002, 12), 1072 => to_unsigned(608, 12), 1073 => to_unsigned(345, 12), 1074 => to_unsigned(581, 12), 1075 => to_unsigned(2703, 12), 1076 => to_unsigned(1126, 12), 1077 => to_unsigned(1830, 12), 1078 => to_unsigned(3891, 12), 1079 => to_unsigned(1168, 12), 1080 => to_unsigned(2505, 12), 1081 => to_unsigned(287, 12), 1082 => to_unsigned(2026, 12), 1083 => to_unsigned(1901, 12), 1084 => to_unsigned(2263, 12), 1085 => to_unsigned(3400, 12), 1086 => to_unsigned(3939, 12), 1087 => to_unsigned(920, 12), 1088 => to_unsigned(4031, 12), 1089 => to_unsigned(3933, 12), 1090 => to_unsigned(2313, 12), 1091 => to_unsigned(643, 12), 1092 => to_unsigned(1290, 12), 1093 => to_unsigned(2930, 12), 1094 => to_unsigned(2635, 12), 1095 => to_unsigned(330, 12), 1096 => to_unsigned(3237, 12), 1097 => to_unsigned(3185, 12), 1098 => to_unsigned(1425, 12), 1099 => to_unsigned(3806, 12), 1100 => to_unsigned(2015, 12), 1101 => to_unsigned(3809, 12), 1102 => to_unsigned(1382, 12), 1103 => to_unsigned(2270, 12), 1104 => to_unsigned(1514, 12), 1105 => to_unsigned(600, 12), 1106 => to_unsigned(2370, 12), 1107 => to_unsigned(708, 12), 1108 => to_unsigned(726, 12), 1109 => to_unsigned(2792, 12), 1110 => to_unsigned(1918, 12), 1111 => to_unsigned(3922, 12), 1112 => to_unsigned(547, 12), 1113 => to_unsigned(2205, 12), 1114 => to_unsigned(2617, 12), 1115 => to_unsigned(1698, 12), 1116 => to_unsigned(212, 12), 1117 => to_unsigned(4079, 12), 1118 => to_unsigned(2018, 12), 1119 => to_unsigned(893, 12), 1120 => to_unsigned(3030, 12), 1121 => to_unsigned(3984, 12), 1122 => to_unsigned(1767, 12), 1123 => to_unsigned(185, 12), 1124 => to_unsigned(3506, 12), 1125 => to_unsigned(294, 12), 1126 => to_unsigned(1762, 12), 1127 => to_unsigned(4023, 12), 1128 => to_unsigned(1434, 12), 1129 => to_unsigned(2274, 12), 1130 => to_unsigned(992, 12), 1131 => to_unsigned(119, 12), 1132 => to_unsigned(1689, 12), 1133 => to_unsigned(3360, 12), 1134 => to_unsigned(240, 12), 1135 => to_unsigned(2348, 12), 1136 => to_unsigned(4076, 12), 1137 => to_unsigned(1152, 12), 1138 => to_unsigned(3289, 12), 1139 => to_unsigned(1366, 12), 1140 => to_unsigned(3120, 12), 1141 => to_unsigned(1821, 12), 1142 => to_unsigned(3492, 12), 1143 => to_unsigned(1499, 12), 1144 => to_unsigned(2972, 12), 1145 => to_unsigned(2704, 12), 1146 => to_unsigned(2056, 12), 1147 => to_unsigned(1872, 12), 1148 => to_unsigned(3618, 12), 1149 => to_unsigned(996, 12), 1150 => to_unsigned(1710, 12), 1151 => to_unsigned(1184, 12), 1152 => to_unsigned(316, 12), 1153 => to_unsigned(2006, 12), 1154 => to_unsigned(1301, 12), 1155 => to_unsigned(3243, 12), 1156 => to_unsigned(224, 12), 1157 => to_unsigned(426, 12), 1158 => to_unsigned(2527, 12), 1159 => to_unsigned(119, 12), 1160 => to_unsigned(4070, 12), 1161 => to_unsigned(1389, 12), 1162 => to_unsigned(3265, 12), 1163 => to_unsigned(1070, 12), 1164 => to_unsigned(1986, 12), 1165 => to_unsigned(3867, 12), 1166 => to_unsigned(3401, 12), 1167 => to_unsigned(1457, 12), 1168 => to_unsigned(2780, 12), 1169 => to_unsigned(2069, 12), 1170 => to_unsigned(3707, 12), 1171 => to_unsigned(2404, 12), 1172 => to_unsigned(2834, 12), 1173 => to_unsigned(2918, 12), 1174 => to_unsigned(2918, 12), 1175 => to_unsigned(972, 12), 1176 => to_unsigned(209, 12), 1177 => to_unsigned(2594, 12), 1178 => to_unsigned(3556, 12), 1179 => to_unsigned(3171, 12), 1180 => to_unsigned(1202, 12), 1181 => to_unsigned(758, 12), 1182 => to_unsigned(1432, 12), 1183 => to_unsigned(2032, 12), 1184 => to_unsigned(2588, 12), 1185 => to_unsigned(1512, 12), 1186 => to_unsigned(1816, 12), 1187 => to_unsigned(1890, 12), 1188 => to_unsigned(871, 12), 1189 => to_unsigned(1564, 12), 1190 => to_unsigned(2526, 12), 1191 => to_unsigned(3223, 12), 1192 => to_unsigned(2672, 12), 1193 => to_unsigned(1477, 12), 1194 => to_unsigned(2373, 12), 1195 => to_unsigned(2721, 12), 1196 => to_unsigned(1698, 12), 1197 => to_unsigned(2787, 12), 1198 => to_unsigned(4017, 12), 1199 => to_unsigned(3190, 12), 1200 => to_unsigned(4020, 12), 1201 => to_unsigned(3892, 12), 1202 => to_unsigned(1087, 12), 1203 => to_unsigned(4051, 12), 1204 => to_unsigned(2036, 12), 1205 => to_unsigned(1453, 12), 1206 => to_unsigned(124, 12), 1207 => to_unsigned(3348, 12), 1208 => to_unsigned(1752, 12), 1209 => to_unsigned(2684, 12), 1210 => to_unsigned(2859, 12), 1211 => to_unsigned(1971, 12), 1212 => to_unsigned(2139, 12), 1213 => to_unsigned(1127, 12), 1214 => to_unsigned(3405, 12), 1215 => to_unsigned(404, 12), 1216 => to_unsigned(436, 12), 1217 => to_unsigned(2228, 12), 1218 => to_unsigned(2030, 12), 1219 => to_unsigned(3750, 12), 1220 => to_unsigned(1002, 12), 1221 => to_unsigned(1642, 12), 1222 => to_unsigned(134, 12), 1223 => to_unsigned(2490, 12), 1224 => to_unsigned(344, 12), 1225 => to_unsigned(1168, 12), 1226 => to_unsigned(1863, 12), 1227 => to_unsigned(1810, 12), 1228 => to_unsigned(1779, 12), 1229 => to_unsigned(3442, 12), 1230 => to_unsigned(1277, 12), 1231 => to_unsigned(1303, 12), 1232 => to_unsigned(2834, 12), 1233 => to_unsigned(2302, 12), 1234 => to_unsigned(1084, 12), 1235 => to_unsigned(1062, 12), 1236 => to_unsigned(3381, 12), 1237 => to_unsigned(3376, 12), 1238 => to_unsigned(3250, 12), 1239 => to_unsigned(2845, 12), 1240 => to_unsigned(1324, 12), 1241 => to_unsigned(2801, 12), 1242 => to_unsigned(604, 12), 1243 => to_unsigned(2838, 12), 1244 => to_unsigned(3713, 12), 1245 => to_unsigned(185, 12), 1246 => to_unsigned(2582, 12), 1247 => to_unsigned(2642, 12), 1248 => to_unsigned(205, 12), 1249 => to_unsigned(2174, 12), 1250 => to_unsigned(3902, 12), 1251 => to_unsigned(3069, 12), 1252 => to_unsigned(3375, 12), 1253 => to_unsigned(347, 12), 1254 => to_unsigned(1256, 12), 1255 => to_unsigned(496, 12), 1256 => to_unsigned(2133, 12), 1257 => to_unsigned(3906, 12), 1258 => to_unsigned(1619, 12), 1259 => to_unsigned(553, 12), 1260 => to_unsigned(435, 12), 1261 => to_unsigned(3316, 12), 1262 => to_unsigned(1577, 12), 1263 => to_unsigned(3847, 12), 1264 => to_unsigned(2628, 12), 1265 => to_unsigned(1090, 12), 1266 => to_unsigned(3043, 12), 1267 => to_unsigned(2367, 12), 1268 => to_unsigned(1421, 12), 1269 => to_unsigned(632, 12), 1270 => to_unsigned(2796, 12), 1271 => to_unsigned(113, 12), 1272 => to_unsigned(1436, 12), 1273 => to_unsigned(1062, 12), 1274 => to_unsigned(1284, 12), 1275 => to_unsigned(3494, 12), 1276 => to_unsigned(445, 12), 1277 => to_unsigned(1803, 12), 1278 => to_unsigned(2950, 12), 1279 => to_unsigned(2383, 12), 1280 => to_unsigned(2880, 12), 1281 => to_unsigned(2779, 12), 1282 => to_unsigned(1698, 12), 1283 => to_unsigned(111, 12), 1284 => to_unsigned(354, 12), 1285 => to_unsigned(1345, 12), 1286 => to_unsigned(2837, 12), 1287 => to_unsigned(2713, 12), 1288 => to_unsigned(2117, 12), 1289 => to_unsigned(3688, 12), 1290 => to_unsigned(791, 12), 1291 => to_unsigned(1618, 12), 1292 => to_unsigned(2203, 12), 1293 => to_unsigned(38, 12), 1294 => to_unsigned(307, 12), 1295 => to_unsigned(2572, 12), 1296 => to_unsigned(1941, 12), 1297 => to_unsigned(353, 12), 1298 => to_unsigned(1709, 12), 1299 => to_unsigned(3720, 12), 1300 => to_unsigned(641, 12), 1301 => to_unsigned(412, 12), 1302 => to_unsigned(1971, 12), 1303 => to_unsigned(2478, 12), 1304 => to_unsigned(2399, 12), 1305 => to_unsigned(1285, 12), 1306 => to_unsigned(3679, 12), 1307 => to_unsigned(358, 12), 1308 => to_unsigned(3857, 12), 1309 => to_unsigned(1655, 12), 1310 => to_unsigned(2989, 12), 1311 => to_unsigned(1314, 12), 1312 => to_unsigned(445, 12), 1313 => to_unsigned(1883, 12), 1314 => to_unsigned(2444, 12), 1315 => to_unsigned(2532, 12), 1316 => to_unsigned(1238, 12), 1317 => to_unsigned(2912, 12), 1318 => to_unsigned(2390, 12), 1319 => to_unsigned(3764, 12), 1320 => to_unsigned(3338, 12), 1321 => to_unsigned(556, 12), 1322 => to_unsigned(1904, 12), 1323 => to_unsigned(81, 12), 1324 => to_unsigned(3974, 12), 1325 => to_unsigned(2922, 12), 1326 => to_unsigned(231, 12), 1327 => to_unsigned(170, 12), 1328 => to_unsigned(601, 12), 1329 => to_unsigned(2596, 12), 1330 => to_unsigned(2657, 12), 1331 => to_unsigned(2864, 12), 1332 => to_unsigned(410, 12), 1333 => to_unsigned(1940, 12), 1334 => to_unsigned(3219, 12), 1335 => to_unsigned(1664, 12), 1336 => to_unsigned(3940, 12), 1337 => to_unsigned(3165, 12), 1338 => to_unsigned(1228, 12), 1339 => to_unsigned(1721, 12), 1340 => to_unsigned(2279, 12), 1341 => to_unsigned(1253, 12), 1342 => to_unsigned(3924, 12), 1343 => to_unsigned(3635, 12), 1344 => to_unsigned(1772, 12), 1345 => to_unsigned(2917, 12), 1346 => to_unsigned(2801, 12), 1347 => to_unsigned(2431, 12), 1348 => to_unsigned(292, 12), 1349 => to_unsigned(1271, 12), 1350 => to_unsigned(3818, 12), 1351 => to_unsigned(2121, 12), 1352 => to_unsigned(944, 12), 1353 => to_unsigned(530, 12), 1354 => to_unsigned(3527, 12), 1355 => to_unsigned(2891, 12), 1356 => to_unsigned(2725, 12), 1357 => to_unsigned(657, 12), 1358 => to_unsigned(845, 12), 1359 => to_unsigned(138, 12), 1360 => to_unsigned(2394, 12), 1361 => to_unsigned(3310, 12), 1362 => to_unsigned(2225, 12), 1363 => to_unsigned(3963, 12), 1364 => to_unsigned(3111, 12), 1365 => to_unsigned(109, 12), 1366 => to_unsigned(2072, 12), 1367 => to_unsigned(2496, 12), 1368 => to_unsigned(3257, 12), 1369 => to_unsigned(3436, 12), 1370 => to_unsigned(546, 12), 1371 => to_unsigned(4021, 12), 1372 => to_unsigned(4011, 12), 1373 => to_unsigned(3290, 12), 1374 => to_unsigned(117, 12), 1375 => to_unsigned(2300, 12), 1376 => to_unsigned(1731, 12), 1377 => to_unsigned(1351, 12), 1378 => to_unsigned(2334, 12), 1379 => to_unsigned(3234, 12), 1380 => to_unsigned(2577, 12), 1381 => to_unsigned(2828, 12), 1382 => to_unsigned(2894, 12), 1383 => to_unsigned(3634, 12), 1384 => to_unsigned(1210, 12), 1385 => to_unsigned(3337, 12), 1386 => to_unsigned(2628, 12), 1387 => to_unsigned(2425, 12), 1388 => to_unsigned(575, 12), 1389 => to_unsigned(3577, 12), 1390 => to_unsigned(3944, 12), 1391 => to_unsigned(3197, 12), 1392 => to_unsigned(1753, 12), 1393 => to_unsigned(790, 12), 1394 => to_unsigned(1051, 12), 1395 => to_unsigned(2593, 12), 1396 => to_unsigned(1047, 12), 1397 => to_unsigned(2743, 12), 1398 => to_unsigned(2166, 12), 1399 => to_unsigned(1700, 12), 1400 => to_unsigned(3570, 12), 1401 => to_unsigned(1307, 12), 1402 => to_unsigned(1968, 12), 1403 => to_unsigned(2202, 12), 1404 => to_unsigned(2921, 12), 1405 => to_unsigned(3042, 12), 1406 => to_unsigned(3903, 12), 1407 => to_unsigned(3116, 12), 1408 => to_unsigned(1513, 12), 1409 => to_unsigned(1858, 12), 1410 => to_unsigned(2453, 12), 1411 => to_unsigned(1281, 12), 1412 => to_unsigned(3588, 12), 1413 => to_unsigned(1509, 12), 1414 => to_unsigned(332, 12), 1415 => to_unsigned(3643, 12), 1416 => to_unsigned(409, 12), 1417 => to_unsigned(2874, 12), 1418 => to_unsigned(2756, 12), 1419 => to_unsigned(747, 12), 1420 => to_unsigned(927, 12), 1421 => to_unsigned(2048, 12), 1422 => to_unsigned(3141, 12), 1423 => to_unsigned(1594, 12), 1424 => to_unsigned(89, 12), 1425 => to_unsigned(1184, 12), 1426 => to_unsigned(396, 12), 1427 => to_unsigned(2035, 12), 1428 => to_unsigned(444, 12), 1429 => to_unsigned(3172, 12), 1430 => to_unsigned(3124, 12), 1431 => to_unsigned(3519, 12), 1432 => to_unsigned(539, 12), 1433 => to_unsigned(1757, 12), 1434 => to_unsigned(3630, 12), 1435 => to_unsigned(172, 12), 1436 => to_unsigned(2447, 12), 1437 => to_unsigned(843, 12), 1438 => to_unsigned(365, 12), 1439 => to_unsigned(2150, 12), 1440 => to_unsigned(487, 12), 1441 => to_unsigned(932, 12), 1442 => to_unsigned(2106, 12), 1443 => to_unsigned(3472, 12), 1444 => to_unsigned(2178, 12), 1445 => to_unsigned(2431, 12), 1446 => to_unsigned(3134, 12), 1447 => to_unsigned(328, 12), 1448 => to_unsigned(330, 12), 1449 => to_unsigned(591, 12), 1450 => to_unsigned(3884, 12), 1451 => to_unsigned(3679, 12), 1452 => to_unsigned(1460, 12), 1453 => to_unsigned(3061, 12), 1454 => to_unsigned(611, 12), 1455 => to_unsigned(3780, 12), 1456 => to_unsigned(1272, 12), 1457 => to_unsigned(534, 12), 1458 => to_unsigned(3186, 12), 1459 => to_unsigned(2744, 12), 1460 => to_unsigned(1640, 12), 1461 => to_unsigned(3318, 12), 1462 => to_unsigned(25, 12), 1463 => to_unsigned(592, 12), 1464 => to_unsigned(3523, 12), 1465 => to_unsigned(2780, 12), 1466 => to_unsigned(1947, 12), 1467 => to_unsigned(3487, 12), 1468 => to_unsigned(3217, 12), 1469 => to_unsigned(513, 12), 1470 => to_unsigned(726, 12), 1471 => to_unsigned(3807, 12), 1472 => to_unsigned(809, 12), 1473 => to_unsigned(173, 12), 1474 => to_unsigned(2028, 12), 1475 => to_unsigned(167, 12), 1476 => to_unsigned(2015, 12), 1477 => to_unsigned(4023, 12), 1478 => to_unsigned(4057, 12), 1479 => to_unsigned(344, 12), 1480 => to_unsigned(2461, 12), 1481 => to_unsigned(141, 12), 1482 => to_unsigned(1266, 12), 1483 => to_unsigned(2422, 12), 1484 => to_unsigned(2608, 12), 1485 => to_unsigned(3778, 12), 1486 => to_unsigned(3604, 12), 1487 => to_unsigned(929, 12), 1488 => to_unsigned(3248, 12), 1489 => to_unsigned(683, 12), 1490 => to_unsigned(2822, 12), 1491 => to_unsigned(2732, 12), 1492 => to_unsigned(3916, 12), 1493 => to_unsigned(3200, 12), 1494 => to_unsigned(410, 12), 1495 => to_unsigned(664, 12), 1496 => to_unsigned(3940, 12), 1497 => to_unsigned(3524, 12), 1498 => to_unsigned(181, 12), 1499 => to_unsigned(651, 12), 1500 => to_unsigned(2689, 12), 1501 => to_unsigned(642, 12), 1502 => to_unsigned(707, 12), 1503 => to_unsigned(1666, 12), 1504 => to_unsigned(1445, 12), 1505 => to_unsigned(3665, 12), 1506 => to_unsigned(3356, 12), 1507 => to_unsigned(2206, 12), 1508 => to_unsigned(1176, 12), 1509 => to_unsigned(3905, 12), 1510 => to_unsigned(195, 12), 1511 => to_unsigned(2662, 12), 1512 => to_unsigned(3026, 12), 1513 => to_unsigned(1254, 12), 1514 => to_unsigned(1313, 12), 1515 => to_unsigned(3791, 12), 1516 => to_unsigned(3162, 12), 1517 => to_unsigned(3976, 12), 1518 => to_unsigned(1089, 12), 1519 => to_unsigned(2840, 12), 1520 => to_unsigned(3271, 12), 1521 => to_unsigned(630, 12), 1522 => to_unsigned(3918, 12), 1523 => to_unsigned(3494, 12), 1524 => to_unsigned(2539, 12), 1525 => to_unsigned(938, 12), 1526 => to_unsigned(1279, 12), 1527 => to_unsigned(694, 12), 1528 => to_unsigned(3571, 12), 1529 => to_unsigned(135, 12), 1530 => to_unsigned(457, 12), 1531 => to_unsigned(2417, 12), 1532 => to_unsigned(2055, 12), 1533 => to_unsigned(2498, 12), 1534 => to_unsigned(3060, 12), 1535 => to_unsigned(2627, 12), 1536 => to_unsigned(133, 12), 1537 => to_unsigned(3079, 12), 1538 => to_unsigned(1094, 12), 1539 => to_unsigned(2959, 12), 1540 => to_unsigned(934, 12), 1541 => to_unsigned(3118, 12), 1542 => to_unsigned(192, 12), 1543 => to_unsigned(663, 12), 1544 => to_unsigned(3665, 12), 1545 => to_unsigned(363, 12), 1546 => to_unsigned(3984, 12), 1547 => to_unsigned(3303, 12), 1548 => to_unsigned(3063, 12), 1549 => to_unsigned(1914, 12), 1550 => to_unsigned(3065, 12), 1551 => to_unsigned(2556, 12), 1552 => to_unsigned(3304, 12), 1553 => to_unsigned(605, 12), 1554 => to_unsigned(3150, 12), 1555 => to_unsigned(1003, 12), 1556 => to_unsigned(2242, 12), 1557 => to_unsigned(831, 12), 1558 => to_unsigned(263, 12), 1559 => to_unsigned(503, 12), 1560 => to_unsigned(2576, 12), 1561 => to_unsigned(3056, 12), 1562 => to_unsigned(3204, 12), 1563 => to_unsigned(3597, 12), 1564 => to_unsigned(169, 12), 1565 => to_unsigned(502, 12), 1566 => to_unsigned(2649, 12), 1567 => to_unsigned(1800, 12), 1568 => to_unsigned(1498, 12), 1569 => to_unsigned(3663, 12), 1570 => to_unsigned(3245, 12), 1571 => to_unsigned(3119, 12), 1572 => to_unsigned(491, 12), 1573 => to_unsigned(2029, 12), 1574 => to_unsigned(4079, 12), 1575 => to_unsigned(1260, 12), 1576 => to_unsigned(713, 12), 1577 => to_unsigned(1396, 12), 1578 => to_unsigned(3581, 12), 1579 => to_unsigned(1212, 12), 1580 => to_unsigned(2001, 12), 1581 => to_unsigned(2543, 12), 1582 => to_unsigned(994, 12), 1583 => to_unsigned(188, 12), 1584 => to_unsigned(3249, 12), 1585 => to_unsigned(2021, 12), 1586 => to_unsigned(2383, 12), 1587 => to_unsigned(2306, 12), 1588 => to_unsigned(751, 12), 1589 => to_unsigned(1788, 12), 1590 => to_unsigned(3846, 12), 1591 => to_unsigned(3595, 12), 1592 => to_unsigned(2847, 12), 1593 => to_unsigned(2015, 12), 1594 => to_unsigned(3669, 12), 1595 => to_unsigned(3610, 12), 1596 => to_unsigned(4092, 12), 1597 => to_unsigned(2502, 12), 1598 => to_unsigned(2628, 12), 1599 => to_unsigned(3762, 12), 1600 => to_unsigned(1599, 12), 1601 => to_unsigned(3410, 12), 1602 => to_unsigned(3559, 12), 1603 => to_unsigned(4083, 12), 1604 => to_unsigned(724, 12), 1605 => to_unsigned(1847, 12), 1606 => to_unsigned(3039, 12), 1607 => to_unsigned(3282, 12), 1608 => to_unsigned(2474, 12), 1609 => to_unsigned(2920, 12), 1610 => to_unsigned(695, 12), 1611 => to_unsigned(3348, 12), 1612 => to_unsigned(724, 12), 1613 => to_unsigned(3976, 12), 1614 => to_unsigned(4006, 12), 1615 => to_unsigned(2507, 12), 1616 => to_unsigned(851, 12), 1617 => to_unsigned(1689, 12), 1618 => to_unsigned(2336, 12), 1619 => to_unsigned(1161, 12), 1620 => to_unsigned(3067, 12), 1621 => to_unsigned(168, 12), 1622 => to_unsigned(3356, 12), 1623 => to_unsigned(2443, 12), 1624 => to_unsigned(482, 12), 1625 => to_unsigned(2201, 12), 1626 => to_unsigned(2578, 12), 1627 => to_unsigned(2804, 12), 1628 => to_unsigned(1273, 12), 1629 => to_unsigned(1313, 12), 1630 => to_unsigned(753, 12), 1631 => to_unsigned(3867, 12), 1632 => to_unsigned(2736, 12), 1633 => to_unsigned(258, 12), 1634 => to_unsigned(1079, 12), 1635 => to_unsigned(2611, 12), 1636 => to_unsigned(1125, 12), 1637 => to_unsigned(90, 12), 1638 => to_unsigned(2719, 12), 1639 => to_unsigned(2767, 12), 1640 => to_unsigned(3926, 12), 1641 => to_unsigned(1224, 12), 1642 => to_unsigned(142, 12), 1643 => to_unsigned(487, 12), 1644 => to_unsigned(273, 12), 1645 => to_unsigned(306, 12), 1646 => to_unsigned(2586, 12), 1647 => to_unsigned(3355, 12), 1648 => to_unsigned(3009, 12), 1649 => to_unsigned(1063, 12), 1650 => to_unsigned(549, 12), 1651 => to_unsigned(4051, 12), 1652 => to_unsigned(3695, 12), 1653 => to_unsigned(3017, 12), 1654 => to_unsigned(3317, 12), 1655 => to_unsigned(2573, 12), 1656 => to_unsigned(1207, 12), 1657 => to_unsigned(1252, 12), 1658 => to_unsigned(1848, 12), 1659 => to_unsigned(3717, 12), 1660 => to_unsigned(459, 12), 1661 => to_unsigned(3655, 12), 1662 => to_unsigned(3885, 12), 1663 => to_unsigned(4029, 12), 1664 => to_unsigned(2372, 12), 1665 => to_unsigned(2199, 12), 1666 => to_unsigned(494, 12), 1667 => to_unsigned(2165, 12), 1668 => to_unsigned(2190, 12), 1669 => to_unsigned(3618, 12), 1670 => to_unsigned(716, 12), 1671 => to_unsigned(3669, 12), 1672 => to_unsigned(2005, 12), 1673 => to_unsigned(400, 12), 1674 => to_unsigned(871, 12), 1675 => to_unsigned(1249, 12), 1676 => to_unsigned(2669, 12), 1677 => to_unsigned(4044, 12), 1678 => to_unsigned(60, 12), 1679 => to_unsigned(1977, 12), 1680 => to_unsigned(1721, 12), 1681 => to_unsigned(1844, 12), 1682 => to_unsigned(4057, 12), 1683 => to_unsigned(1570, 12), 1684 => to_unsigned(248, 12), 1685 => to_unsigned(103, 12), 1686 => to_unsigned(9, 12), 1687 => to_unsigned(2778, 12), 1688 => to_unsigned(2009, 12), 1689 => to_unsigned(1452, 12), 1690 => to_unsigned(3429, 12), 1691 => to_unsigned(952, 12), 1692 => to_unsigned(1709, 12), 1693 => to_unsigned(2571, 12), 1694 => to_unsigned(303, 12), 1695 => to_unsigned(2376, 12), 1696 => to_unsigned(3216, 12), 1697 => to_unsigned(2493, 12), 1698 => to_unsigned(267, 12), 1699 => to_unsigned(2454, 12), 1700 => to_unsigned(866, 12), 1701 => to_unsigned(4038, 12), 1702 => to_unsigned(45, 12), 1703 => to_unsigned(1298, 12), 1704 => to_unsigned(2554, 12), 1705 => to_unsigned(3736, 12), 1706 => to_unsigned(554, 12), 1707 => to_unsigned(1587, 12), 1708 => to_unsigned(1178, 12), 1709 => to_unsigned(1882, 12), 1710 => to_unsigned(3261, 12), 1711 => to_unsigned(109, 12), 1712 => to_unsigned(1628, 12), 1713 => to_unsigned(178, 12), 1714 => to_unsigned(3691, 12), 1715 => to_unsigned(3084, 12), 1716 => to_unsigned(3748, 12), 1717 => to_unsigned(1444, 12), 1718 => to_unsigned(647, 12), 1719 => to_unsigned(439, 12), 1720 => to_unsigned(3229, 12), 1721 => to_unsigned(731, 12), 1722 => to_unsigned(1072, 12), 1723 => to_unsigned(638, 12), 1724 => to_unsigned(59, 12), 1725 => to_unsigned(3638, 12), 1726 => to_unsigned(1837, 12), 1727 => to_unsigned(4052, 12), 1728 => to_unsigned(624, 12), 1729 => to_unsigned(2257, 12), 1730 => to_unsigned(215, 12), 1731 => to_unsigned(553, 12), 1732 => to_unsigned(1491, 12), 1733 => to_unsigned(49, 12), 1734 => to_unsigned(1359, 12), 1735 => to_unsigned(2982, 12), 1736 => to_unsigned(2842, 12), 1737 => to_unsigned(1634, 12), 1738 => to_unsigned(473, 12), 1739 => to_unsigned(2445, 12), 1740 => to_unsigned(376, 12), 1741 => to_unsigned(1390, 12), 1742 => to_unsigned(710, 12), 1743 => to_unsigned(959, 12), 1744 => to_unsigned(1048, 12), 1745 => to_unsigned(2850, 12), 1746 => to_unsigned(1599, 12), 1747 => to_unsigned(398, 12), 1748 => to_unsigned(1194, 12), 1749 => to_unsigned(336, 12), 1750 => to_unsigned(985, 12), 1751 => to_unsigned(2269, 12), 1752 => to_unsigned(2211, 12), 1753 => to_unsigned(418, 12), 1754 => to_unsigned(3469, 12), 1755 => to_unsigned(233, 12), 1756 => to_unsigned(3297, 12), 1757 => to_unsigned(2995, 12), 1758 => to_unsigned(3080, 12), 1759 => to_unsigned(3164, 12), 1760 => to_unsigned(3347, 12), 1761 => to_unsigned(2078, 12), 1762 => to_unsigned(450, 12), 1763 => to_unsigned(3811, 12), 1764 => to_unsigned(1922, 12), 1765 => to_unsigned(938, 12), 1766 => to_unsigned(53, 12), 1767 => to_unsigned(882, 12), 1768 => to_unsigned(1485, 12), 1769 => to_unsigned(793, 12), 1770 => to_unsigned(2951, 12), 1771 => to_unsigned(742, 12), 1772 => to_unsigned(4024, 12), 1773 => to_unsigned(3828, 12), 1774 => to_unsigned(2909, 12), 1775 => to_unsigned(3344, 12), 1776 => to_unsigned(2881, 12), 1777 => to_unsigned(439, 12), 1778 => to_unsigned(2769, 12), 1779 => to_unsigned(3457, 12), 1780 => to_unsigned(2785, 12), 1781 => to_unsigned(1310, 12), 1782 => to_unsigned(773, 12), 1783 => to_unsigned(3637, 12), 1784 => to_unsigned(3344, 12), 1785 => to_unsigned(3971, 12), 1786 => to_unsigned(2515, 12), 1787 => to_unsigned(3951, 12), 1788 => to_unsigned(242, 12), 1789 => to_unsigned(500, 12), 1790 => to_unsigned(1916, 12), 1791 => to_unsigned(2035, 12), 1792 => to_unsigned(3659, 12), 1793 => to_unsigned(3821, 12), 1794 => to_unsigned(2122, 12), 1795 => to_unsigned(966, 12), 1796 => to_unsigned(2795, 12), 1797 => to_unsigned(3483, 12), 1798 => to_unsigned(1413, 12), 1799 => to_unsigned(3267, 12), 1800 => to_unsigned(2485, 12), 1801 => to_unsigned(1043, 12), 1802 => to_unsigned(1572, 12), 1803 => to_unsigned(516, 12), 1804 => to_unsigned(755, 12), 1805 => to_unsigned(3483, 12), 1806 => to_unsigned(2246, 12), 1807 => to_unsigned(3830, 12), 1808 => to_unsigned(2279, 12), 1809 => to_unsigned(2431, 12), 1810 => to_unsigned(2805, 12), 1811 => to_unsigned(3787, 12), 1812 => to_unsigned(1475, 12), 1813 => to_unsigned(978, 12), 1814 => to_unsigned(1690, 12), 1815 => to_unsigned(267, 12), 1816 => to_unsigned(1422, 12), 1817 => to_unsigned(85, 12), 1818 => to_unsigned(487, 12), 1819 => to_unsigned(1795, 12), 1820 => to_unsigned(3933, 12), 1821 => to_unsigned(133, 12), 1822 => to_unsigned(1173, 12), 1823 => to_unsigned(3936, 12), 1824 => to_unsigned(3864, 12), 1825 => to_unsigned(2699, 12), 1826 => to_unsigned(1055, 12), 1827 => to_unsigned(1423, 12), 1828 => to_unsigned(2170, 12), 1829 => to_unsigned(712, 12), 1830 => to_unsigned(1714, 12), 1831 => to_unsigned(363, 12), 1832 => to_unsigned(3845, 12), 1833 => to_unsigned(1422, 12), 1834 => to_unsigned(26, 12), 1835 => to_unsigned(472, 12), 1836 => to_unsigned(2725, 12), 1837 => to_unsigned(1394, 12), 1838 => to_unsigned(2810, 12), 1839 => to_unsigned(3992, 12), 1840 => to_unsigned(413, 12), 1841 => to_unsigned(3895, 12), 1842 => to_unsigned(1171, 12), 1843 => to_unsigned(2209, 12), 1844 => to_unsigned(1734, 12), 1845 => to_unsigned(2889, 12), 1846 => to_unsigned(2141, 12), 1847 => to_unsigned(3178, 12), 1848 => to_unsigned(3237, 12), 1849 => to_unsigned(2235, 12), 1850 => to_unsigned(3861, 12), 1851 => to_unsigned(4015, 12), 1852 => to_unsigned(2956, 12), 1853 => to_unsigned(3516, 12), 1854 => to_unsigned(1781, 12), 1855 => to_unsigned(349, 12), 1856 => to_unsigned(532, 12), 1857 => to_unsigned(1610, 12), 1858 => to_unsigned(1012, 12), 1859 => to_unsigned(717, 12), 1860 => to_unsigned(2687, 12), 1861 => to_unsigned(452, 12), 1862 => to_unsigned(3819, 12), 1863 => to_unsigned(2722, 12), 1864 => to_unsigned(4078, 12), 1865 => to_unsigned(3122, 12), 1866 => to_unsigned(783, 12), 1867 => to_unsigned(4028, 12), 1868 => to_unsigned(1829, 12), 1869 => to_unsigned(1716, 12), 1870 => to_unsigned(892, 12), 1871 => to_unsigned(1925, 12), 1872 => to_unsigned(1413, 12), 1873 => to_unsigned(1999, 12), 1874 => to_unsigned(345, 12), 1875 => to_unsigned(3506, 12), 1876 => to_unsigned(2621, 12), 1877 => to_unsigned(856, 12), 1878 => to_unsigned(449, 12), 1879 => to_unsigned(2243, 12), 1880 => to_unsigned(209, 12), 1881 => to_unsigned(3680, 12), 1882 => to_unsigned(1334, 12), 1883 => to_unsigned(3997, 12), 1884 => to_unsigned(781, 12), 1885 => to_unsigned(3751, 12), 1886 => to_unsigned(1431, 12), 1887 => to_unsigned(3428, 12), 1888 => to_unsigned(2840, 12), 1889 => to_unsigned(1194, 12), 1890 => to_unsigned(820, 12), 1891 => to_unsigned(2183, 12), 1892 => to_unsigned(3723, 12), 1893 => to_unsigned(3324, 12), 1894 => to_unsigned(1770, 12), 1895 => to_unsigned(1938, 12), 1896 => to_unsigned(3794, 12), 1897 => to_unsigned(3359, 12), 1898 => to_unsigned(51, 12), 1899 => to_unsigned(1574, 12), 1900 => to_unsigned(1146, 12), 1901 => to_unsigned(419, 12), 1902 => to_unsigned(2666, 12), 1903 => to_unsigned(3806, 12), 1904 => to_unsigned(1734, 12), 1905 => to_unsigned(3563, 12), 1906 => to_unsigned(2666, 12), 1907 => to_unsigned(436, 12), 1908 => to_unsigned(167, 12), 1909 => to_unsigned(2140, 12), 1910 => to_unsigned(3460, 12), 1911 => to_unsigned(2009, 12), 1912 => to_unsigned(2173, 12), 1913 => to_unsigned(666, 12), 1914 => to_unsigned(1638, 12), 1915 => to_unsigned(2700, 12), 1916 => to_unsigned(2652, 12), 1917 => to_unsigned(528, 12), 1918 => to_unsigned(1715, 12), 1919 => to_unsigned(2983, 12), 1920 => to_unsigned(1748, 12), 1921 => to_unsigned(1210, 12), 1922 => to_unsigned(3209, 12), 1923 => to_unsigned(1012, 12), 1924 => to_unsigned(2879, 12), 1925 => to_unsigned(1711, 12), 1926 => to_unsigned(2775, 12), 1927 => to_unsigned(1701, 12), 1928 => to_unsigned(711, 12), 1929 => to_unsigned(3870, 12), 1930 => to_unsigned(781, 12), 1931 => to_unsigned(2360, 12), 1932 => to_unsigned(2178, 12), 1933 => to_unsigned(480, 12), 1934 => to_unsigned(3252, 12), 1935 => to_unsigned(2710, 12), 1936 => to_unsigned(1758, 12), 1937 => to_unsigned(2968, 12), 1938 => to_unsigned(1118, 12), 1939 => to_unsigned(282, 12), 1940 => to_unsigned(2361, 12), 1941 => to_unsigned(1518, 12), 1942 => to_unsigned(2280, 12), 1943 => to_unsigned(1933, 12), 1944 => to_unsigned(2246, 12), 1945 => to_unsigned(229, 12), 1946 => to_unsigned(2243, 12), 1947 => to_unsigned(912, 12), 1948 => to_unsigned(2573, 12), 1949 => to_unsigned(650, 12), 1950 => to_unsigned(208, 12), 1951 => to_unsigned(3569, 12), 1952 => to_unsigned(2965, 12), 1953 => to_unsigned(340, 12), 1954 => to_unsigned(1232, 12), 1955 => to_unsigned(1644, 12), 1956 => to_unsigned(2596, 12), 1957 => to_unsigned(2804, 12), 1958 => to_unsigned(2099, 12), 1959 => to_unsigned(2034, 12), 1960 => to_unsigned(305, 12), 1961 => to_unsigned(1552, 12), 1962 => to_unsigned(3490, 12), 1963 => to_unsigned(489, 12), 1964 => to_unsigned(199, 12), 1965 => to_unsigned(3551, 12), 1966 => to_unsigned(1398, 12), 1967 => to_unsigned(362, 12), 1968 => to_unsigned(1917, 12), 1969 => to_unsigned(3495, 12), 1970 => to_unsigned(1034, 12), 1971 => to_unsigned(3666, 12), 1972 => to_unsigned(892, 12), 1973 => to_unsigned(2587, 12), 1974 => to_unsigned(2407, 12), 1975 => to_unsigned(1280, 12), 1976 => to_unsigned(2228, 12), 1977 => to_unsigned(3913, 12), 1978 => to_unsigned(3410, 12), 1979 => to_unsigned(1925, 12), 1980 => to_unsigned(980, 12), 1981 => to_unsigned(1675, 12), 1982 => to_unsigned(3456, 12), 1983 => to_unsigned(2825, 12), 1984 => to_unsigned(3369, 12), 1985 => to_unsigned(1544, 12), 1986 => to_unsigned(372, 12), 1987 => to_unsigned(1221, 12), 1988 => to_unsigned(2558, 12), 1989 => to_unsigned(25, 12), 1990 => to_unsigned(1515, 12), 1991 => to_unsigned(2597, 12), 1992 => to_unsigned(860, 12), 1993 => to_unsigned(2494, 12), 1994 => to_unsigned(3921, 12), 1995 => to_unsigned(1196, 12), 1996 => to_unsigned(2825, 12), 1997 => to_unsigned(1999, 12), 1998 => to_unsigned(838, 12), 1999 => to_unsigned(315, 12), 2000 => to_unsigned(3826, 12), 2001 => to_unsigned(3466, 12), 2002 => to_unsigned(139, 12), 2003 => to_unsigned(1286, 12), 2004 => to_unsigned(1939, 12), 2005 => to_unsigned(863, 12), 2006 => to_unsigned(3927, 12), 2007 => to_unsigned(2179, 12), 2008 => to_unsigned(747, 12), 2009 => to_unsigned(2414, 12), 2010 => to_unsigned(3950, 12), 2011 => to_unsigned(375, 12), 2012 => to_unsigned(3122, 12), 2013 => to_unsigned(389, 12), 2014 => to_unsigned(4002, 12), 2015 => to_unsigned(246, 12), 2016 => to_unsigned(3575, 12), 2017 => to_unsigned(1259, 12), 2018 => to_unsigned(1116, 12), 2019 => to_unsigned(784, 12), 2020 => to_unsigned(3445, 12), 2021 => to_unsigned(44, 12), 2022 => to_unsigned(263, 12), 2023 => to_unsigned(100, 12), 2024 => to_unsigned(3662, 12), 2025 => to_unsigned(1201, 12), 2026 => to_unsigned(2053, 12), 2027 => to_unsigned(1750, 12), 2028 => to_unsigned(2072, 12), 2029 => to_unsigned(4021, 12), 2030 => to_unsigned(3171, 12), 2031 => to_unsigned(141, 12), 2032 => to_unsigned(3299, 12), 2033 => to_unsigned(1542, 12), 2034 => to_unsigned(1928, 12), 2035 => to_unsigned(2691, 12), 2036 => to_unsigned(828, 12), 2037 => to_unsigned(3709, 12), 2038 => to_unsigned(806, 12), 2039 => to_unsigned(1710, 12), 2040 => to_unsigned(2413, 12), 2041 => to_unsigned(3201, 12), 2042 => to_unsigned(918, 12), 2043 => to_unsigned(3505, 12), 2044 => to_unsigned(674, 12), 2045 => to_unsigned(2189, 12), 2046 => to_unsigned(1359, 12), 2047 => to_unsigned(2483, 12)),
            7 => (0 => to_unsigned(3413, 12), 1 => to_unsigned(1039, 12), 2 => to_unsigned(3845, 12), 3 => to_unsigned(3389, 12), 4 => to_unsigned(3100, 12), 5 => to_unsigned(1494, 12), 6 => to_unsigned(2563, 12), 7 => to_unsigned(2662, 12), 8 => to_unsigned(3696, 12), 9 => to_unsigned(181, 12), 10 => to_unsigned(2768, 12), 11 => to_unsigned(4019, 12), 12 => to_unsigned(2874, 12), 13 => to_unsigned(3456, 12), 14 => to_unsigned(3082, 12), 15 => to_unsigned(1909, 12), 16 => to_unsigned(2007, 12), 17 => to_unsigned(1182, 12), 18 => to_unsigned(850, 12), 19 => to_unsigned(2053, 12), 20 => to_unsigned(1460, 12), 21 => to_unsigned(1544, 12), 22 => to_unsigned(2062, 12), 23 => to_unsigned(3356, 12), 24 => to_unsigned(1678, 12), 25 => to_unsigned(441, 12), 26 => to_unsigned(2708, 12), 27 => to_unsigned(909, 12), 28 => to_unsigned(2958, 12), 29 => to_unsigned(1989, 12), 30 => to_unsigned(609, 12), 31 => to_unsigned(423, 12), 32 => to_unsigned(369, 12), 33 => to_unsigned(1557, 12), 34 => to_unsigned(1059, 12), 35 => to_unsigned(22, 12), 36 => to_unsigned(2529, 12), 37 => to_unsigned(2032, 12), 38 => to_unsigned(679, 12), 39 => to_unsigned(3305, 12), 40 => to_unsigned(1274, 12), 41 => to_unsigned(1152, 12), 42 => to_unsigned(3695, 12), 43 => to_unsigned(419, 12), 44 => to_unsigned(2305, 12), 45 => to_unsigned(3025, 12), 46 => to_unsigned(2694, 12), 47 => to_unsigned(3889, 12), 48 => to_unsigned(3442, 12), 49 => to_unsigned(3782, 12), 50 => to_unsigned(2466, 12), 51 => to_unsigned(2322, 12), 52 => to_unsigned(2468, 12), 53 => to_unsigned(1360, 12), 54 => to_unsigned(669, 12), 55 => to_unsigned(3720, 12), 56 => to_unsigned(3048, 12), 57 => to_unsigned(3883, 12), 58 => to_unsigned(2976, 12), 59 => to_unsigned(2978, 12), 60 => to_unsigned(3985, 12), 61 => to_unsigned(3515, 12), 62 => to_unsigned(1405, 12), 63 => to_unsigned(2672, 12), 64 => to_unsigned(3141, 12), 65 => to_unsigned(1289, 12), 66 => to_unsigned(522, 12), 67 => to_unsigned(2604, 12), 68 => to_unsigned(2537, 12), 69 => to_unsigned(3561, 12), 70 => to_unsigned(976, 12), 71 => to_unsigned(1523, 12), 72 => to_unsigned(3544, 12), 73 => to_unsigned(2072, 12), 74 => to_unsigned(3670, 12), 75 => to_unsigned(1860, 12), 76 => to_unsigned(1286, 12), 77 => to_unsigned(916, 12), 78 => to_unsigned(1856, 12), 79 => to_unsigned(3888, 12), 80 => to_unsigned(2798, 12), 81 => to_unsigned(1462, 12), 82 => to_unsigned(2507, 12), 83 => to_unsigned(3431, 12), 84 => to_unsigned(2189, 12), 85 => to_unsigned(2527, 12), 86 => to_unsigned(3345, 12), 87 => to_unsigned(1735, 12), 88 => to_unsigned(3647, 12), 89 => to_unsigned(2107, 12), 90 => to_unsigned(1354, 12), 91 => to_unsigned(3004, 12), 92 => to_unsigned(3055, 12), 93 => to_unsigned(2562, 12), 94 => to_unsigned(3170, 12), 95 => to_unsigned(1491, 12), 96 => to_unsigned(1550, 12), 97 => to_unsigned(3154, 12), 98 => to_unsigned(3869, 12), 99 => to_unsigned(2751, 12), 100 => to_unsigned(1277, 12), 101 => to_unsigned(3232, 12), 102 => to_unsigned(586, 12), 103 => to_unsigned(3544, 12), 104 => to_unsigned(3237, 12), 105 => to_unsigned(2904, 12), 106 => to_unsigned(1842, 12), 107 => to_unsigned(4004, 12), 108 => to_unsigned(598, 12), 109 => to_unsigned(629, 12), 110 => to_unsigned(2966, 12), 111 => to_unsigned(273, 12), 112 => to_unsigned(2161, 12), 113 => to_unsigned(81, 12), 114 => to_unsigned(1083, 12), 115 => to_unsigned(1546, 12), 116 => to_unsigned(2842, 12), 117 => to_unsigned(2460, 12), 118 => to_unsigned(1039, 12), 119 => to_unsigned(1970, 12), 120 => to_unsigned(3658, 12), 121 => to_unsigned(1936, 12), 122 => to_unsigned(244, 12), 123 => to_unsigned(1728, 12), 124 => to_unsigned(1750, 12), 125 => to_unsigned(3630, 12), 126 => to_unsigned(1503, 12), 127 => to_unsigned(2334, 12), 128 => to_unsigned(4014, 12), 129 => to_unsigned(3847, 12), 130 => to_unsigned(510, 12), 131 => to_unsigned(464, 12), 132 => to_unsigned(2967, 12), 133 => to_unsigned(1866, 12), 134 => to_unsigned(889, 12), 135 => to_unsigned(64, 12), 136 => to_unsigned(2175, 12), 137 => to_unsigned(615, 12), 138 => to_unsigned(2051, 12), 139 => to_unsigned(1638, 12), 140 => to_unsigned(3078, 12), 141 => to_unsigned(1800, 12), 142 => to_unsigned(2497, 12), 143 => to_unsigned(2262, 12), 144 => to_unsigned(704, 12), 145 => to_unsigned(1159, 12), 146 => to_unsigned(807, 12), 147 => to_unsigned(3725, 12), 148 => to_unsigned(1308, 12), 149 => to_unsigned(2153, 12), 150 => to_unsigned(2430, 12), 151 => to_unsigned(3665, 12), 152 => to_unsigned(3166, 12), 153 => to_unsigned(2435, 12), 154 => to_unsigned(2370, 12), 155 => to_unsigned(1299, 12), 156 => to_unsigned(2244, 12), 157 => to_unsigned(3683, 12), 158 => to_unsigned(1452, 12), 159 => to_unsigned(2249, 12), 160 => to_unsigned(3351, 12), 161 => to_unsigned(1759, 12), 162 => to_unsigned(3074, 12), 163 => to_unsigned(1995, 12), 164 => to_unsigned(1090, 12), 165 => to_unsigned(1686, 12), 166 => to_unsigned(1217, 12), 167 => to_unsigned(3525, 12), 168 => to_unsigned(3637, 12), 169 => to_unsigned(3482, 12), 170 => to_unsigned(936, 12), 171 => to_unsigned(390, 12), 172 => to_unsigned(653, 12), 173 => to_unsigned(948, 12), 174 => to_unsigned(1205, 12), 175 => to_unsigned(1389, 12), 176 => to_unsigned(3333, 12), 177 => to_unsigned(2746, 12), 178 => to_unsigned(422, 12), 179 => to_unsigned(3913, 12), 180 => to_unsigned(1605, 12), 181 => to_unsigned(3542, 12), 182 => to_unsigned(666, 12), 183 => to_unsigned(1582, 12), 184 => to_unsigned(903, 12), 185 => to_unsigned(798, 12), 186 => to_unsigned(2406, 12), 187 => to_unsigned(1911, 12), 188 => to_unsigned(1414, 12), 189 => to_unsigned(3751, 12), 190 => to_unsigned(3604, 12), 191 => to_unsigned(3570, 12), 192 => to_unsigned(560, 12), 193 => to_unsigned(3034, 12), 194 => to_unsigned(2113, 12), 195 => to_unsigned(420, 12), 196 => to_unsigned(900, 12), 197 => to_unsigned(1693, 12), 198 => to_unsigned(3579, 12), 199 => to_unsigned(2519, 12), 200 => to_unsigned(225, 12), 201 => to_unsigned(351, 12), 202 => to_unsigned(3282, 12), 203 => to_unsigned(3859, 12), 204 => to_unsigned(1795, 12), 205 => to_unsigned(2481, 12), 206 => to_unsigned(2371, 12), 207 => to_unsigned(1036, 12), 208 => to_unsigned(1961, 12), 209 => to_unsigned(4043, 12), 210 => to_unsigned(2080, 12), 211 => to_unsigned(4019, 12), 212 => to_unsigned(2069, 12), 213 => to_unsigned(224, 12), 214 => to_unsigned(2696, 12), 215 => to_unsigned(351, 12), 216 => to_unsigned(2140, 12), 217 => to_unsigned(1856, 12), 218 => to_unsigned(900, 12), 219 => to_unsigned(1947, 12), 220 => to_unsigned(3886, 12), 221 => to_unsigned(267, 12), 222 => to_unsigned(2009, 12), 223 => to_unsigned(3795, 12), 224 => to_unsigned(1544, 12), 225 => to_unsigned(104, 12), 226 => to_unsigned(387, 12), 227 => to_unsigned(468, 12), 228 => to_unsigned(1033, 12), 229 => to_unsigned(1622, 12), 230 => to_unsigned(1571, 12), 231 => to_unsigned(901, 12), 232 => to_unsigned(469, 12), 233 => to_unsigned(2016, 12), 234 => to_unsigned(1084, 12), 235 => to_unsigned(2835, 12), 236 => to_unsigned(2266, 12), 237 => to_unsigned(148, 12), 238 => to_unsigned(3758, 12), 239 => to_unsigned(1620, 12), 240 => to_unsigned(2239, 12), 241 => to_unsigned(2063, 12), 242 => to_unsigned(2392, 12), 243 => to_unsigned(149, 12), 244 => to_unsigned(340, 12), 245 => to_unsigned(358, 12), 246 => to_unsigned(3661, 12), 247 => to_unsigned(3193, 12), 248 => to_unsigned(1102, 12), 249 => to_unsigned(2899, 12), 250 => to_unsigned(1799, 12), 251 => to_unsigned(921, 12), 252 => to_unsigned(1222, 12), 253 => to_unsigned(2600, 12), 254 => to_unsigned(337, 12), 255 => to_unsigned(2735, 12), 256 => to_unsigned(2743, 12), 257 => to_unsigned(2426, 12), 258 => to_unsigned(1871, 12), 259 => to_unsigned(2843, 12), 260 => to_unsigned(1617, 12), 261 => to_unsigned(3653, 12), 262 => to_unsigned(2056, 12), 263 => to_unsigned(464, 12), 264 => to_unsigned(466, 12), 265 => to_unsigned(1063, 12), 266 => to_unsigned(1603, 12), 267 => to_unsigned(2824, 12), 268 => to_unsigned(910, 12), 269 => to_unsigned(1532, 12), 270 => to_unsigned(3266, 12), 271 => to_unsigned(88, 12), 272 => to_unsigned(3629, 12), 273 => to_unsigned(2494, 12), 274 => to_unsigned(2887, 12), 275 => to_unsigned(2687, 12), 276 => to_unsigned(3851, 12), 277 => to_unsigned(740, 12), 278 => to_unsigned(2901, 12), 279 => to_unsigned(1702, 12), 280 => to_unsigned(488, 12), 281 => to_unsigned(2564, 12), 282 => to_unsigned(1704, 12), 283 => to_unsigned(2925, 12), 284 => to_unsigned(3558, 12), 285 => to_unsigned(1588, 12), 286 => to_unsigned(39, 12), 287 => to_unsigned(419, 12), 288 => to_unsigned(3218, 12), 289 => to_unsigned(3427, 12), 290 => to_unsigned(1708, 12), 291 => to_unsigned(4018, 12), 292 => to_unsigned(734, 12), 293 => to_unsigned(3414, 12), 294 => to_unsigned(3743, 12), 295 => to_unsigned(3223, 12), 296 => to_unsigned(2948, 12), 297 => to_unsigned(3088, 12), 298 => to_unsigned(1428, 12), 299 => to_unsigned(622, 12), 300 => to_unsigned(260, 12), 301 => to_unsigned(1773, 12), 302 => to_unsigned(2510, 12), 303 => to_unsigned(2944, 12), 304 => to_unsigned(1174, 12), 305 => to_unsigned(2869, 12), 306 => to_unsigned(926, 12), 307 => to_unsigned(579, 12), 308 => to_unsigned(4042, 12), 309 => to_unsigned(2992, 12), 310 => to_unsigned(241, 12), 311 => to_unsigned(3541, 12), 312 => to_unsigned(2274, 12), 313 => to_unsigned(2704, 12), 314 => to_unsigned(2103, 12), 315 => to_unsigned(3467, 12), 316 => to_unsigned(3818, 12), 317 => to_unsigned(1672, 12), 318 => to_unsigned(1400, 12), 319 => to_unsigned(3774, 12), 320 => to_unsigned(983, 12), 321 => to_unsigned(3337, 12), 322 => to_unsigned(1119, 12), 323 => to_unsigned(3922, 12), 324 => to_unsigned(71, 12), 325 => to_unsigned(2600, 12), 326 => to_unsigned(3972, 12), 327 => to_unsigned(2025, 12), 328 => to_unsigned(580, 12), 329 => to_unsigned(2943, 12), 330 => to_unsigned(131, 12), 331 => to_unsigned(2181, 12), 332 => to_unsigned(427, 12), 333 => to_unsigned(2008, 12), 334 => to_unsigned(340, 12), 335 => to_unsigned(1498, 12), 336 => to_unsigned(1300, 12), 337 => to_unsigned(2129, 12), 338 => to_unsigned(2501, 12), 339 => to_unsigned(2759, 12), 340 => to_unsigned(2948, 12), 341 => to_unsigned(2788, 12), 342 => to_unsigned(4002, 12), 343 => to_unsigned(3062, 12), 344 => to_unsigned(741, 12), 345 => to_unsigned(2660, 12), 346 => to_unsigned(3585, 12), 347 => to_unsigned(3841, 12), 348 => to_unsigned(1014, 12), 349 => to_unsigned(935, 12), 350 => to_unsigned(2675, 12), 351 => to_unsigned(2484, 12), 352 => to_unsigned(3410, 12), 353 => to_unsigned(1523, 12), 354 => to_unsigned(3192, 12), 355 => to_unsigned(3156, 12), 356 => to_unsigned(86, 12), 357 => to_unsigned(3869, 12), 358 => to_unsigned(2762, 12), 359 => to_unsigned(531, 12), 360 => to_unsigned(1319, 12), 361 => to_unsigned(708, 12), 362 => to_unsigned(1192, 12), 363 => to_unsigned(2494, 12), 364 => to_unsigned(856, 12), 365 => to_unsigned(2960, 12), 366 => to_unsigned(2026, 12), 367 => to_unsigned(3275, 12), 368 => to_unsigned(784, 12), 369 => to_unsigned(2970, 12), 370 => to_unsigned(2338, 12), 371 => to_unsigned(741, 12), 372 => to_unsigned(734, 12), 373 => to_unsigned(3224, 12), 374 => to_unsigned(894, 12), 375 => to_unsigned(2065, 12), 376 => to_unsigned(383, 12), 377 => to_unsigned(533, 12), 378 => to_unsigned(2336, 12), 379 => to_unsigned(2771, 12), 380 => to_unsigned(769, 12), 381 => to_unsigned(2450, 12), 382 => to_unsigned(621, 12), 383 => to_unsigned(189, 12), 384 => to_unsigned(2996, 12), 385 => to_unsigned(1346, 12), 386 => to_unsigned(3884, 12), 387 => to_unsigned(3197, 12), 388 => to_unsigned(2947, 12), 389 => to_unsigned(1424, 12), 390 => to_unsigned(3753, 12), 391 => to_unsigned(3127, 12), 392 => to_unsigned(996, 12), 393 => to_unsigned(3347, 12), 394 => to_unsigned(45, 12), 395 => to_unsigned(1819, 12), 396 => to_unsigned(407, 12), 397 => to_unsigned(3164, 12), 398 => to_unsigned(3675, 12), 399 => to_unsigned(2741, 12), 400 => to_unsigned(2316, 12), 401 => to_unsigned(3639, 12), 402 => to_unsigned(3667, 12), 403 => to_unsigned(2821, 12), 404 => to_unsigned(2591, 12), 405 => to_unsigned(12, 12), 406 => to_unsigned(2817, 12), 407 => to_unsigned(3445, 12), 408 => to_unsigned(977, 12), 409 => to_unsigned(3002, 12), 410 => to_unsigned(2575, 12), 411 => to_unsigned(734, 12), 412 => to_unsigned(545, 12), 413 => to_unsigned(2724, 12), 414 => to_unsigned(1405, 12), 415 => to_unsigned(2314, 12), 416 => to_unsigned(3863, 12), 417 => to_unsigned(3924, 12), 418 => to_unsigned(3410, 12), 419 => to_unsigned(2649, 12), 420 => to_unsigned(3382, 12), 421 => to_unsigned(2329, 12), 422 => to_unsigned(1061, 12), 423 => to_unsigned(572, 12), 424 => to_unsigned(2800, 12), 425 => to_unsigned(2319, 12), 426 => to_unsigned(1484, 12), 427 => to_unsigned(1051, 12), 428 => to_unsigned(3301, 12), 429 => to_unsigned(2116, 12), 430 => to_unsigned(4074, 12), 431 => to_unsigned(1553, 12), 432 => to_unsigned(1001, 12), 433 => to_unsigned(3369, 12), 434 => to_unsigned(3151, 12), 435 => to_unsigned(2476, 12), 436 => to_unsigned(2526, 12), 437 => to_unsigned(1020, 12), 438 => to_unsigned(306, 12), 439 => to_unsigned(1502, 12), 440 => to_unsigned(3116, 12), 441 => to_unsigned(1548, 12), 442 => to_unsigned(3279, 12), 443 => to_unsigned(2257, 12), 444 => to_unsigned(3801, 12), 445 => to_unsigned(477, 12), 446 => to_unsigned(2881, 12), 447 => to_unsigned(3049, 12), 448 => to_unsigned(414, 12), 449 => to_unsigned(2872, 12), 450 => to_unsigned(3561, 12), 451 => to_unsigned(3510, 12), 452 => to_unsigned(1519, 12), 453 => to_unsigned(1225, 12), 454 => to_unsigned(911, 12), 455 => to_unsigned(4012, 12), 456 => to_unsigned(1352, 12), 457 => to_unsigned(3111, 12), 458 => to_unsigned(1341, 12), 459 => to_unsigned(1549, 12), 460 => to_unsigned(389, 12), 461 => to_unsigned(1648, 12), 462 => to_unsigned(1379, 12), 463 => to_unsigned(2850, 12), 464 => to_unsigned(1528, 12), 465 => to_unsigned(425, 12), 466 => to_unsigned(3551, 12), 467 => to_unsigned(2749, 12), 468 => to_unsigned(1261, 12), 469 => to_unsigned(933, 12), 470 => to_unsigned(725, 12), 471 => to_unsigned(1398, 12), 472 => to_unsigned(2301, 12), 473 => to_unsigned(3144, 12), 474 => to_unsigned(2549, 12), 475 => to_unsigned(1429, 12), 476 => to_unsigned(2186, 12), 477 => to_unsigned(3941, 12), 478 => to_unsigned(2682, 12), 479 => to_unsigned(3125, 12), 480 => to_unsigned(2115, 12), 481 => to_unsigned(3670, 12), 482 => to_unsigned(3091, 12), 483 => to_unsigned(2575, 12), 484 => to_unsigned(152, 12), 485 => to_unsigned(2894, 12), 486 => to_unsigned(1888, 12), 487 => to_unsigned(1447, 12), 488 => to_unsigned(669, 12), 489 => to_unsigned(3508, 12), 490 => to_unsigned(2511, 12), 491 => to_unsigned(2009, 12), 492 => to_unsigned(2564, 12), 493 => to_unsigned(1077, 12), 494 => to_unsigned(3570, 12), 495 => to_unsigned(314, 12), 496 => to_unsigned(2249, 12), 497 => to_unsigned(2665, 12), 498 => to_unsigned(2773, 12), 499 => to_unsigned(2148, 12), 500 => to_unsigned(1775, 12), 501 => to_unsigned(3464, 12), 502 => to_unsigned(1001, 12), 503 => to_unsigned(2599, 12), 504 => to_unsigned(2342, 12), 505 => to_unsigned(299, 12), 506 => to_unsigned(2662, 12), 507 => to_unsigned(2520, 12), 508 => to_unsigned(4091, 12), 509 => to_unsigned(3928, 12), 510 => to_unsigned(3594, 12), 511 => to_unsigned(3252, 12), 512 => to_unsigned(1852, 12), 513 => to_unsigned(1299, 12), 514 => to_unsigned(873, 12), 515 => to_unsigned(2061, 12), 516 => to_unsigned(203, 12), 517 => to_unsigned(660, 12), 518 => to_unsigned(2136, 12), 519 => to_unsigned(400, 12), 520 => to_unsigned(1640, 12), 521 => to_unsigned(4005, 12), 522 => to_unsigned(2753, 12), 523 => to_unsigned(2041, 12), 524 => to_unsigned(2800, 12), 525 => to_unsigned(219, 12), 526 => to_unsigned(1363, 12), 527 => to_unsigned(1164, 12), 528 => to_unsigned(1859, 12), 529 => to_unsigned(825, 12), 530 => to_unsigned(2609, 12), 531 => to_unsigned(1750, 12), 532 => to_unsigned(4045, 12), 533 => to_unsigned(2205, 12), 534 => to_unsigned(1011, 12), 535 => to_unsigned(1272, 12), 536 => to_unsigned(2597, 12), 537 => to_unsigned(2737, 12), 538 => to_unsigned(4060, 12), 539 => to_unsigned(3002, 12), 540 => to_unsigned(1261, 12), 541 => to_unsigned(3867, 12), 542 => to_unsigned(3203, 12), 543 => to_unsigned(2079, 12), 544 => to_unsigned(358, 12), 545 => to_unsigned(4040, 12), 546 => to_unsigned(3013, 12), 547 => to_unsigned(3318, 12), 548 => to_unsigned(335, 12), 549 => to_unsigned(1883, 12), 550 => to_unsigned(2545, 12), 551 => to_unsigned(614, 12), 552 => to_unsigned(2157, 12), 553 => to_unsigned(626, 12), 554 => to_unsigned(224, 12), 555 => to_unsigned(2401, 12), 556 => to_unsigned(792, 12), 557 => to_unsigned(1504, 12), 558 => to_unsigned(2742, 12), 559 => to_unsigned(2514, 12), 560 => to_unsigned(3304, 12), 561 => to_unsigned(3705, 12), 562 => to_unsigned(3348, 12), 563 => to_unsigned(948, 12), 564 => to_unsigned(920, 12), 565 => to_unsigned(1538, 12), 566 => to_unsigned(2850, 12), 567 => to_unsigned(3543, 12), 568 => to_unsigned(3599, 12), 569 => to_unsigned(1306, 12), 570 => to_unsigned(145, 12), 571 => to_unsigned(607, 12), 572 => to_unsigned(1492, 12), 573 => to_unsigned(2520, 12), 574 => to_unsigned(744, 12), 575 => to_unsigned(3865, 12), 576 => to_unsigned(1195, 12), 577 => to_unsigned(1432, 12), 578 => to_unsigned(3706, 12), 579 => to_unsigned(2650, 12), 580 => to_unsigned(4092, 12), 581 => to_unsigned(3531, 12), 582 => to_unsigned(1243, 12), 583 => to_unsigned(412, 12), 584 => to_unsigned(3344, 12), 585 => to_unsigned(1318, 12), 586 => to_unsigned(3131, 12), 587 => to_unsigned(1660, 12), 588 => to_unsigned(1187, 12), 589 => to_unsigned(300, 12), 590 => to_unsigned(223, 12), 591 => to_unsigned(2547, 12), 592 => to_unsigned(2727, 12), 593 => to_unsigned(1849, 12), 594 => to_unsigned(712, 12), 595 => to_unsigned(1098, 12), 596 => to_unsigned(1445, 12), 597 => to_unsigned(2110, 12), 598 => to_unsigned(2123, 12), 599 => to_unsigned(405, 12), 600 => to_unsigned(2870, 12), 601 => to_unsigned(2946, 12), 602 => to_unsigned(489, 12), 603 => to_unsigned(1318, 12), 604 => to_unsigned(2307, 12), 605 => to_unsigned(597, 12), 606 => to_unsigned(2851, 12), 607 => to_unsigned(1251, 12), 608 => to_unsigned(3960, 12), 609 => to_unsigned(1988, 12), 610 => to_unsigned(1590, 12), 611 => to_unsigned(3635, 12), 612 => to_unsigned(269, 12), 613 => to_unsigned(3140, 12), 614 => to_unsigned(439, 12), 615 => to_unsigned(3656, 12), 616 => to_unsigned(3188, 12), 617 => to_unsigned(850, 12), 618 => to_unsigned(2015, 12), 619 => to_unsigned(1230, 12), 620 => to_unsigned(2656, 12), 621 => to_unsigned(421, 12), 622 => to_unsigned(581, 12), 623 => to_unsigned(1012, 12), 624 => to_unsigned(1641, 12), 625 => to_unsigned(1714, 12), 626 => to_unsigned(2418, 12), 627 => to_unsigned(4019, 12), 628 => to_unsigned(3860, 12), 629 => to_unsigned(1184, 12), 630 => to_unsigned(3324, 12), 631 => to_unsigned(3658, 12), 632 => to_unsigned(3892, 12), 633 => to_unsigned(2223, 12), 634 => to_unsigned(3140, 12), 635 => to_unsigned(2117, 12), 636 => to_unsigned(1436, 12), 637 => to_unsigned(1898, 12), 638 => to_unsigned(1565, 12), 639 => to_unsigned(645, 12), 640 => to_unsigned(2522, 12), 641 => to_unsigned(78, 12), 642 => to_unsigned(2998, 12), 643 => to_unsigned(2713, 12), 644 => to_unsigned(2468, 12), 645 => to_unsigned(1034, 12), 646 => to_unsigned(2754, 12), 647 => to_unsigned(3247, 12), 648 => to_unsigned(1406, 12), 649 => to_unsigned(1573, 12), 650 => to_unsigned(3783, 12), 651 => to_unsigned(2445, 12), 652 => to_unsigned(2911, 12), 653 => to_unsigned(489, 12), 654 => to_unsigned(3869, 12), 655 => to_unsigned(2181, 12), 656 => to_unsigned(1485, 12), 657 => to_unsigned(1371, 12), 658 => to_unsigned(3494, 12), 659 => to_unsigned(2576, 12), 660 => to_unsigned(798, 12), 661 => to_unsigned(3736, 12), 662 => to_unsigned(3128, 12), 663 => to_unsigned(2257, 12), 664 => to_unsigned(1331, 12), 665 => to_unsigned(225, 12), 666 => to_unsigned(1360, 12), 667 => to_unsigned(3337, 12), 668 => to_unsigned(570, 12), 669 => to_unsigned(822, 12), 670 => to_unsigned(3009, 12), 671 => to_unsigned(3118, 12), 672 => to_unsigned(2411, 12), 673 => to_unsigned(414, 12), 674 => to_unsigned(733, 12), 675 => to_unsigned(658, 12), 676 => to_unsigned(83, 12), 677 => to_unsigned(2100, 12), 678 => to_unsigned(305, 12), 679 => to_unsigned(2812, 12), 680 => to_unsigned(1742, 12), 681 => to_unsigned(2298, 12), 682 => to_unsigned(3914, 12), 683 => to_unsigned(1778, 12), 684 => to_unsigned(4045, 12), 685 => to_unsigned(2115, 12), 686 => to_unsigned(2783, 12), 687 => to_unsigned(3270, 12), 688 => to_unsigned(4023, 12), 689 => to_unsigned(1999, 12), 690 => to_unsigned(2000, 12), 691 => to_unsigned(629, 12), 692 => to_unsigned(123, 12), 693 => to_unsigned(1058, 12), 694 => to_unsigned(1743, 12), 695 => to_unsigned(2243, 12), 696 => to_unsigned(2998, 12), 697 => to_unsigned(3691, 12), 698 => to_unsigned(3090, 12), 699 => to_unsigned(2334, 12), 700 => to_unsigned(299, 12), 701 => to_unsigned(3243, 12), 702 => to_unsigned(2963, 12), 703 => to_unsigned(2481, 12), 704 => to_unsigned(69, 12), 705 => to_unsigned(2417, 12), 706 => to_unsigned(326, 12), 707 => to_unsigned(1483, 12), 708 => to_unsigned(259, 12), 709 => to_unsigned(3985, 12), 710 => to_unsigned(1939, 12), 711 => to_unsigned(1862, 12), 712 => to_unsigned(377, 12), 713 => to_unsigned(3225, 12), 714 => to_unsigned(3829, 12), 715 => to_unsigned(2648, 12), 716 => to_unsigned(2114, 12), 717 => to_unsigned(2198, 12), 718 => to_unsigned(2294, 12), 719 => to_unsigned(1873, 12), 720 => to_unsigned(3823, 12), 721 => to_unsigned(3830, 12), 722 => to_unsigned(278, 12), 723 => to_unsigned(2446, 12), 724 => to_unsigned(1636, 12), 725 => to_unsigned(1298, 12), 726 => to_unsigned(1874, 12), 727 => to_unsigned(495, 12), 728 => to_unsigned(1749, 12), 729 => to_unsigned(1938, 12), 730 => to_unsigned(1615, 12), 731 => to_unsigned(2326, 12), 732 => to_unsigned(3447, 12), 733 => to_unsigned(398, 12), 734 => to_unsigned(4038, 12), 735 => to_unsigned(2548, 12), 736 => to_unsigned(2196, 12), 737 => to_unsigned(1356, 12), 738 => to_unsigned(3110, 12), 739 => to_unsigned(3094, 12), 740 => to_unsigned(2602, 12), 741 => to_unsigned(1091, 12), 742 => to_unsigned(1207, 12), 743 => to_unsigned(3353, 12), 744 => to_unsigned(3618, 12), 745 => to_unsigned(2974, 12), 746 => to_unsigned(962, 12), 747 => to_unsigned(2667, 12), 748 => to_unsigned(2705, 12), 749 => to_unsigned(1908, 12), 750 => to_unsigned(1309, 12), 751 => to_unsigned(3096, 12), 752 => to_unsigned(3441, 12), 753 => to_unsigned(1131, 12), 754 => to_unsigned(4052, 12), 755 => to_unsigned(1852, 12), 756 => to_unsigned(2963, 12), 757 => to_unsigned(818, 12), 758 => to_unsigned(2862, 12), 759 => to_unsigned(3277, 12), 760 => to_unsigned(3503, 12), 761 => to_unsigned(3764, 12), 762 => to_unsigned(1398, 12), 763 => to_unsigned(2063, 12), 764 => to_unsigned(317, 12), 765 => to_unsigned(1771, 12), 766 => to_unsigned(2948, 12), 767 => to_unsigned(3951, 12), 768 => to_unsigned(3538, 12), 769 => to_unsigned(2979, 12), 770 => to_unsigned(2207, 12), 771 => to_unsigned(1952, 12), 772 => to_unsigned(261, 12), 773 => to_unsigned(1757, 12), 774 => to_unsigned(2427, 12), 775 => to_unsigned(1885, 12), 776 => to_unsigned(3662, 12), 777 => to_unsigned(292, 12), 778 => to_unsigned(769, 12), 779 => to_unsigned(3217, 12), 780 => to_unsigned(72, 12), 781 => to_unsigned(1560, 12), 782 => to_unsigned(2364, 12), 783 => to_unsigned(1813, 12), 784 => to_unsigned(3608, 12), 785 => to_unsigned(1588, 12), 786 => to_unsigned(1154, 12), 787 => to_unsigned(1262, 12), 788 => to_unsigned(2506, 12), 789 => to_unsigned(722, 12), 790 => to_unsigned(2670, 12), 791 => to_unsigned(434, 12), 792 => to_unsigned(4063, 12), 793 => to_unsigned(562, 12), 794 => to_unsigned(1987, 12), 795 => to_unsigned(253, 12), 796 => to_unsigned(3242, 12), 797 => to_unsigned(3899, 12), 798 => to_unsigned(3400, 12), 799 => to_unsigned(2150, 12), 800 => to_unsigned(1780, 12), 801 => to_unsigned(2039, 12), 802 => to_unsigned(813, 12), 803 => to_unsigned(1120, 12), 804 => to_unsigned(847, 12), 805 => to_unsigned(1104, 12), 806 => to_unsigned(3463, 12), 807 => to_unsigned(95, 12), 808 => to_unsigned(670, 12), 809 => to_unsigned(869, 12), 810 => to_unsigned(641, 12), 811 => to_unsigned(1044, 12), 812 => to_unsigned(2393, 12), 813 => to_unsigned(1203, 12), 814 => to_unsigned(1260, 12), 815 => to_unsigned(2677, 12), 816 => to_unsigned(1611, 12), 817 => to_unsigned(1945, 12), 818 => to_unsigned(639, 12), 819 => to_unsigned(938, 12), 820 => to_unsigned(1663, 12), 821 => to_unsigned(819, 12), 822 => to_unsigned(1190, 12), 823 => to_unsigned(1926, 12), 824 => to_unsigned(1430, 12), 825 => to_unsigned(2404, 12), 826 => to_unsigned(2209, 12), 827 => to_unsigned(2539, 12), 828 => to_unsigned(394, 12), 829 => to_unsigned(2865, 12), 830 => to_unsigned(1059, 12), 831 => to_unsigned(442, 12), 832 => to_unsigned(3131, 12), 833 => to_unsigned(3615, 12), 834 => to_unsigned(3976, 12), 835 => to_unsigned(1668, 12), 836 => to_unsigned(3593, 12), 837 => to_unsigned(3200, 12), 838 => to_unsigned(342, 12), 839 => to_unsigned(2152, 12), 840 => to_unsigned(822, 12), 841 => to_unsigned(601, 12), 842 => to_unsigned(1834, 12), 843 => to_unsigned(1830, 12), 844 => to_unsigned(1162, 12), 845 => to_unsigned(1895, 12), 846 => to_unsigned(247, 12), 847 => to_unsigned(1885, 12), 848 => to_unsigned(2349, 12), 849 => to_unsigned(2066, 12), 850 => to_unsigned(3605, 12), 851 => to_unsigned(3765, 12), 852 => to_unsigned(2442, 12), 853 => to_unsigned(1445, 12), 854 => to_unsigned(3502, 12), 855 => to_unsigned(2355, 12), 856 => to_unsigned(133, 12), 857 => to_unsigned(2550, 12), 858 => to_unsigned(3331, 12), 859 => to_unsigned(3055, 12), 860 => to_unsigned(2869, 12), 861 => to_unsigned(90, 12), 862 => to_unsigned(2756, 12), 863 => to_unsigned(2894, 12), 864 => to_unsigned(378, 12), 865 => to_unsigned(1182, 12), 866 => to_unsigned(3070, 12), 867 => to_unsigned(3906, 12), 868 => to_unsigned(63, 12), 869 => to_unsigned(4082, 12), 870 => to_unsigned(2669, 12), 871 => to_unsigned(1241, 12), 872 => to_unsigned(854, 12), 873 => to_unsigned(3003, 12), 874 => to_unsigned(499, 12), 875 => to_unsigned(1157, 12), 876 => to_unsigned(1961, 12), 877 => to_unsigned(1489, 12), 878 => to_unsigned(270, 12), 879 => to_unsigned(3674, 12), 880 => to_unsigned(3631, 12), 881 => to_unsigned(797, 12), 882 => to_unsigned(2125, 12), 883 => to_unsigned(3165, 12), 884 => to_unsigned(2715, 12), 885 => to_unsigned(1557, 12), 886 => to_unsigned(2027, 12), 887 => to_unsigned(3622, 12), 888 => to_unsigned(320, 12), 889 => to_unsigned(2611, 12), 890 => to_unsigned(810, 12), 891 => to_unsigned(3127, 12), 892 => to_unsigned(2765, 12), 893 => to_unsigned(2515, 12), 894 => to_unsigned(3346, 12), 895 => to_unsigned(2658, 12), 896 => to_unsigned(476, 12), 897 => to_unsigned(3000, 12), 898 => to_unsigned(1527, 12), 899 => to_unsigned(1184, 12), 900 => to_unsigned(1641, 12), 901 => to_unsigned(159, 12), 902 => to_unsigned(2751, 12), 903 => to_unsigned(2307, 12), 904 => to_unsigned(908, 12), 905 => to_unsigned(2102, 12), 906 => to_unsigned(1545, 12), 907 => to_unsigned(567, 12), 908 => to_unsigned(1398, 12), 909 => to_unsigned(4095, 12), 910 => to_unsigned(1822, 12), 911 => to_unsigned(1196, 12), 912 => to_unsigned(2830, 12), 913 => to_unsigned(2148, 12), 914 => to_unsigned(2153, 12), 915 => to_unsigned(2817, 12), 916 => to_unsigned(3177, 12), 917 => to_unsigned(1476, 12), 918 => to_unsigned(28, 12), 919 => to_unsigned(506, 12), 920 => to_unsigned(1039, 12), 921 => to_unsigned(1273, 12), 922 => to_unsigned(4042, 12), 923 => to_unsigned(2453, 12), 924 => to_unsigned(2074, 12), 925 => to_unsigned(2529, 12), 926 => to_unsigned(610, 12), 927 => to_unsigned(2763, 12), 928 => to_unsigned(3811, 12), 929 => to_unsigned(3833, 12), 930 => to_unsigned(892, 12), 931 => to_unsigned(1583, 12), 932 => to_unsigned(3665, 12), 933 => to_unsigned(582, 12), 934 => to_unsigned(912, 12), 935 => to_unsigned(1203, 12), 936 => to_unsigned(1408, 12), 937 => to_unsigned(2824, 12), 938 => to_unsigned(400, 12), 939 => to_unsigned(392, 12), 940 => to_unsigned(3532, 12), 941 => to_unsigned(2729, 12), 942 => to_unsigned(2466, 12), 943 => to_unsigned(2537, 12), 944 => to_unsigned(181, 12), 945 => to_unsigned(1108, 12), 946 => to_unsigned(363, 12), 947 => to_unsigned(116, 12), 948 => to_unsigned(1558, 12), 949 => to_unsigned(2469, 12), 950 => to_unsigned(1294, 12), 951 => to_unsigned(2675, 12), 952 => to_unsigned(1318, 12), 953 => to_unsigned(2848, 12), 954 => to_unsigned(2239, 12), 955 => to_unsigned(1494, 12), 956 => to_unsigned(3789, 12), 957 => to_unsigned(423, 12), 958 => to_unsigned(2700, 12), 959 => to_unsigned(239, 12), 960 => to_unsigned(2434, 12), 961 => to_unsigned(303, 12), 962 => to_unsigned(2584, 12), 963 => to_unsigned(1978, 12), 964 => to_unsigned(2842, 12), 965 => to_unsigned(2198, 12), 966 => to_unsigned(2050, 12), 967 => to_unsigned(4020, 12), 968 => to_unsigned(3870, 12), 969 => to_unsigned(1705, 12), 970 => to_unsigned(2212, 12), 971 => to_unsigned(3624, 12), 972 => to_unsigned(3276, 12), 973 => to_unsigned(1737, 12), 974 => to_unsigned(1259, 12), 975 => to_unsigned(88, 12), 976 => to_unsigned(1146, 12), 977 => to_unsigned(884, 12), 978 => to_unsigned(2839, 12), 979 => to_unsigned(885, 12), 980 => to_unsigned(3489, 12), 981 => to_unsigned(1692, 12), 982 => to_unsigned(97, 12), 983 => to_unsigned(1258, 12), 984 => to_unsigned(660, 12), 985 => to_unsigned(2118, 12), 986 => to_unsigned(498, 12), 987 => to_unsigned(1510, 12), 988 => to_unsigned(244, 12), 989 => to_unsigned(2480, 12), 990 => to_unsigned(4027, 12), 991 => to_unsigned(901, 12), 992 => to_unsigned(100, 12), 993 => to_unsigned(1938, 12), 994 => to_unsigned(933, 12), 995 => to_unsigned(734, 12), 996 => to_unsigned(1948, 12), 997 => to_unsigned(3465, 12), 998 => to_unsigned(1168, 12), 999 => to_unsigned(2549, 12), 1000 => to_unsigned(2264, 12), 1001 => to_unsigned(3412, 12), 1002 => to_unsigned(521, 12), 1003 => to_unsigned(1176, 12), 1004 => to_unsigned(569, 12), 1005 => to_unsigned(3003, 12), 1006 => to_unsigned(2515, 12), 1007 => to_unsigned(2573, 12), 1008 => to_unsigned(2076, 12), 1009 => to_unsigned(390, 12), 1010 => to_unsigned(1085, 12), 1011 => to_unsigned(2139, 12), 1012 => to_unsigned(1459, 12), 1013 => to_unsigned(2224, 12), 1014 => to_unsigned(3902, 12), 1015 => to_unsigned(3856, 12), 1016 => to_unsigned(1247, 12), 1017 => to_unsigned(1058, 12), 1018 => to_unsigned(483, 12), 1019 => to_unsigned(1246, 12), 1020 => to_unsigned(1609, 12), 1021 => to_unsigned(1304, 12), 1022 => to_unsigned(1875, 12), 1023 => to_unsigned(2923, 12), 1024 => to_unsigned(3772, 12), 1025 => to_unsigned(3828, 12), 1026 => to_unsigned(336, 12), 1027 => to_unsigned(2038, 12), 1028 => to_unsigned(4018, 12), 1029 => to_unsigned(1728, 12), 1030 => to_unsigned(1672, 12), 1031 => to_unsigned(3006, 12), 1032 => to_unsigned(3540, 12), 1033 => to_unsigned(2127, 12), 1034 => to_unsigned(2624, 12), 1035 => to_unsigned(3972, 12), 1036 => to_unsigned(651, 12), 1037 => to_unsigned(1211, 12), 1038 => to_unsigned(694, 12), 1039 => to_unsigned(965, 12), 1040 => to_unsigned(1216, 12), 1041 => to_unsigned(568, 12), 1042 => to_unsigned(451, 12), 1043 => to_unsigned(2623, 12), 1044 => to_unsigned(1096, 12), 1045 => to_unsigned(39, 12), 1046 => to_unsigned(117, 12), 1047 => to_unsigned(3588, 12), 1048 => to_unsigned(2400, 12), 1049 => to_unsigned(3970, 12), 1050 => to_unsigned(2741, 12), 1051 => to_unsigned(1130, 12), 1052 => to_unsigned(336, 12), 1053 => to_unsigned(1492, 12), 1054 => to_unsigned(3352, 12), 1055 => to_unsigned(2132, 12), 1056 => to_unsigned(1614, 12), 1057 => to_unsigned(2042, 12), 1058 => to_unsigned(1808, 12), 1059 => to_unsigned(3290, 12), 1060 => to_unsigned(4028, 12), 1061 => to_unsigned(715, 12), 1062 => to_unsigned(1012, 12), 1063 => to_unsigned(3753, 12), 1064 => to_unsigned(3741, 12), 1065 => to_unsigned(3830, 12), 1066 => to_unsigned(1603, 12), 1067 => to_unsigned(446, 12), 1068 => to_unsigned(1301, 12), 1069 => to_unsigned(3094, 12), 1070 => to_unsigned(3511, 12), 1071 => to_unsigned(1422, 12), 1072 => to_unsigned(1472, 12), 1073 => to_unsigned(35, 12), 1074 => to_unsigned(1481, 12), 1075 => to_unsigned(1343, 12), 1076 => to_unsigned(3854, 12), 1077 => to_unsigned(60, 12), 1078 => to_unsigned(1784, 12), 1079 => to_unsigned(3807, 12), 1080 => to_unsigned(210, 12), 1081 => to_unsigned(2496, 12), 1082 => to_unsigned(2646, 12), 1083 => to_unsigned(1913, 12), 1084 => to_unsigned(3181, 12), 1085 => to_unsigned(3105, 12), 1086 => to_unsigned(2358, 12), 1087 => to_unsigned(2462, 12), 1088 => to_unsigned(3087, 12), 1089 => to_unsigned(2591, 12), 1090 => to_unsigned(1964, 12), 1091 => to_unsigned(1058, 12), 1092 => to_unsigned(1161, 12), 1093 => to_unsigned(3257, 12), 1094 => to_unsigned(206, 12), 1095 => to_unsigned(1304, 12), 1096 => to_unsigned(710, 12), 1097 => to_unsigned(1624, 12), 1098 => to_unsigned(617, 12), 1099 => to_unsigned(2566, 12), 1100 => to_unsigned(2966, 12), 1101 => to_unsigned(2282, 12), 1102 => to_unsigned(2383, 12), 1103 => to_unsigned(39, 12), 1104 => to_unsigned(1205, 12), 1105 => to_unsigned(2358, 12), 1106 => to_unsigned(1472, 12), 1107 => to_unsigned(513, 12), 1108 => to_unsigned(1944, 12), 1109 => to_unsigned(3955, 12), 1110 => to_unsigned(3457, 12), 1111 => to_unsigned(1170, 12), 1112 => to_unsigned(778, 12), 1113 => to_unsigned(112, 12), 1114 => to_unsigned(3585, 12), 1115 => to_unsigned(2277, 12), 1116 => to_unsigned(1815, 12), 1117 => to_unsigned(1342, 12), 1118 => to_unsigned(3668, 12), 1119 => to_unsigned(1863, 12), 1120 => to_unsigned(1011, 12), 1121 => to_unsigned(1155, 12), 1122 => to_unsigned(26, 12), 1123 => to_unsigned(1550, 12), 1124 => to_unsigned(2051, 12), 1125 => to_unsigned(3439, 12), 1126 => to_unsigned(1449, 12), 1127 => to_unsigned(4084, 12), 1128 => to_unsigned(3496, 12), 1129 => to_unsigned(3804, 12), 1130 => to_unsigned(2198, 12), 1131 => to_unsigned(712, 12), 1132 => to_unsigned(896, 12), 1133 => to_unsigned(545, 12), 1134 => to_unsigned(337, 12), 1135 => to_unsigned(754, 12), 1136 => to_unsigned(3533, 12), 1137 => to_unsigned(380, 12), 1138 => to_unsigned(2793, 12), 1139 => to_unsigned(1813, 12), 1140 => to_unsigned(2469, 12), 1141 => to_unsigned(3914, 12), 1142 => to_unsigned(3897, 12), 1143 => to_unsigned(3796, 12), 1144 => to_unsigned(2163, 12), 1145 => to_unsigned(1847, 12), 1146 => to_unsigned(2706, 12), 1147 => to_unsigned(2360, 12), 1148 => to_unsigned(11, 12), 1149 => to_unsigned(1276, 12), 1150 => to_unsigned(1471, 12), 1151 => to_unsigned(3001, 12), 1152 => to_unsigned(2234, 12), 1153 => to_unsigned(455, 12), 1154 => to_unsigned(1508, 12), 1155 => to_unsigned(2119, 12), 1156 => to_unsigned(2733, 12), 1157 => to_unsigned(3862, 12), 1158 => to_unsigned(2255, 12), 1159 => to_unsigned(3491, 12), 1160 => to_unsigned(1652, 12), 1161 => to_unsigned(1863, 12), 1162 => to_unsigned(3989, 12), 1163 => to_unsigned(1090, 12), 1164 => to_unsigned(263, 12), 1165 => to_unsigned(3692, 12), 1166 => to_unsigned(1710, 12), 1167 => to_unsigned(536, 12), 1168 => to_unsigned(2837, 12), 1169 => to_unsigned(4092, 12), 1170 => to_unsigned(2427, 12), 1171 => to_unsigned(2385, 12), 1172 => to_unsigned(1275, 12), 1173 => to_unsigned(3350, 12), 1174 => to_unsigned(22, 12), 1175 => to_unsigned(3236, 12), 1176 => to_unsigned(1408, 12), 1177 => to_unsigned(2760, 12), 1178 => to_unsigned(2522, 12), 1179 => to_unsigned(2418, 12), 1180 => to_unsigned(3145, 12), 1181 => to_unsigned(1749, 12), 1182 => to_unsigned(1316, 12), 1183 => to_unsigned(776, 12), 1184 => to_unsigned(1346, 12), 1185 => to_unsigned(3495, 12), 1186 => to_unsigned(2871, 12), 1187 => to_unsigned(1883, 12), 1188 => to_unsigned(2628, 12), 1189 => to_unsigned(3569, 12), 1190 => to_unsigned(2302, 12), 1191 => to_unsigned(1337, 12), 1192 => to_unsigned(1605, 12), 1193 => to_unsigned(108, 12), 1194 => to_unsigned(1887, 12), 1195 => to_unsigned(2894, 12), 1196 => to_unsigned(2228, 12), 1197 => to_unsigned(3352, 12), 1198 => to_unsigned(3663, 12), 1199 => to_unsigned(2167, 12), 1200 => to_unsigned(2356, 12), 1201 => to_unsigned(3715, 12), 1202 => to_unsigned(2027, 12), 1203 => to_unsigned(3312, 12), 1204 => to_unsigned(1940, 12), 1205 => to_unsigned(2914, 12), 1206 => to_unsigned(1671, 12), 1207 => to_unsigned(866, 12), 1208 => to_unsigned(1914, 12), 1209 => to_unsigned(1685, 12), 1210 => to_unsigned(1540, 12), 1211 => to_unsigned(1366, 12), 1212 => to_unsigned(1545, 12), 1213 => to_unsigned(1778, 12), 1214 => to_unsigned(2036, 12), 1215 => to_unsigned(1749, 12), 1216 => to_unsigned(1068, 12), 1217 => to_unsigned(1086, 12), 1218 => to_unsigned(3668, 12), 1219 => to_unsigned(2947, 12), 1220 => to_unsigned(3209, 12), 1221 => to_unsigned(1497, 12), 1222 => to_unsigned(3888, 12), 1223 => to_unsigned(3262, 12), 1224 => to_unsigned(234, 12), 1225 => to_unsigned(1545, 12), 1226 => to_unsigned(2544, 12), 1227 => to_unsigned(2189, 12), 1228 => to_unsigned(2800, 12), 1229 => to_unsigned(2830, 12), 1230 => to_unsigned(2246, 12), 1231 => to_unsigned(675, 12), 1232 => to_unsigned(1753, 12), 1233 => to_unsigned(594, 12), 1234 => to_unsigned(1772, 12), 1235 => to_unsigned(3465, 12), 1236 => to_unsigned(859, 12), 1237 => to_unsigned(2871, 12), 1238 => to_unsigned(772, 12), 1239 => to_unsigned(1793, 12), 1240 => to_unsigned(1379, 12), 1241 => to_unsigned(3975, 12), 1242 => to_unsigned(448, 12), 1243 => to_unsigned(2871, 12), 1244 => to_unsigned(3710, 12), 1245 => to_unsigned(3143, 12), 1246 => to_unsigned(3437, 12), 1247 => to_unsigned(2397, 12), 1248 => to_unsigned(2628, 12), 1249 => to_unsigned(2822, 12), 1250 => to_unsigned(592, 12), 1251 => to_unsigned(987, 12), 1252 => to_unsigned(2627, 12), 1253 => to_unsigned(2091, 12), 1254 => to_unsigned(2625, 12), 1255 => to_unsigned(2607, 12), 1256 => to_unsigned(2658, 12), 1257 => to_unsigned(494, 12), 1258 => to_unsigned(2961, 12), 1259 => to_unsigned(1317, 12), 1260 => to_unsigned(1773, 12), 1261 => to_unsigned(2874, 12), 1262 => to_unsigned(3621, 12), 1263 => to_unsigned(1328, 12), 1264 => to_unsigned(2043, 12), 1265 => to_unsigned(934, 12), 1266 => to_unsigned(1005, 12), 1267 => to_unsigned(2605, 12), 1268 => to_unsigned(2554, 12), 1269 => to_unsigned(1060, 12), 1270 => to_unsigned(343, 12), 1271 => to_unsigned(761, 12), 1272 => to_unsigned(666, 12), 1273 => to_unsigned(1953, 12), 1274 => to_unsigned(1834, 12), 1275 => to_unsigned(2931, 12), 1276 => to_unsigned(1247, 12), 1277 => to_unsigned(209, 12), 1278 => to_unsigned(1429, 12), 1279 => to_unsigned(1141, 12), 1280 => to_unsigned(748, 12), 1281 => to_unsigned(3999, 12), 1282 => to_unsigned(907, 12), 1283 => to_unsigned(1858, 12), 1284 => to_unsigned(298, 12), 1285 => to_unsigned(1633, 12), 1286 => to_unsigned(2838, 12), 1287 => to_unsigned(3467, 12), 1288 => to_unsigned(2536, 12), 1289 => to_unsigned(1531, 12), 1290 => to_unsigned(2989, 12), 1291 => to_unsigned(2736, 12), 1292 => to_unsigned(1886, 12), 1293 => to_unsigned(3859, 12), 1294 => to_unsigned(1318, 12), 1295 => to_unsigned(2918, 12), 1296 => to_unsigned(3012, 12), 1297 => to_unsigned(2421, 12), 1298 => to_unsigned(269, 12), 1299 => to_unsigned(2861, 12), 1300 => to_unsigned(3696, 12), 1301 => to_unsigned(3567, 12), 1302 => to_unsigned(1114, 12), 1303 => to_unsigned(4090, 12), 1304 => to_unsigned(1397, 12), 1305 => to_unsigned(38, 12), 1306 => to_unsigned(350, 12), 1307 => to_unsigned(1550, 12), 1308 => to_unsigned(3516, 12), 1309 => to_unsigned(611, 12), 1310 => to_unsigned(607, 12), 1311 => to_unsigned(3254, 12), 1312 => to_unsigned(3274, 12), 1313 => to_unsigned(3683, 12), 1314 => to_unsigned(2026, 12), 1315 => to_unsigned(2510, 12), 1316 => to_unsigned(1299, 12), 1317 => to_unsigned(3497, 12), 1318 => to_unsigned(1819, 12), 1319 => to_unsigned(490, 12), 1320 => to_unsigned(389, 12), 1321 => to_unsigned(439, 12), 1322 => to_unsigned(2776, 12), 1323 => to_unsigned(3656, 12), 1324 => to_unsigned(4078, 12), 1325 => to_unsigned(1811, 12), 1326 => to_unsigned(2341, 12), 1327 => to_unsigned(3405, 12), 1328 => to_unsigned(2270, 12), 1329 => to_unsigned(2927, 12), 1330 => to_unsigned(3072, 12), 1331 => to_unsigned(651, 12), 1332 => to_unsigned(1058, 12), 1333 => to_unsigned(1036, 12), 1334 => to_unsigned(3635, 12), 1335 => to_unsigned(1691, 12), 1336 => to_unsigned(1651, 12), 1337 => to_unsigned(377, 12), 1338 => to_unsigned(679, 12), 1339 => to_unsigned(3616, 12), 1340 => to_unsigned(2459, 12), 1341 => to_unsigned(2822, 12), 1342 => to_unsigned(2742, 12), 1343 => to_unsigned(1628, 12), 1344 => to_unsigned(1297, 12), 1345 => to_unsigned(2756, 12), 1346 => to_unsigned(2200, 12), 1347 => to_unsigned(3803, 12), 1348 => to_unsigned(1042, 12), 1349 => to_unsigned(1106, 12), 1350 => to_unsigned(990, 12), 1351 => to_unsigned(3973, 12), 1352 => to_unsigned(1182, 12), 1353 => to_unsigned(1768, 12), 1354 => to_unsigned(1535, 12), 1355 => to_unsigned(2635, 12), 1356 => to_unsigned(953, 12), 1357 => to_unsigned(2021, 12), 1358 => to_unsigned(2110, 12), 1359 => to_unsigned(3388, 12), 1360 => to_unsigned(439, 12), 1361 => to_unsigned(734, 12), 1362 => to_unsigned(129, 12), 1363 => to_unsigned(2326, 12), 1364 => to_unsigned(1541, 12), 1365 => to_unsigned(228, 12), 1366 => to_unsigned(1746, 12), 1367 => to_unsigned(2818, 12), 1368 => to_unsigned(1328, 12), 1369 => to_unsigned(46, 12), 1370 => to_unsigned(498, 12), 1371 => to_unsigned(427, 12), 1372 => to_unsigned(445, 12), 1373 => to_unsigned(521, 12), 1374 => to_unsigned(2466, 12), 1375 => to_unsigned(3953, 12), 1376 => to_unsigned(841, 12), 1377 => to_unsigned(2955, 12), 1378 => to_unsigned(1447, 12), 1379 => to_unsigned(2599, 12), 1380 => to_unsigned(993, 12), 1381 => to_unsigned(22, 12), 1382 => to_unsigned(1512, 12), 1383 => to_unsigned(2484, 12), 1384 => to_unsigned(1779, 12), 1385 => to_unsigned(2153, 12), 1386 => to_unsigned(449, 12), 1387 => to_unsigned(543, 12), 1388 => to_unsigned(2045, 12), 1389 => to_unsigned(1555, 12), 1390 => to_unsigned(1336, 12), 1391 => to_unsigned(1562, 12), 1392 => to_unsigned(3836, 12), 1393 => to_unsigned(190, 12), 1394 => to_unsigned(2068, 12), 1395 => to_unsigned(997, 12), 1396 => to_unsigned(2340, 12), 1397 => to_unsigned(1857, 12), 1398 => to_unsigned(1901, 12), 1399 => to_unsigned(1298, 12), 1400 => to_unsigned(71, 12), 1401 => to_unsigned(1635, 12), 1402 => to_unsigned(577, 12), 1403 => to_unsigned(248, 12), 1404 => to_unsigned(3707, 12), 1405 => to_unsigned(2490, 12), 1406 => to_unsigned(2732, 12), 1407 => to_unsigned(221, 12), 1408 => to_unsigned(1868, 12), 1409 => to_unsigned(1016, 12), 1410 => to_unsigned(2622, 12), 1411 => to_unsigned(2231, 12), 1412 => to_unsigned(3861, 12), 1413 => to_unsigned(2466, 12), 1414 => to_unsigned(2469, 12), 1415 => to_unsigned(194, 12), 1416 => to_unsigned(2848, 12), 1417 => to_unsigned(888, 12), 1418 => to_unsigned(1399, 12), 1419 => to_unsigned(3318, 12), 1420 => to_unsigned(4036, 12), 1421 => to_unsigned(878, 12), 1422 => to_unsigned(1246, 12), 1423 => to_unsigned(2741, 12), 1424 => to_unsigned(2292, 12), 1425 => to_unsigned(2483, 12), 1426 => to_unsigned(3603, 12), 1427 => to_unsigned(1345, 12), 1428 => to_unsigned(1259, 12), 1429 => to_unsigned(281, 12), 1430 => to_unsigned(1072, 12), 1431 => to_unsigned(3036, 12), 1432 => to_unsigned(3978, 12), 1433 => to_unsigned(2700, 12), 1434 => to_unsigned(3917, 12), 1435 => to_unsigned(1470, 12), 1436 => to_unsigned(3142, 12), 1437 => to_unsigned(1890, 12), 1438 => to_unsigned(574, 12), 1439 => to_unsigned(2472, 12), 1440 => to_unsigned(141, 12), 1441 => to_unsigned(594, 12), 1442 => to_unsigned(3445, 12), 1443 => to_unsigned(3020, 12), 1444 => to_unsigned(3996, 12), 1445 => to_unsigned(632, 12), 1446 => to_unsigned(2063, 12), 1447 => to_unsigned(1547, 12), 1448 => to_unsigned(1729, 12), 1449 => to_unsigned(874, 12), 1450 => to_unsigned(1548, 12), 1451 => to_unsigned(649, 12), 1452 => to_unsigned(2463, 12), 1453 => to_unsigned(2707, 12), 1454 => to_unsigned(1321, 12), 1455 => to_unsigned(3569, 12), 1456 => to_unsigned(3670, 12), 1457 => to_unsigned(3487, 12), 1458 => to_unsigned(2394, 12), 1459 => to_unsigned(3557, 12), 1460 => to_unsigned(2207, 12), 1461 => to_unsigned(2797, 12), 1462 => to_unsigned(3113, 12), 1463 => to_unsigned(1055, 12), 1464 => to_unsigned(1406, 12), 1465 => to_unsigned(2515, 12), 1466 => to_unsigned(531, 12), 1467 => to_unsigned(3820, 12), 1468 => to_unsigned(3304, 12), 1469 => to_unsigned(2136, 12), 1470 => to_unsigned(1326, 12), 1471 => to_unsigned(684, 12), 1472 => to_unsigned(1580, 12), 1473 => to_unsigned(3213, 12), 1474 => to_unsigned(3882, 12), 1475 => to_unsigned(3871, 12), 1476 => to_unsigned(2150, 12), 1477 => to_unsigned(3206, 12), 1478 => to_unsigned(748, 12), 1479 => to_unsigned(2504, 12), 1480 => to_unsigned(973, 12), 1481 => to_unsigned(2737, 12), 1482 => to_unsigned(743, 12), 1483 => to_unsigned(2220, 12), 1484 => to_unsigned(1466, 12), 1485 => to_unsigned(2499, 12), 1486 => to_unsigned(376, 12), 1487 => to_unsigned(3498, 12), 1488 => to_unsigned(3274, 12), 1489 => to_unsigned(582, 12), 1490 => to_unsigned(148, 12), 1491 => to_unsigned(1416, 12), 1492 => to_unsigned(3356, 12), 1493 => to_unsigned(1205, 12), 1494 => to_unsigned(208, 12), 1495 => to_unsigned(3483, 12), 1496 => to_unsigned(3578, 12), 1497 => to_unsigned(1466, 12), 1498 => to_unsigned(1443, 12), 1499 => to_unsigned(1645, 12), 1500 => to_unsigned(3736, 12), 1501 => to_unsigned(2817, 12), 1502 => to_unsigned(641, 12), 1503 => to_unsigned(820, 12), 1504 => to_unsigned(3774, 12), 1505 => to_unsigned(1141, 12), 1506 => to_unsigned(3225, 12), 1507 => to_unsigned(3226, 12), 1508 => to_unsigned(1985, 12), 1509 => to_unsigned(3019, 12), 1510 => to_unsigned(1120, 12), 1511 => to_unsigned(1228, 12), 1512 => to_unsigned(698, 12), 1513 => to_unsigned(3164, 12), 1514 => to_unsigned(3393, 12), 1515 => to_unsigned(454, 12), 1516 => to_unsigned(2891, 12), 1517 => to_unsigned(71, 12), 1518 => to_unsigned(3269, 12), 1519 => to_unsigned(3084, 12), 1520 => to_unsigned(1056, 12), 1521 => to_unsigned(3162, 12), 1522 => to_unsigned(2799, 12), 1523 => to_unsigned(2752, 12), 1524 => to_unsigned(597, 12), 1525 => to_unsigned(4056, 12), 1526 => to_unsigned(1869, 12), 1527 => to_unsigned(294, 12), 1528 => to_unsigned(2328, 12), 1529 => to_unsigned(1394, 12), 1530 => to_unsigned(2478, 12), 1531 => to_unsigned(2149, 12), 1532 => to_unsigned(2633, 12), 1533 => to_unsigned(1567, 12), 1534 => to_unsigned(2737, 12), 1535 => to_unsigned(2052, 12), 1536 => to_unsigned(347, 12), 1537 => to_unsigned(1725, 12), 1538 => to_unsigned(1052, 12), 1539 => to_unsigned(1872, 12), 1540 => to_unsigned(1716, 12), 1541 => to_unsigned(3735, 12), 1542 => to_unsigned(1363, 12), 1543 => to_unsigned(3439, 12), 1544 => to_unsigned(200, 12), 1545 => to_unsigned(368, 12), 1546 => to_unsigned(2580, 12), 1547 => to_unsigned(307, 12), 1548 => to_unsigned(1783, 12), 1549 => to_unsigned(3325, 12), 1550 => to_unsigned(557, 12), 1551 => to_unsigned(1514, 12), 1552 => to_unsigned(1560, 12), 1553 => to_unsigned(3772, 12), 1554 => to_unsigned(1651, 12), 1555 => to_unsigned(278, 12), 1556 => to_unsigned(1555, 12), 1557 => to_unsigned(1435, 12), 1558 => to_unsigned(1410, 12), 1559 => to_unsigned(2685, 12), 1560 => to_unsigned(3890, 12), 1561 => to_unsigned(2038, 12), 1562 => to_unsigned(852, 12), 1563 => to_unsigned(3277, 12), 1564 => to_unsigned(4095, 12), 1565 => to_unsigned(4003, 12), 1566 => to_unsigned(1913, 12), 1567 => to_unsigned(294, 12), 1568 => to_unsigned(976, 12), 1569 => to_unsigned(3757, 12), 1570 => to_unsigned(1184, 12), 1571 => to_unsigned(2242, 12), 1572 => to_unsigned(530, 12), 1573 => to_unsigned(3289, 12), 1574 => to_unsigned(2987, 12), 1575 => to_unsigned(515, 12), 1576 => to_unsigned(1171, 12), 1577 => to_unsigned(3888, 12), 1578 => to_unsigned(312, 12), 1579 => to_unsigned(3985, 12), 1580 => to_unsigned(1812, 12), 1581 => to_unsigned(3029, 12), 1582 => to_unsigned(424, 12), 1583 => to_unsigned(4073, 12), 1584 => to_unsigned(2096, 12), 1585 => to_unsigned(4038, 12), 1586 => to_unsigned(3344, 12), 1587 => to_unsigned(1217, 12), 1588 => to_unsigned(2508, 12), 1589 => to_unsigned(1966, 12), 1590 => to_unsigned(2229, 12), 1591 => to_unsigned(272, 12), 1592 => to_unsigned(2709, 12), 1593 => to_unsigned(2802, 12), 1594 => to_unsigned(3405, 12), 1595 => to_unsigned(514, 12), 1596 => to_unsigned(195, 12), 1597 => to_unsigned(1937, 12), 1598 => to_unsigned(1865, 12), 1599 => to_unsigned(3639, 12), 1600 => to_unsigned(804, 12), 1601 => to_unsigned(2317, 12), 1602 => to_unsigned(3089, 12), 1603 => to_unsigned(1981, 12), 1604 => to_unsigned(692, 12), 1605 => to_unsigned(380, 12), 1606 => to_unsigned(2465, 12), 1607 => to_unsigned(962, 12), 1608 => to_unsigned(2325, 12), 1609 => to_unsigned(433, 12), 1610 => to_unsigned(4070, 12), 1611 => to_unsigned(1970, 12), 1612 => to_unsigned(1262, 12), 1613 => to_unsigned(3986, 12), 1614 => to_unsigned(218, 12), 1615 => to_unsigned(1100, 12), 1616 => to_unsigned(4032, 12), 1617 => to_unsigned(575, 12), 1618 => to_unsigned(2549, 12), 1619 => to_unsigned(1167, 12), 1620 => to_unsigned(2676, 12), 1621 => to_unsigned(1542, 12), 1622 => to_unsigned(1799, 12), 1623 => to_unsigned(307, 12), 1624 => to_unsigned(3172, 12), 1625 => to_unsigned(3960, 12), 1626 => to_unsigned(559, 12), 1627 => to_unsigned(3089, 12), 1628 => to_unsigned(390, 12), 1629 => to_unsigned(3729, 12), 1630 => to_unsigned(452, 12), 1631 => to_unsigned(3087, 12), 1632 => to_unsigned(720, 12), 1633 => to_unsigned(3825, 12), 1634 => to_unsigned(2602, 12), 1635 => to_unsigned(3022, 12), 1636 => to_unsigned(709, 12), 1637 => to_unsigned(3788, 12), 1638 => to_unsigned(3539, 12), 1639 => to_unsigned(3685, 12), 1640 => to_unsigned(3918, 12), 1641 => to_unsigned(2518, 12), 1642 => to_unsigned(2282, 12), 1643 => to_unsigned(2245, 12), 1644 => to_unsigned(2241, 12), 1645 => to_unsigned(1397, 12), 1646 => to_unsigned(1603, 12), 1647 => to_unsigned(1982, 12), 1648 => to_unsigned(3405, 12), 1649 => to_unsigned(511, 12), 1650 => to_unsigned(1210, 12), 1651 => to_unsigned(3353, 12), 1652 => to_unsigned(255, 12), 1653 => to_unsigned(1798, 12), 1654 => to_unsigned(3214, 12), 1655 => to_unsigned(2829, 12), 1656 => to_unsigned(1741, 12), 1657 => to_unsigned(989, 12), 1658 => to_unsigned(3456, 12), 1659 => to_unsigned(959, 12), 1660 => to_unsigned(1129, 12), 1661 => to_unsigned(347, 12), 1662 => to_unsigned(606, 12), 1663 => to_unsigned(1053, 12), 1664 => to_unsigned(1429, 12), 1665 => to_unsigned(532, 12), 1666 => to_unsigned(1435, 12), 1667 => to_unsigned(4005, 12), 1668 => to_unsigned(3604, 12), 1669 => to_unsigned(177, 12), 1670 => to_unsigned(3289, 12), 1671 => to_unsigned(2168, 12), 1672 => to_unsigned(629, 12), 1673 => to_unsigned(3875, 12), 1674 => to_unsigned(52, 12), 1675 => to_unsigned(3180, 12), 1676 => to_unsigned(2146, 12), 1677 => to_unsigned(760, 12), 1678 => to_unsigned(2432, 12), 1679 => to_unsigned(2128, 12), 1680 => to_unsigned(3865, 12), 1681 => to_unsigned(3097, 12), 1682 => to_unsigned(2401, 12), 1683 => to_unsigned(3758, 12), 1684 => to_unsigned(462, 12), 1685 => to_unsigned(2866, 12), 1686 => to_unsigned(3307, 12), 1687 => to_unsigned(3519, 12), 1688 => to_unsigned(2244, 12), 1689 => to_unsigned(263, 12), 1690 => to_unsigned(3082, 12), 1691 => to_unsigned(35, 12), 1692 => to_unsigned(4018, 12), 1693 => to_unsigned(2876, 12), 1694 => to_unsigned(3273, 12), 1695 => to_unsigned(3969, 12), 1696 => to_unsigned(1526, 12), 1697 => to_unsigned(454, 12), 1698 => to_unsigned(1549, 12), 1699 => to_unsigned(3271, 12), 1700 => to_unsigned(301, 12), 1701 => to_unsigned(1457, 12), 1702 => to_unsigned(3226, 12), 1703 => to_unsigned(340, 12), 1704 => to_unsigned(2947, 12), 1705 => to_unsigned(2372, 12), 1706 => to_unsigned(3558, 12), 1707 => to_unsigned(3030, 12), 1708 => to_unsigned(1698, 12), 1709 => to_unsigned(584, 12), 1710 => to_unsigned(3946, 12), 1711 => to_unsigned(1667, 12), 1712 => to_unsigned(1216, 12), 1713 => to_unsigned(2814, 12), 1714 => to_unsigned(2646, 12), 1715 => to_unsigned(513, 12), 1716 => to_unsigned(1575, 12), 1717 => to_unsigned(3411, 12), 1718 => to_unsigned(2225, 12), 1719 => to_unsigned(1460, 12), 1720 => to_unsigned(1093, 12), 1721 => to_unsigned(2474, 12), 1722 => to_unsigned(3904, 12), 1723 => to_unsigned(3371, 12), 1724 => to_unsigned(1450, 12), 1725 => to_unsigned(3596, 12), 1726 => to_unsigned(1878, 12), 1727 => to_unsigned(1386, 12), 1728 => to_unsigned(2990, 12), 1729 => to_unsigned(558, 12), 1730 => to_unsigned(3658, 12), 1731 => to_unsigned(3365, 12), 1732 => to_unsigned(3776, 12), 1733 => to_unsigned(755, 12), 1734 => to_unsigned(290, 12), 1735 => to_unsigned(648, 12), 1736 => to_unsigned(2128, 12), 1737 => to_unsigned(1086, 12), 1738 => to_unsigned(1358, 12), 1739 => to_unsigned(2454, 12), 1740 => to_unsigned(2149, 12), 1741 => to_unsigned(4053, 12), 1742 => to_unsigned(563, 12), 1743 => to_unsigned(3626, 12), 1744 => to_unsigned(1158, 12), 1745 => to_unsigned(162, 12), 1746 => to_unsigned(1543, 12), 1747 => to_unsigned(3990, 12), 1748 => to_unsigned(584, 12), 1749 => to_unsigned(3593, 12), 1750 => to_unsigned(1287, 12), 1751 => to_unsigned(3383, 12), 1752 => to_unsigned(1886, 12), 1753 => to_unsigned(2792, 12), 1754 => to_unsigned(1042, 12), 1755 => to_unsigned(1548, 12), 1756 => to_unsigned(191, 12), 1757 => to_unsigned(3304, 12), 1758 => to_unsigned(1436, 12), 1759 => to_unsigned(4073, 12), 1760 => to_unsigned(2087, 12), 1761 => to_unsigned(3263, 12), 1762 => to_unsigned(1906, 12), 1763 => to_unsigned(1674, 12), 1764 => to_unsigned(2754, 12), 1765 => to_unsigned(1010, 12), 1766 => to_unsigned(355, 12), 1767 => to_unsigned(2114, 12), 1768 => to_unsigned(3577, 12), 1769 => to_unsigned(220, 12), 1770 => to_unsigned(1382, 12), 1771 => to_unsigned(2065, 12), 1772 => to_unsigned(922, 12), 1773 => to_unsigned(3636, 12), 1774 => to_unsigned(1706, 12), 1775 => to_unsigned(922, 12), 1776 => to_unsigned(2099, 12), 1777 => to_unsigned(1738, 12), 1778 => to_unsigned(3228, 12), 1779 => to_unsigned(733, 12), 1780 => to_unsigned(3174, 12), 1781 => to_unsigned(569, 12), 1782 => to_unsigned(3676, 12), 1783 => to_unsigned(3398, 12), 1784 => to_unsigned(334, 12), 1785 => to_unsigned(1275, 12), 1786 => to_unsigned(2028, 12), 1787 => to_unsigned(2504, 12), 1788 => to_unsigned(926, 12), 1789 => to_unsigned(2567, 12), 1790 => to_unsigned(2516, 12), 1791 => to_unsigned(1882, 12), 1792 => to_unsigned(221, 12), 1793 => to_unsigned(458, 12), 1794 => to_unsigned(764, 12), 1795 => to_unsigned(678, 12), 1796 => to_unsigned(3095, 12), 1797 => to_unsigned(1496, 12), 1798 => to_unsigned(3889, 12), 1799 => to_unsigned(604, 12), 1800 => to_unsigned(3457, 12), 1801 => to_unsigned(909, 12), 1802 => to_unsigned(1218, 12), 1803 => to_unsigned(1321, 12), 1804 => to_unsigned(560, 12), 1805 => to_unsigned(172, 12), 1806 => to_unsigned(2299, 12), 1807 => to_unsigned(4046, 12), 1808 => to_unsigned(1129, 12), 1809 => to_unsigned(2835, 12), 1810 => to_unsigned(3556, 12), 1811 => to_unsigned(1631, 12), 1812 => to_unsigned(1647, 12), 1813 => to_unsigned(283, 12), 1814 => to_unsigned(2782, 12), 1815 => to_unsigned(1, 12), 1816 => to_unsigned(1105, 12), 1817 => to_unsigned(2453, 12), 1818 => to_unsigned(457, 12), 1819 => to_unsigned(1807, 12), 1820 => to_unsigned(3164, 12), 1821 => to_unsigned(3091, 12), 1822 => to_unsigned(956, 12), 1823 => to_unsigned(1173, 12), 1824 => to_unsigned(1110, 12), 1825 => to_unsigned(1508, 12), 1826 => to_unsigned(1400, 12), 1827 => to_unsigned(3216, 12), 1828 => to_unsigned(1395, 12), 1829 => to_unsigned(2738, 12), 1830 => to_unsigned(235, 12), 1831 => to_unsigned(3429, 12), 1832 => to_unsigned(2393, 12), 1833 => to_unsigned(2554, 12), 1834 => to_unsigned(1268, 12), 1835 => to_unsigned(93, 12), 1836 => to_unsigned(1743, 12), 1837 => to_unsigned(2201, 12), 1838 => to_unsigned(1663, 12), 1839 => to_unsigned(2346, 12), 1840 => to_unsigned(3900, 12), 1841 => to_unsigned(3071, 12), 1842 => to_unsigned(2145, 12), 1843 => to_unsigned(3264, 12), 1844 => to_unsigned(1278, 12), 1845 => to_unsigned(3058, 12), 1846 => to_unsigned(1367, 12), 1847 => to_unsigned(3386, 12), 1848 => to_unsigned(1731, 12), 1849 => to_unsigned(2007, 12), 1850 => to_unsigned(2718, 12), 1851 => to_unsigned(350, 12), 1852 => to_unsigned(188, 12), 1853 => to_unsigned(113, 12), 1854 => to_unsigned(3804, 12), 1855 => to_unsigned(1859, 12), 1856 => to_unsigned(2601, 12), 1857 => to_unsigned(2826, 12), 1858 => to_unsigned(46, 12), 1859 => to_unsigned(2213, 12), 1860 => to_unsigned(2935, 12), 1861 => to_unsigned(2051, 12), 1862 => to_unsigned(1510, 12), 1863 => to_unsigned(2470, 12), 1864 => to_unsigned(2836, 12), 1865 => to_unsigned(2752, 12), 1866 => to_unsigned(3809, 12), 1867 => to_unsigned(4077, 12), 1868 => to_unsigned(2746, 12), 1869 => to_unsigned(750, 12), 1870 => to_unsigned(633, 12), 1871 => to_unsigned(883, 12), 1872 => to_unsigned(2606, 12), 1873 => to_unsigned(392, 12), 1874 => to_unsigned(3595, 12), 1875 => to_unsigned(1385, 12), 1876 => to_unsigned(3537, 12), 1877 => to_unsigned(3785, 12), 1878 => to_unsigned(549, 12), 1879 => to_unsigned(778, 12), 1880 => to_unsigned(3233, 12), 1881 => to_unsigned(3140, 12), 1882 => to_unsigned(234, 12), 1883 => to_unsigned(3983, 12), 1884 => to_unsigned(218, 12), 1885 => to_unsigned(98, 12), 1886 => to_unsigned(3209, 12), 1887 => to_unsigned(338, 12), 1888 => to_unsigned(2579, 12), 1889 => to_unsigned(128, 12), 1890 => to_unsigned(2464, 12), 1891 => to_unsigned(720, 12), 1892 => to_unsigned(3745, 12), 1893 => to_unsigned(2278, 12), 1894 => to_unsigned(2551, 12), 1895 => to_unsigned(664, 12), 1896 => to_unsigned(313, 12), 1897 => to_unsigned(1818, 12), 1898 => to_unsigned(2018, 12), 1899 => to_unsigned(396, 12), 1900 => to_unsigned(130, 12), 1901 => to_unsigned(3621, 12), 1902 => to_unsigned(2188, 12), 1903 => to_unsigned(802, 12), 1904 => to_unsigned(2777, 12), 1905 => to_unsigned(1395, 12), 1906 => to_unsigned(2707, 12), 1907 => to_unsigned(692, 12), 1908 => to_unsigned(13, 12), 1909 => to_unsigned(769, 12), 1910 => to_unsigned(580, 12), 1911 => to_unsigned(1108, 12), 1912 => to_unsigned(1306, 12), 1913 => to_unsigned(2137, 12), 1914 => to_unsigned(407, 12), 1915 => to_unsigned(2789, 12), 1916 => to_unsigned(3238, 12), 1917 => to_unsigned(2623, 12), 1918 => to_unsigned(1972, 12), 1919 => to_unsigned(3980, 12), 1920 => to_unsigned(1110, 12), 1921 => to_unsigned(1950, 12), 1922 => to_unsigned(203, 12), 1923 => to_unsigned(4011, 12), 1924 => to_unsigned(245, 12), 1925 => to_unsigned(2108, 12), 1926 => to_unsigned(2363, 12), 1927 => to_unsigned(1240, 12), 1928 => to_unsigned(3613, 12), 1929 => to_unsigned(831, 12), 1930 => to_unsigned(1726, 12), 1931 => to_unsigned(3791, 12), 1932 => to_unsigned(236, 12), 1933 => to_unsigned(479, 12), 1934 => to_unsigned(3549, 12), 1935 => to_unsigned(3715, 12), 1936 => to_unsigned(669, 12), 1937 => to_unsigned(1398, 12), 1938 => to_unsigned(3297, 12), 1939 => to_unsigned(3523, 12), 1940 => to_unsigned(2844, 12), 1941 => to_unsigned(873, 12), 1942 => to_unsigned(3025, 12), 1943 => to_unsigned(1391, 12), 1944 => to_unsigned(3071, 12), 1945 => to_unsigned(1619, 12), 1946 => to_unsigned(1955, 12), 1947 => to_unsigned(3483, 12), 1948 => to_unsigned(213, 12), 1949 => to_unsigned(247, 12), 1950 => to_unsigned(1967, 12), 1951 => to_unsigned(2035, 12), 1952 => to_unsigned(328, 12), 1953 => to_unsigned(258, 12), 1954 => to_unsigned(3382, 12), 1955 => to_unsigned(965, 12), 1956 => to_unsigned(4057, 12), 1957 => to_unsigned(2339, 12), 1958 => to_unsigned(3081, 12), 1959 => to_unsigned(1687, 12), 1960 => to_unsigned(2672, 12), 1961 => to_unsigned(2127, 12), 1962 => to_unsigned(1241, 12), 1963 => to_unsigned(3925, 12), 1964 => to_unsigned(108, 12), 1965 => to_unsigned(2103, 12), 1966 => to_unsigned(3457, 12), 1967 => to_unsigned(1371, 12), 1968 => to_unsigned(2482, 12), 1969 => to_unsigned(3036, 12), 1970 => to_unsigned(372, 12), 1971 => to_unsigned(3914, 12), 1972 => to_unsigned(2035, 12), 1973 => to_unsigned(343, 12), 1974 => to_unsigned(2498, 12), 1975 => to_unsigned(2130, 12), 1976 => to_unsigned(1187, 12), 1977 => to_unsigned(2950, 12), 1978 => to_unsigned(1899, 12), 1979 => to_unsigned(842, 12), 1980 => to_unsigned(1127, 12), 1981 => to_unsigned(1766, 12), 1982 => to_unsigned(3050, 12), 1983 => to_unsigned(2275, 12), 1984 => to_unsigned(3427, 12), 1985 => to_unsigned(3614, 12), 1986 => to_unsigned(775, 12), 1987 => to_unsigned(2974, 12), 1988 => to_unsigned(2388, 12), 1989 => to_unsigned(1773, 12), 1990 => to_unsigned(1010, 12), 1991 => to_unsigned(404, 12), 1992 => to_unsigned(1142, 12), 1993 => to_unsigned(1901, 12), 1994 => to_unsigned(1569, 12), 1995 => to_unsigned(3053, 12), 1996 => to_unsigned(518, 12), 1997 => to_unsigned(918, 12), 1998 => to_unsigned(3447, 12), 1999 => to_unsigned(3539, 12), 2000 => to_unsigned(3896, 12), 2001 => to_unsigned(33, 12), 2002 => to_unsigned(278, 12), 2003 => to_unsigned(444, 12), 2004 => to_unsigned(3533, 12), 2005 => to_unsigned(383, 12), 2006 => to_unsigned(2740, 12), 2007 => to_unsigned(2527, 12), 2008 => to_unsigned(2516, 12), 2009 => to_unsigned(1678, 12), 2010 => to_unsigned(286, 12), 2011 => to_unsigned(2064, 12), 2012 => to_unsigned(2118, 12), 2013 => to_unsigned(1680, 12), 2014 => to_unsigned(1057, 12), 2015 => to_unsigned(126, 12), 2016 => to_unsigned(2406, 12), 2017 => to_unsigned(2683, 12), 2018 => to_unsigned(3871, 12), 2019 => to_unsigned(182, 12), 2020 => to_unsigned(1361, 12), 2021 => to_unsigned(3326, 12), 2022 => to_unsigned(1796, 12), 2023 => to_unsigned(2401, 12), 2024 => to_unsigned(1895, 12), 2025 => to_unsigned(3383, 12), 2026 => to_unsigned(3279, 12), 2027 => to_unsigned(4015, 12), 2028 => to_unsigned(3911, 12), 2029 => to_unsigned(3133, 12), 2030 => to_unsigned(1577, 12), 2031 => to_unsigned(1206, 12), 2032 => to_unsigned(2868, 12), 2033 => to_unsigned(324, 12), 2034 => to_unsigned(1835, 12), 2035 => to_unsigned(2750, 12), 2036 => to_unsigned(3111, 12), 2037 => to_unsigned(2542, 12), 2038 => to_unsigned(2912, 12), 2039 => to_unsigned(1235, 12), 2040 => to_unsigned(1113, 12), 2041 => to_unsigned(1743, 12), 2042 => to_unsigned(3724, 12), 2043 => to_unsigned(1172, 12), 2044 => to_unsigned(892, 12), 2045 => to_unsigned(3755, 12), 2046 => to_unsigned(3021, 12), 2047 => to_unsigned(1421, 12)),
            8 => (0 => to_unsigned(2865, 12), 1 => to_unsigned(2190, 12), 2 => to_unsigned(2240, 12), 3 => to_unsigned(3365, 12), 4 => to_unsigned(983, 12), 5 => to_unsigned(2597, 12), 6 => to_unsigned(1701, 12), 7 => to_unsigned(3332, 12), 8 => to_unsigned(1629, 12), 9 => to_unsigned(535, 12), 10 => to_unsigned(366, 12), 11 => to_unsigned(873, 12), 12 => to_unsigned(1297, 12), 13 => to_unsigned(686, 12), 14 => to_unsigned(3650, 12), 15 => to_unsigned(2099, 12), 16 => to_unsigned(1267, 12), 17 => to_unsigned(3595, 12), 18 => to_unsigned(2992, 12), 19 => to_unsigned(3446, 12), 20 => to_unsigned(2815, 12), 21 => to_unsigned(3391, 12), 22 => to_unsigned(132, 12), 23 => to_unsigned(2054, 12), 24 => to_unsigned(298, 12), 25 => to_unsigned(678, 12), 26 => to_unsigned(1096, 12), 27 => to_unsigned(2116, 12), 28 => to_unsigned(1580, 12), 29 => to_unsigned(3631, 12), 30 => to_unsigned(991, 12), 31 => to_unsigned(3639, 12), 32 => to_unsigned(1712, 12), 33 => to_unsigned(114, 12), 34 => to_unsigned(2878, 12), 35 => to_unsigned(3289, 12), 36 => to_unsigned(1673, 12), 37 => to_unsigned(363, 12), 38 => to_unsigned(1341, 12), 39 => to_unsigned(318, 12), 40 => to_unsigned(561, 12), 41 => to_unsigned(304, 12), 42 => to_unsigned(1892, 12), 43 => to_unsigned(3451, 12), 44 => to_unsigned(2574, 12), 45 => to_unsigned(1249, 12), 46 => to_unsigned(3595, 12), 47 => to_unsigned(401, 12), 48 => to_unsigned(1698, 12), 49 => to_unsigned(3764, 12), 50 => to_unsigned(3518, 12), 51 => to_unsigned(2018, 12), 52 => to_unsigned(3047, 12), 53 => to_unsigned(1039, 12), 54 => to_unsigned(1349, 12), 55 => to_unsigned(2718, 12), 56 => to_unsigned(728, 12), 57 => to_unsigned(930, 12), 58 => to_unsigned(959, 12), 59 => to_unsigned(1725, 12), 60 => to_unsigned(1988, 12), 61 => to_unsigned(85, 12), 62 => to_unsigned(2660, 12), 63 => to_unsigned(3062, 12), 64 => to_unsigned(929, 12), 65 => to_unsigned(2558, 12), 66 => to_unsigned(644, 12), 67 => to_unsigned(3222, 12), 68 => to_unsigned(2856, 12), 69 => to_unsigned(3859, 12), 70 => to_unsigned(928, 12), 71 => to_unsigned(3753, 12), 72 => to_unsigned(97, 12), 73 => to_unsigned(3475, 12), 74 => to_unsigned(1951, 12), 75 => to_unsigned(1131, 12), 76 => to_unsigned(1434, 12), 77 => to_unsigned(3142, 12), 78 => to_unsigned(1111, 12), 79 => to_unsigned(207, 12), 80 => to_unsigned(40, 12), 81 => to_unsigned(564, 12), 82 => to_unsigned(2117, 12), 83 => to_unsigned(1471, 12), 84 => to_unsigned(1788, 12), 85 => to_unsigned(2938, 12), 86 => to_unsigned(1421, 12), 87 => to_unsigned(3841, 12), 88 => to_unsigned(1347, 12), 89 => to_unsigned(872, 12), 90 => to_unsigned(2821, 12), 91 => to_unsigned(4004, 12), 92 => to_unsigned(1801, 12), 93 => to_unsigned(3401, 12), 94 => to_unsigned(1324, 12), 95 => to_unsigned(1676, 12), 96 => to_unsigned(933, 12), 97 => to_unsigned(933, 12), 98 => to_unsigned(2785, 12), 99 => to_unsigned(844, 12), 100 => to_unsigned(2712, 12), 101 => to_unsigned(2488, 12), 102 => to_unsigned(2404, 12), 103 => to_unsigned(2353, 12), 104 => to_unsigned(2217, 12), 105 => to_unsigned(3865, 12), 106 => to_unsigned(116, 12), 107 => to_unsigned(2204, 12), 108 => to_unsigned(725, 12), 109 => to_unsigned(2786, 12), 110 => to_unsigned(3538, 12), 111 => to_unsigned(314, 12), 112 => to_unsigned(3637, 12), 113 => to_unsigned(1939, 12), 114 => to_unsigned(1233, 12), 115 => to_unsigned(3253, 12), 116 => to_unsigned(269, 12), 117 => to_unsigned(1640, 12), 118 => to_unsigned(2449, 12), 119 => to_unsigned(2306, 12), 120 => to_unsigned(2151, 12), 121 => to_unsigned(2909, 12), 122 => to_unsigned(1723, 12), 123 => to_unsigned(3051, 12), 124 => to_unsigned(1998, 12), 125 => to_unsigned(3219, 12), 126 => to_unsigned(805, 12), 127 => to_unsigned(4034, 12), 128 => to_unsigned(1641, 12), 129 => to_unsigned(3145, 12), 130 => to_unsigned(2404, 12), 131 => to_unsigned(2066, 12), 132 => to_unsigned(3552, 12), 133 => to_unsigned(3248, 12), 134 => to_unsigned(321, 12), 135 => to_unsigned(529, 12), 136 => to_unsigned(2027, 12), 137 => to_unsigned(2873, 12), 138 => to_unsigned(3305, 12), 139 => to_unsigned(3178, 12), 140 => to_unsigned(3896, 12), 141 => to_unsigned(2677, 12), 142 => to_unsigned(2091, 12), 143 => to_unsigned(3657, 12), 144 => to_unsigned(2914, 12), 145 => to_unsigned(77, 12), 146 => to_unsigned(618, 12), 147 => to_unsigned(849, 12), 148 => to_unsigned(2479, 12), 149 => to_unsigned(687, 12), 150 => to_unsigned(46, 12), 151 => to_unsigned(2557, 12), 152 => to_unsigned(3770, 12), 153 => to_unsigned(3053, 12), 154 => to_unsigned(3765, 12), 155 => to_unsigned(12, 12), 156 => to_unsigned(957, 12), 157 => to_unsigned(4018, 12), 158 => to_unsigned(3969, 12), 159 => to_unsigned(461, 12), 160 => to_unsigned(3356, 12), 161 => to_unsigned(2314, 12), 162 => to_unsigned(3321, 12), 163 => to_unsigned(278, 12), 164 => to_unsigned(3274, 12), 165 => to_unsigned(1807, 12), 166 => to_unsigned(1090, 12), 167 => to_unsigned(1245, 12), 168 => to_unsigned(2879, 12), 169 => to_unsigned(2075, 12), 170 => to_unsigned(2240, 12), 171 => to_unsigned(2896, 12), 172 => to_unsigned(3552, 12), 173 => to_unsigned(233, 12), 174 => to_unsigned(506, 12), 175 => to_unsigned(666, 12), 176 => to_unsigned(790, 12), 177 => to_unsigned(377, 12), 178 => to_unsigned(1472, 12), 179 => to_unsigned(1974, 12), 180 => to_unsigned(609, 12), 181 => to_unsigned(3731, 12), 182 => to_unsigned(3844, 12), 183 => to_unsigned(1040, 12), 184 => to_unsigned(1760, 12), 185 => to_unsigned(2574, 12), 186 => to_unsigned(1390, 12), 187 => to_unsigned(3788, 12), 188 => to_unsigned(1429, 12), 189 => to_unsigned(2859, 12), 190 => to_unsigned(29, 12), 191 => to_unsigned(3069, 12), 192 => to_unsigned(2457, 12), 193 => to_unsigned(1871, 12), 194 => to_unsigned(3312, 12), 195 => to_unsigned(3101, 12), 196 => to_unsigned(609, 12), 197 => to_unsigned(4047, 12), 198 => to_unsigned(3232, 12), 199 => to_unsigned(3608, 12), 200 => to_unsigned(1097, 12), 201 => to_unsigned(1756, 12), 202 => to_unsigned(3220, 12), 203 => to_unsigned(666, 12), 204 => to_unsigned(3780, 12), 205 => to_unsigned(1037, 12), 206 => to_unsigned(2665, 12), 207 => to_unsigned(2836, 12), 208 => to_unsigned(1208, 12), 209 => to_unsigned(1150, 12), 210 => to_unsigned(2035, 12), 211 => to_unsigned(2096, 12), 212 => to_unsigned(3816, 12), 213 => to_unsigned(1079, 12), 214 => to_unsigned(3218, 12), 215 => to_unsigned(1383, 12), 216 => to_unsigned(1517, 12), 217 => to_unsigned(3780, 12), 218 => to_unsigned(934, 12), 219 => to_unsigned(2090, 12), 220 => to_unsigned(2647, 12), 221 => to_unsigned(398, 12), 222 => to_unsigned(22, 12), 223 => to_unsigned(1981, 12), 224 => to_unsigned(8, 12), 225 => to_unsigned(1924, 12), 226 => to_unsigned(3893, 12), 227 => to_unsigned(3671, 12), 228 => to_unsigned(2823, 12), 229 => to_unsigned(3894, 12), 230 => to_unsigned(3991, 12), 231 => to_unsigned(2121, 12), 232 => to_unsigned(714, 12), 233 => to_unsigned(2658, 12), 234 => to_unsigned(2096, 12), 235 => to_unsigned(2906, 12), 236 => to_unsigned(3637, 12), 237 => to_unsigned(2697, 12), 238 => to_unsigned(2272, 12), 239 => to_unsigned(1058, 12), 240 => to_unsigned(3056, 12), 241 => to_unsigned(3401, 12), 242 => to_unsigned(352, 12), 243 => to_unsigned(232, 12), 244 => to_unsigned(2878, 12), 245 => to_unsigned(834, 12), 246 => to_unsigned(672, 12), 247 => to_unsigned(1455, 12), 248 => to_unsigned(2085, 12), 249 => to_unsigned(3646, 12), 250 => to_unsigned(1859, 12), 251 => to_unsigned(1536, 12), 252 => to_unsigned(2846, 12), 253 => to_unsigned(3532, 12), 254 => to_unsigned(7, 12), 255 => to_unsigned(1652, 12), 256 => to_unsigned(3623, 12), 257 => to_unsigned(3590, 12), 258 => to_unsigned(709, 12), 259 => to_unsigned(2474, 12), 260 => to_unsigned(1201, 12), 261 => to_unsigned(3307, 12), 262 => to_unsigned(3895, 12), 263 => to_unsigned(2435, 12), 264 => to_unsigned(1570, 12), 265 => to_unsigned(1476, 12), 266 => to_unsigned(749, 12), 267 => to_unsigned(3697, 12), 268 => to_unsigned(1582, 12), 269 => to_unsigned(2914, 12), 270 => to_unsigned(3015, 12), 271 => to_unsigned(2348, 12), 272 => to_unsigned(2994, 12), 273 => to_unsigned(2590, 12), 274 => to_unsigned(3073, 12), 275 => to_unsigned(1573, 12), 276 => to_unsigned(1303, 12), 277 => to_unsigned(2998, 12), 278 => to_unsigned(1467, 12), 279 => to_unsigned(1164, 12), 280 => to_unsigned(3203, 12), 281 => to_unsigned(3716, 12), 282 => to_unsigned(260, 12), 283 => to_unsigned(3555, 12), 284 => to_unsigned(2835, 12), 285 => to_unsigned(3756, 12), 286 => to_unsigned(2558, 12), 287 => to_unsigned(2538, 12), 288 => to_unsigned(314, 12), 289 => to_unsigned(1607, 12), 290 => to_unsigned(65, 12), 291 => to_unsigned(4067, 12), 292 => to_unsigned(3588, 12), 293 => to_unsigned(1757, 12), 294 => to_unsigned(1587, 12), 295 => to_unsigned(51, 12), 296 => to_unsigned(258, 12), 297 => to_unsigned(307, 12), 298 => to_unsigned(1861, 12), 299 => to_unsigned(3314, 12), 300 => to_unsigned(2440, 12), 301 => to_unsigned(1526, 12), 302 => to_unsigned(2362, 12), 303 => to_unsigned(2014, 12), 304 => to_unsigned(165, 12), 305 => to_unsigned(3776, 12), 306 => to_unsigned(3751, 12), 307 => to_unsigned(239, 12), 308 => to_unsigned(1566, 12), 309 => to_unsigned(570, 12), 310 => to_unsigned(228, 12), 311 => to_unsigned(2652, 12), 312 => to_unsigned(709, 12), 313 => to_unsigned(4091, 12), 314 => to_unsigned(4033, 12), 315 => to_unsigned(428, 12), 316 => to_unsigned(3460, 12), 317 => to_unsigned(3220, 12), 318 => to_unsigned(1282, 12), 319 => to_unsigned(1281, 12), 320 => to_unsigned(2061, 12), 321 => to_unsigned(1573, 12), 322 => to_unsigned(1878, 12), 323 => to_unsigned(2731, 12), 324 => to_unsigned(2144, 12), 325 => to_unsigned(3739, 12), 326 => to_unsigned(3918, 12), 327 => to_unsigned(2698, 12), 328 => to_unsigned(3292, 12), 329 => to_unsigned(2335, 12), 330 => to_unsigned(1364, 12), 331 => to_unsigned(3455, 12), 332 => to_unsigned(1465, 12), 333 => to_unsigned(2676, 12), 334 => to_unsigned(2124, 12), 335 => to_unsigned(202, 12), 336 => to_unsigned(2032, 12), 337 => to_unsigned(919, 12), 338 => to_unsigned(645, 12), 339 => to_unsigned(1813, 12), 340 => to_unsigned(2480, 12), 341 => to_unsigned(807, 12), 342 => to_unsigned(1619, 12), 343 => to_unsigned(2970, 12), 344 => to_unsigned(619, 12), 345 => to_unsigned(244, 12), 346 => to_unsigned(496, 12), 347 => to_unsigned(3611, 12), 348 => to_unsigned(1755, 12), 349 => to_unsigned(3313, 12), 350 => to_unsigned(2103, 12), 351 => to_unsigned(397, 12), 352 => to_unsigned(3207, 12), 353 => to_unsigned(4042, 12), 354 => to_unsigned(2456, 12), 355 => to_unsigned(2767, 12), 356 => to_unsigned(2986, 12), 357 => to_unsigned(1259, 12), 358 => to_unsigned(1759, 12), 359 => to_unsigned(2869, 12), 360 => to_unsigned(527, 12), 361 => to_unsigned(1353, 12), 362 => to_unsigned(3747, 12), 363 => to_unsigned(1452, 12), 364 => to_unsigned(1315, 12), 365 => to_unsigned(1081, 12), 366 => to_unsigned(1122, 12), 367 => to_unsigned(1313, 12), 368 => to_unsigned(1937, 12), 369 => to_unsigned(1102, 12), 370 => to_unsigned(1302, 12), 371 => to_unsigned(1035, 12), 372 => to_unsigned(3482, 12), 373 => to_unsigned(2011, 12), 374 => to_unsigned(483, 12), 375 => to_unsigned(1253, 12), 376 => to_unsigned(2799, 12), 377 => to_unsigned(821, 12), 378 => to_unsigned(558, 12), 379 => to_unsigned(683, 12), 380 => to_unsigned(1564, 12), 381 => to_unsigned(2298, 12), 382 => to_unsigned(2687, 12), 383 => to_unsigned(3301, 12), 384 => to_unsigned(368, 12), 385 => to_unsigned(2078, 12), 386 => to_unsigned(1711, 12), 387 => to_unsigned(2303, 12), 388 => to_unsigned(2885, 12), 389 => to_unsigned(41, 12), 390 => to_unsigned(1386, 12), 391 => to_unsigned(518, 12), 392 => to_unsigned(1828, 12), 393 => to_unsigned(587, 12), 394 => to_unsigned(3045, 12), 395 => to_unsigned(2609, 12), 396 => to_unsigned(2131, 12), 397 => to_unsigned(1376, 12), 398 => to_unsigned(2170, 12), 399 => to_unsigned(1420, 12), 400 => to_unsigned(3525, 12), 401 => to_unsigned(415, 12), 402 => to_unsigned(377, 12), 403 => to_unsigned(1818, 12), 404 => to_unsigned(4033, 12), 405 => to_unsigned(2861, 12), 406 => to_unsigned(2587, 12), 407 => to_unsigned(3456, 12), 408 => to_unsigned(632, 12), 409 => to_unsigned(2460, 12), 410 => to_unsigned(2715, 12), 411 => to_unsigned(308, 12), 412 => to_unsigned(565, 12), 413 => to_unsigned(2535, 12), 414 => to_unsigned(2811, 12), 415 => to_unsigned(2243, 12), 416 => to_unsigned(2983, 12), 417 => to_unsigned(2697, 12), 418 => to_unsigned(234, 12), 419 => to_unsigned(3048, 12), 420 => to_unsigned(252, 12), 421 => to_unsigned(2741, 12), 422 => to_unsigned(1045, 12), 423 => to_unsigned(2191, 12), 424 => to_unsigned(3509, 12), 425 => to_unsigned(2668, 12), 426 => to_unsigned(2525, 12), 427 => to_unsigned(3902, 12), 428 => to_unsigned(205, 12), 429 => to_unsigned(1701, 12), 430 => to_unsigned(90, 12), 431 => to_unsigned(1904, 12), 432 => to_unsigned(520, 12), 433 => to_unsigned(3348, 12), 434 => to_unsigned(1591, 12), 435 => to_unsigned(3563, 12), 436 => to_unsigned(2931, 12), 437 => to_unsigned(2437, 12), 438 => to_unsigned(3136, 12), 439 => to_unsigned(184, 12), 440 => to_unsigned(2760, 12), 441 => to_unsigned(2923, 12), 442 => to_unsigned(1646, 12), 443 => to_unsigned(2466, 12), 444 => to_unsigned(2282, 12), 445 => to_unsigned(2787, 12), 446 => to_unsigned(952, 12), 447 => to_unsigned(793, 12), 448 => to_unsigned(3424, 12), 449 => to_unsigned(1971, 12), 450 => to_unsigned(1366, 12), 451 => to_unsigned(99, 12), 452 => to_unsigned(4025, 12), 453 => to_unsigned(1773, 12), 454 => to_unsigned(442, 12), 455 => to_unsigned(2502, 12), 456 => to_unsigned(2977, 12), 457 => to_unsigned(3574, 12), 458 => to_unsigned(3966, 12), 459 => to_unsigned(2640, 12), 460 => to_unsigned(2077, 12), 461 => to_unsigned(2318, 12), 462 => to_unsigned(1623, 12), 463 => to_unsigned(456, 12), 464 => to_unsigned(1151, 12), 465 => to_unsigned(2950, 12), 466 => to_unsigned(3391, 12), 467 => to_unsigned(72, 12), 468 => to_unsigned(1516, 12), 469 => to_unsigned(3513, 12), 470 => to_unsigned(1048, 12), 471 => to_unsigned(2247, 12), 472 => to_unsigned(2899, 12), 473 => to_unsigned(2442, 12), 474 => to_unsigned(861, 12), 475 => to_unsigned(1712, 12), 476 => to_unsigned(2883, 12), 477 => to_unsigned(1173, 12), 478 => to_unsigned(636, 12), 479 => to_unsigned(237, 12), 480 => to_unsigned(2580, 12), 481 => to_unsigned(3575, 12), 482 => to_unsigned(1483, 12), 483 => to_unsigned(1559, 12), 484 => to_unsigned(883, 12), 485 => to_unsigned(1124, 12), 486 => to_unsigned(2352, 12), 487 => to_unsigned(1924, 12), 488 => to_unsigned(3672, 12), 489 => to_unsigned(1931, 12), 490 => to_unsigned(2415, 12), 491 => to_unsigned(3018, 12), 492 => to_unsigned(1204, 12), 493 => to_unsigned(3871, 12), 494 => to_unsigned(2862, 12), 495 => to_unsigned(2390, 12), 496 => to_unsigned(2902, 12), 497 => to_unsigned(2721, 12), 498 => to_unsigned(1486, 12), 499 => to_unsigned(651, 12), 500 => to_unsigned(1117, 12), 501 => to_unsigned(3540, 12), 502 => to_unsigned(1476, 12), 503 => to_unsigned(1654, 12), 504 => to_unsigned(3126, 12), 505 => to_unsigned(4072, 12), 506 => to_unsigned(1476, 12), 507 => to_unsigned(2755, 12), 508 => to_unsigned(437, 12), 509 => to_unsigned(4003, 12), 510 => to_unsigned(2459, 12), 511 => to_unsigned(1243, 12), 512 => to_unsigned(3475, 12), 513 => to_unsigned(3212, 12), 514 => to_unsigned(74, 12), 515 => to_unsigned(1050, 12), 516 => to_unsigned(612, 12), 517 => to_unsigned(2919, 12), 518 => to_unsigned(1896, 12), 519 => to_unsigned(1222, 12), 520 => to_unsigned(2453, 12), 521 => to_unsigned(2023, 12), 522 => to_unsigned(623, 12), 523 => to_unsigned(29, 12), 524 => to_unsigned(806, 12), 525 => to_unsigned(1145, 12), 526 => to_unsigned(1460, 12), 527 => to_unsigned(625, 12), 528 => to_unsigned(2190, 12), 529 => to_unsigned(331, 12), 530 => to_unsigned(451, 12), 531 => to_unsigned(3390, 12), 532 => to_unsigned(2176, 12), 533 => to_unsigned(2086, 12), 534 => to_unsigned(3039, 12), 535 => to_unsigned(2090, 12), 536 => to_unsigned(2690, 12), 537 => to_unsigned(3876, 12), 538 => to_unsigned(3182, 12), 539 => to_unsigned(385, 12), 540 => to_unsigned(2894, 12), 541 => to_unsigned(713, 12), 542 => to_unsigned(3121, 12), 543 => to_unsigned(2136, 12), 544 => to_unsigned(2365, 12), 545 => to_unsigned(864, 12), 546 => to_unsigned(2060, 12), 547 => to_unsigned(3475, 12), 548 => to_unsigned(2800, 12), 549 => to_unsigned(1222, 12), 550 => to_unsigned(3606, 12), 551 => to_unsigned(3147, 12), 552 => to_unsigned(1706, 12), 553 => to_unsigned(3025, 12), 554 => to_unsigned(2502, 12), 555 => to_unsigned(2536, 12), 556 => to_unsigned(1482, 12), 557 => to_unsigned(1538, 12), 558 => to_unsigned(2128, 12), 559 => to_unsigned(3423, 12), 560 => to_unsigned(263, 12), 561 => to_unsigned(4045, 12), 562 => to_unsigned(3861, 12), 563 => to_unsigned(2651, 12), 564 => to_unsigned(49, 12), 565 => to_unsigned(1357, 12), 566 => to_unsigned(2185, 12), 567 => to_unsigned(4027, 12), 568 => to_unsigned(2473, 12), 569 => to_unsigned(1406, 12), 570 => to_unsigned(222, 12), 571 => to_unsigned(1609, 12), 572 => to_unsigned(62, 12), 573 => to_unsigned(1835, 12), 574 => to_unsigned(803, 12), 575 => to_unsigned(118, 12), 576 => to_unsigned(373, 12), 577 => to_unsigned(1034, 12), 578 => to_unsigned(3701, 12), 579 => to_unsigned(1320, 12), 580 => to_unsigned(2121, 12), 581 => to_unsigned(58, 12), 582 => to_unsigned(3043, 12), 583 => to_unsigned(3824, 12), 584 => to_unsigned(484, 12), 585 => to_unsigned(2328, 12), 586 => to_unsigned(2860, 12), 587 => to_unsigned(2863, 12), 588 => to_unsigned(2886, 12), 589 => to_unsigned(2087, 12), 590 => to_unsigned(3459, 12), 591 => to_unsigned(2026, 12), 592 => to_unsigned(2294, 12), 593 => to_unsigned(2435, 12), 594 => to_unsigned(9, 12), 595 => to_unsigned(2082, 12), 596 => to_unsigned(1639, 12), 597 => to_unsigned(2221, 12), 598 => to_unsigned(1069, 12), 599 => to_unsigned(2785, 12), 600 => to_unsigned(2084, 12), 601 => to_unsigned(818, 12), 602 => to_unsigned(2192, 12), 603 => to_unsigned(633, 12), 604 => to_unsigned(2854, 12), 605 => to_unsigned(555, 12), 606 => to_unsigned(3689, 12), 607 => to_unsigned(742, 12), 608 => to_unsigned(1127, 12), 609 => to_unsigned(1312, 12), 610 => to_unsigned(3317, 12), 611 => to_unsigned(1321, 12), 612 => to_unsigned(418, 12), 613 => to_unsigned(2092, 12), 614 => to_unsigned(491, 12), 615 => to_unsigned(1304, 12), 616 => to_unsigned(942, 12), 617 => to_unsigned(1686, 12), 618 => to_unsigned(3786, 12), 619 => to_unsigned(2192, 12), 620 => to_unsigned(97, 12), 621 => to_unsigned(630, 12), 622 => to_unsigned(1196, 12), 623 => to_unsigned(302, 12), 624 => to_unsigned(1269, 12), 625 => to_unsigned(2777, 12), 626 => to_unsigned(3072, 12), 627 => to_unsigned(885, 12), 628 => to_unsigned(480, 12), 629 => to_unsigned(2932, 12), 630 => to_unsigned(2906, 12), 631 => to_unsigned(63, 12), 632 => to_unsigned(3292, 12), 633 => to_unsigned(1974, 12), 634 => to_unsigned(3861, 12), 635 => to_unsigned(4000, 12), 636 => to_unsigned(1583, 12), 637 => to_unsigned(1776, 12), 638 => to_unsigned(2019, 12), 639 => to_unsigned(1774, 12), 640 => to_unsigned(2676, 12), 641 => to_unsigned(659, 12), 642 => to_unsigned(2168, 12), 643 => to_unsigned(4035, 12), 644 => to_unsigned(3344, 12), 645 => to_unsigned(1378, 12), 646 => to_unsigned(497, 12), 647 => to_unsigned(3458, 12), 648 => to_unsigned(1329, 12), 649 => to_unsigned(1706, 12), 650 => to_unsigned(3022, 12), 651 => to_unsigned(3960, 12), 652 => to_unsigned(1251, 12), 653 => to_unsigned(1200, 12), 654 => to_unsigned(643, 12), 655 => to_unsigned(1642, 12), 656 => to_unsigned(2171, 12), 657 => to_unsigned(1853, 12), 658 => to_unsigned(2577, 12), 659 => to_unsigned(2839, 12), 660 => to_unsigned(2022, 12), 661 => to_unsigned(1679, 12), 662 => to_unsigned(1822, 12), 663 => to_unsigned(2917, 12), 664 => to_unsigned(3963, 12), 665 => to_unsigned(3237, 12), 666 => to_unsigned(2163, 12), 667 => to_unsigned(1449, 12), 668 => to_unsigned(3272, 12), 669 => to_unsigned(2027, 12), 670 => to_unsigned(2003, 12), 671 => to_unsigned(221, 12), 672 => to_unsigned(3405, 12), 673 => to_unsigned(1468, 12), 674 => to_unsigned(3032, 12), 675 => to_unsigned(2869, 12), 676 => to_unsigned(2077, 12), 677 => to_unsigned(2430, 12), 678 => to_unsigned(3402, 12), 679 => to_unsigned(3543, 12), 680 => to_unsigned(3528, 12), 681 => to_unsigned(3335, 12), 682 => to_unsigned(2695, 12), 683 => to_unsigned(976, 12), 684 => to_unsigned(924, 12), 685 => to_unsigned(3681, 12), 686 => to_unsigned(1041, 12), 687 => to_unsigned(1816, 12), 688 => to_unsigned(3136, 12), 689 => to_unsigned(930, 12), 690 => to_unsigned(1183, 12), 691 => to_unsigned(1212, 12), 692 => to_unsigned(1759, 12), 693 => to_unsigned(2634, 12), 694 => to_unsigned(2903, 12), 695 => to_unsigned(1653, 12), 696 => to_unsigned(1836, 12), 697 => to_unsigned(535, 12), 698 => to_unsigned(1609, 12), 699 => to_unsigned(2637, 12), 700 => to_unsigned(1648, 12), 701 => to_unsigned(2309, 12), 702 => to_unsigned(3369, 12), 703 => to_unsigned(2830, 12), 704 => to_unsigned(1418, 12), 705 => to_unsigned(692, 12), 706 => to_unsigned(925, 12), 707 => to_unsigned(3702, 12), 708 => to_unsigned(3035, 12), 709 => to_unsigned(3620, 12), 710 => to_unsigned(1551, 12), 711 => to_unsigned(4049, 12), 712 => to_unsigned(3065, 12), 713 => to_unsigned(3112, 12), 714 => to_unsigned(156, 12), 715 => to_unsigned(3, 12), 716 => to_unsigned(2335, 12), 717 => to_unsigned(54, 12), 718 => to_unsigned(1778, 12), 719 => to_unsigned(614, 12), 720 => to_unsigned(1827, 12), 721 => to_unsigned(2217, 12), 722 => to_unsigned(1322, 12), 723 => to_unsigned(1581, 12), 724 => to_unsigned(3346, 12), 725 => to_unsigned(833, 12), 726 => to_unsigned(114, 12), 727 => to_unsigned(2669, 12), 728 => to_unsigned(3581, 12), 729 => to_unsigned(4067, 12), 730 => to_unsigned(241, 12), 731 => to_unsigned(3369, 12), 732 => to_unsigned(1399, 12), 733 => to_unsigned(114, 12), 734 => to_unsigned(2951, 12), 735 => to_unsigned(2322, 12), 736 => to_unsigned(3428, 12), 737 => to_unsigned(4062, 12), 738 => to_unsigned(856, 12), 739 => to_unsigned(3101, 12), 740 => to_unsigned(1188, 12), 741 => to_unsigned(1334, 12), 742 => to_unsigned(1580, 12), 743 => to_unsigned(3249, 12), 744 => to_unsigned(1600, 12), 745 => to_unsigned(2262, 12), 746 => to_unsigned(2894, 12), 747 => to_unsigned(2262, 12), 748 => to_unsigned(3984, 12), 749 => to_unsigned(3576, 12), 750 => to_unsigned(1050, 12), 751 => to_unsigned(2086, 12), 752 => to_unsigned(1195, 12), 753 => to_unsigned(2852, 12), 754 => to_unsigned(3275, 12), 755 => to_unsigned(2102, 12), 756 => to_unsigned(2536, 12), 757 => to_unsigned(2947, 12), 758 => to_unsigned(3772, 12), 759 => to_unsigned(3348, 12), 760 => to_unsigned(2233, 12), 761 => to_unsigned(506, 12), 762 => to_unsigned(1547, 12), 763 => to_unsigned(2989, 12), 764 => to_unsigned(705, 12), 765 => to_unsigned(3942, 12), 766 => to_unsigned(2394, 12), 767 => to_unsigned(145, 12), 768 => to_unsigned(2052, 12), 769 => to_unsigned(1652, 12), 770 => to_unsigned(2468, 12), 771 => to_unsigned(951, 12), 772 => to_unsigned(2180, 12), 773 => to_unsigned(534, 12), 774 => to_unsigned(2116, 12), 775 => to_unsigned(592, 12), 776 => to_unsigned(72, 12), 777 => to_unsigned(2807, 12), 778 => to_unsigned(256, 12), 779 => to_unsigned(3591, 12), 780 => to_unsigned(3727, 12), 781 => to_unsigned(384, 12), 782 => to_unsigned(3750, 12), 783 => to_unsigned(660, 12), 784 => to_unsigned(3045, 12), 785 => to_unsigned(1819, 12), 786 => to_unsigned(3573, 12), 787 => to_unsigned(1813, 12), 788 => to_unsigned(3918, 12), 789 => to_unsigned(312, 12), 790 => to_unsigned(2916, 12), 791 => to_unsigned(1292, 12), 792 => to_unsigned(3335, 12), 793 => to_unsigned(3823, 12), 794 => to_unsigned(3830, 12), 795 => to_unsigned(1900, 12), 796 => to_unsigned(3364, 12), 797 => to_unsigned(2903, 12), 798 => to_unsigned(1915, 12), 799 => to_unsigned(1443, 12), 800 => to_unsigned(341, 12), 801 => to_unsigned(1819, 12), 802 => to_unsigned(1271, 12), 803 => to_unsigned(1234, 12), 804 => to_unsigned(75, 12), 805 => to_unsigned(1277, 12), 806 => to_unsigned(3154, 12), 807 => to_unsigned(1070, 12), 808 => to_unsigned(2268, 12), 809 => to_unsigned(507, 12), 810 => to_unsigned(452, 12), 811 => to_unsigned(1437, 12), 812 => to_unsigned(1948, 12), 813 => to_unsigned(3331, 12), 814 => to_unsigned(872, 12), 815 => to_unsigned(256, 12), 816 => to_unsigned(1160, 12), 817 => to_unsigned(1292, 12), 818 => to_unsigned(1428, 12), 819 => to_unsigned(2676, 12), 820 => to_unsigned(234, 12), 821 => to_unsigned(2815, 12), 822 => to_unsigned(2386, 12), 823 => to_unsigned(2645, 12), 824 => to_unsigned(2126, 12), 825 => to_unsigned(545, 12), 826 => to_unsigned(2679, 12), 827 => to_unsigned(280, 12), 828 => to_unsigned(733, 12), 829 => to_unsigned(3209, 12), 830 => to_unsigned(2217, 12), 831 => to_unsigned(2579, 12), 832 => to_unsigned(3444, 12), 833 => to_unsigned(3031, 12), 834 => to_unsigned(234, 12), 835 => to_unsigned(3279, 12), 836 => to_unsigned(851, 12), 837 => to_unsigned(1360, 12), 838 => to_unsigned(577, 12), 839 => to_unsigned(3773, 12), 840 => to_unsigned(2263, 12), 841 => to_unsigned(123, 12), 842 => to_unsigned(2461, 12), 843 => to_unsigned(1583, 12), 844 => to_unsigned(3075, 12), 845 => to_unsigned(2290, 12), 846 => to_unsigned(3564, 12), 847 => to_unsigned(462, 12), 848 => to_unsigned(662, 12), 849 => to_unsigned(567, 12), 850 => to_unsigned(1717, 12), 851 => to_unsigned(475, 12), 852 => to_unsigned(562, 12), 853 => to_unsigned(3563, 12), 854 => to_unsigned(1688, 12), 855 => to_unsigned(2396, 12), 856 => to_unsigned(979, 12), 857 => to_unsigned(3295, 12), 858 => to_unsigned(1561, 12), 859 => to_unsigned(1210, 12), 860 => to_unsigned(2930, 12), 861 => to_unsigned(2434, 12), 862 => to_unsigned(2461, 12), 863 => to_unsigned(817, 12), 864 => to_unsigned(2611, 12), 865 => to_unsigned(1749, 12), 866 => to_unsigned(3380, 12), 867 => to_unsigned(2068, 12), 868 => to_unsigned(1043, 12), 869 => to_unsigned(3042, 12), 870 => to_unsigned(2902, 12), 871 => to_unsigned(2951, 12), 872 => to_unsigned(2612, 12), 873 => to_unsigned(2265, 12), 874 => to_unsigned(10, 12), 875 => to_unsigned(1716, 12), 876 => to_unsigned(432, 12), 877 => to_unsigned(370, 12), 878 => to_unsigned(999, 12), 879 => to_unsigned(2174, 12), 880 => to_unsigned(854, 12), 881 => to_unsigned(1554, 12), 882 => to_unsigned(151, 12), 883 => to_unsigned(850, 12), 884 => to_unsigned(3542, 12), 885 => to_unsigned(2932, 12), 886 => to_unsigned(868, 12), 887 => to_unsigned(2484, 12), 888 => to_unsigned(2683, 12), 889 => to_unsigned(2919, 12), 890 => to_unsigned(2304, 12), 891 => to_unsigned(828, 12), 892 => to_unsigned(3292, 12), 893 => to_unsigned(2308, 12), 894 => to_unsigned(1914, 12), 895 => to_unsigned(810, 12), 896 => to_unsigned(3154, 12), 897 => to_unsigned(70, 12), 898 => to_unsigned(1916, 12), 899 => to_unsigned(4001, 12), 900 => to_unsigned(614, 12), 901 => to_unsigned(2084, 12), 902 => to_unsigned(3421, 12), 903 => to_unsigned(1782, 12), 904 => to_unsigned(3884, 12), 905 => to_unsigned(3954, 12), 906 => to_unsigned(1383, 12), 907 => to_unsigned(1080, 12), 908 => to_unsigned(2944, 12), 909 => to_unsigned(3064, 12), 910 => to_unsigned(688, 12), 911 => to_unsigned(2925, 12), 912 => to_unsigned(536, 12), 913 => to_unsigned(3865, 12), 914 => to_unsigned(3889, 12), 915 => to_unsigned(2965, 12), 916 => to_unsigned(3388, 12), 917 => to_unsigned(129, 12), 918 => to_unsigned(2656, 12), 919 => to_unsigned(62, 12), 920 => to_unsigned(828, 12), 921 => to_unsigned(1928, 12), 922 => to_unsigned(633, 12), 923 => to_unsigned(3325, 12), 924 => to_unsigned(2056, 12), 925 => to_unsigned(699, 12), 926 => to_unsigned(887, 12), 927 => to_unsigned(2336, 12), 928 => to_unsigned(1247, 12), 929 => to_unsigned(1080, 12), 930 => to_unsigned(3927, 12), 931 => to_unsigned(279, 12), 932 => to_unsigned(441, 12), 933 => to_unsigned(2447, 12), 934 => to_unsigned(3583, 12), 935 => to_unsigned(1190, 12), 936 => to_unsigned(2597, 12), 937 => to_unsigned(2358, 12), 938 => to_unsigned(480, 12), 939 => to_unsigned(3894, 12), 940 => to_unsigned(1120, 12), 941 => to_unsigned(2729, 12), 942 => to_unsigned(1134, 12), 943 => to_unsigned(3357, 12), 944 => to_unsigned(380, 12), 945 => to_unsigned(3629, 12), 946 => to_unsigned(255, 12), 947 => to_unsigned(2945, 12), 948 => to_unsigned(1695, 12), 949 => to_unsigned(3710, 12), 950 => to_unsigned(798, 12), 951 => to_unsigned(217, 12), 952 => to_unsigned(1571, 12), 953 => to_unsigned(786, 12), 954 => to_unsigned(1055, 12), 955 => to_unsigned(1732, 12), 956 => to_unsigned(6, 12), 957 => to_unsigned(3017, 12), 958 => to_unsigned(3186, 12), 959 => to_unsigned(3783, 12), 960 => to_unsigned(2181, 12), 961 => to_unsigned(4011, 12), 962 => to_unsigned(3774, 12), 963 => to_unsigned(1657, 12), 964 => to_unsigned(2402, 12), 965 => to_unsigned(1755, 12), 966 => to_unsigned(969, 12), 967 => to_unsigned(3811, 12), 968 => to_unsigned(176, 12), 969 => to_unsigned(238, 12), 970 => to_unsigned(598, 12), 971 => to_unsigned(356, 12), 972 => to_unsigned(1399, 12), 973 => to_unsigned(1539, 12), 974 => to_unsigned(467, 12), 975 => to_unsigned(2235, 12), 976 => to_unsigned(3348, 12), 977 => to_unsigned(3984, 12), 978 => to_unsigned(2341, 12), 979 => to_unsigned(1709, 12), 980 => to_unsigned(2307, 12), 981 => to_unsigned(895, 12), 982 => to_unsigned(536, 12), 983 => to_unsigned(1900, 12), 984 => to_unsigned(1599, 12), 985 => to_unsigned(1312, 12), 986 => to_unsigned(1096, 12), 987 => to_unsigned(3925, 12), 988 => to_unsigned(792, 12), 989 => to_unsigned(1988, 12), 990 => to_unsigned(3079, 12), 991 => to_unsigned(1948, 12), 992 => to_unsigned(359, 12), 993 => to_unsigned(1073, 12), 994 => to_unsigned(2526, 12), 995 => to_unsigned(610, 12), 996 => to_unsigned(3302, 12), 997 => to_unsigned(1636, 12), 998 => to_unsigned(3520, 12), 999 => to_unsigned(1859, 12), 1000 => to_unsigned(2142, 12), 1001 => to_unsigned(613, 12), 1002 => to_unsigned(1715, 12), 1003 => to_unsigned(2866, 12), 1004 => to_unsigned(2236, 12), 1005 => to_unsigned(970, 12), 1006 => to_unsigned(2618, 12), 1007 => to_unsigned(2512, 12), 1008 => to_unsigned(3924, 12), 1009 => to_unsigned(652, 12), 1010 => to_unsigned(2046, 12), 1011 => to_unsigned(1672, 12), 1012 => to_unsigned(579, 12), 1013 => to_unsigned(3683, 12), 1014 => to_unsigned(635, 12), 1015 => to_unsigned(1525, 12), 1016 => to_unsigned(1449, 12), 1017 => to_unsigned(348, 12), 1018 => to_unsigned(1825, 12), 1019 => to_unsigned(3336, 12), 1020 => to_unsigned(1251, 12), 1021 => to_unsigned(3116, 12), 1022 => to_unsigned(2320, 12), 1023 => to_unsigned(3976, 12), 1024 => to_unsigned(2061, 12), 1025 => to_unsigned(820, 12), 1026 => to_unsigned(1674, 12), 1027 => to_unsigned(3186, 12), 1028 => to_unsigned(374, 12), 1029 => to_unsigned(1520, 12), 1030 => to_unsigned(1216, 12), 1031 => to_unsigned(1722, 12), 1032 => to_unsigned(3088, 12), 1033 => to_unsigned(2727, 12), 1034 => to_unsigned(972, 12), 1035 => to_unsigned(2077, 12), 1036 => to_unsigned(20, 12), 1037 => to_unsigned(3700, 12), 1038 => to_unsigned(1440, 12), 1039 => to_unsigned(2683, 12), 1040 => to_unsigned(3159, 12), 1041 => to_unsigned(2570, 12), 1042 => to_unsigned(1042, 12), 1043 => to_unsigned(3467, 12), 1044 => to_unsigned(1066, 12), 1045 => to_unsigned(3339, 12), 1046 => to_unsigned(1479, 12), 1047 => to_unsigned(4038, 12), 1048 => to_unsigned(2455, 12), 1049 => to_unsigned(1911, 12), 1050 => to_unsigned(1216, 12), 1051 => to_unsigned(1632, 12), 1052 => to_unsigned(3464, 12), 1053 => to_unsigned(54, 12), 1054 => to_unsigned(387, 12), 1055 => to_unsigned(646, 12), 1056 => to_unsigned(3694, 12), 1057 => to_unsigned(1170, 12), 1058 => to_unsigned(3524, 12), 1059 => to_unsigned(3408, 12), 1060 => to_unsigned(2524, 12), 1061 => to_unsigned(2867, 12), 1062 => to_unsigned(3144, 12), 1063 => to_unsigned(2906, 12), 1064 => to_unsigned(2227, 12), 1065 => to_unsigned(2675, 12), 1066 => to_unsigned(3204, 12), 1067 => to_unsigned(3181, 12), 1068 => to_unsigned(243, 12), 1069 => to_unsigned(3227, 12), 1070 => to_unsigned(1792, 12), 1071 => to_unsigned(1820, 12), 1072 => to_unsigned(606, 12), 1073 => to_unsigned(3870, 12), 1074 => to_unsigned(3117, 12), 1075 => to_unsigned(584, 12), 1076 => to_unsigned(60, 12), 1077 => to_unsigned(3729, 12), 1078 => to_unsigned(1234, 12), 1079 => to_unsigned(2098, 12), 1080 => to_unsigned(1274, 12), 1081 => to_unsigned(3166, 12), 1082 => to_unsigned(1998, 12), 1083 => to_unsigned(559, 12), 1084 => to_unsigned(3606, 12), 1085 => to_unsigned(143, 12), 1086 => to_unsigned(4055, 12), 1087 => to_unsigned(894, 12), 1088 => to_unsigned(2587, 12), 1089 => to_unsigned(1825, 12), 1090 => to_unsigned(245, 12), 1091 => to_unsigned(2750, 12), 1092 => to_unsigned(3013, 12), 1093 => to_unsigned(3544, 12), 1094 => to_unsigned(956, 12), 1095 => to_unsigned(3407, 12), 1096 => to_unsigned(3387, 12), 1097 => to_unsigned(375, 12), 1098 => to_unsigned(130, 12), 1099 => to_unsigned(1674, 12), 1100 => to_unsigned(3214, 12), 1101 => to_unsigned(1152, 12), 1102 => to_unsigned(3559, 12), 1103 => to_unsigned(423, 12), 1104 => to_unsigned(2063, 12), 1105 => to_unsigned(850, 12), 1106 => to_unsigned(1264, 12), 1107 => to_unsigned(799, 12), 1108 => to_unsigned(1737, 12), 1109 => to_unsigned(1001, 12), 1110 => to_unsigned(3449, 12), 1111 => to_unsigned(2858, 12), 1112 => to_unsigned(3535, 12), 1113 => to_unsigned(633, 12), 1114 => to_unsigned(1127, 12), 1115 => to_unsigned(2936, 12), 1116 => to_unsigned(1636, 12), 1117 => to_unsigned(835, 12), 1118 => to_unsigned(2971, 12), 1119 => to_unsigned(944, 12), 1120 => to_unsigned(789, 12), 1121 => to_unsigned(164, 12), 1122 => to_unsigned(916, 12), 1123 => to_unsigned(871, 12), 1124 => to_unsigned(4063, 12), 1125 => to_unsigned(3057, 12), 1126 => to_unsigned(395, 12), 1127 => to_unsigned(2042, 12), 1128 => to_unsigned(664, 12), 1129 => to_unsigned(2001, 12), 1130 => to_unsigned(3404, 12), 1131 => to_unsigned(3010, 12), 1132 => to_unsigned(1658, 12), 1133 => to_unsigned(193, 12), 1134 => to_unsigned(2554, 12), 1135 => to_unsigned(2961, 12), 1136 => to_unsigned(1649, 12), 1137 => to_unsigned(3660, 12), 1138 => to_unsigned(2469, 12), 1139 => to_unsigned(1460, 12), 1140 => to_unsigned(1715, 12), 1141 => to_unsigned(1070, 12), 1142 => to_unsigned(3564, 12), 1143 => to_unsigned(3173, 12), 1144 => to_unsigned(2603, 12), 1145 => to_unsigned(2820, 12), 1146 => to_unsigned(1443, 12), 1147 => to_unsigned(175, 12), 1148 => to_unsigned(702, 12), 1149 => to_unsigned(2582, 12), 1150 => to_unsigned(3935, 12), 1151 => to_unsigned(2432, 12), 1152 => to_unsigned(3506, 12), 1153 => to_unsigned(3528, 12), 1154 => to_unsigned(1820, 12), 1155 => to_unsigned(1336, 12), 1156 => to_unsigned(2033, 12), 1157 => to_unsigned(2283, 12), 1158 => to_unsigned(1527, 12), 1159 => to_unsigned(3770, 12), 1160 => to_unsigned(3853, 12), 1161 => to_unsigned(946, 12), 1162 => to_unsigned(3436, 12), 1163 => to_unsigned(1859, 12), 1164 => to_unsigned(3704, 12), 1165 => to_unsigned(501, 12), 1166 => to_unsigned(1831, 12), 1167 => to_unsigned(2404, 12), 1168 => to_unsigned(697, 12), 1169 => to_unsigned(2230, 12), 1170 => to_unsigned(263, 12), 1171 => to_unsigned(3715, 12), 1172 => to_unsigned(3638, 12), 1173 => to_unsigned(2731, 12), 1174 => to_unsigned(2024, 12), 1175 => to_unsigned(2118, 12), 1176 => to_unsigned(1472, 12), 1177 => to_unsigned(3734, 12), 1178 => to_unsigned(3169, 12), 1179 => to_unsigned(3294, 12), 1180 => to_unsigned(968, 12), 1181 => to_unsigned(462, 12), 1182 => to_unsigned(3280, 12), 1183 => to_unsigned(3022, 12), 1184 => to_unsigned(3378, 12), 1185 => to_unsigned(897, 12), 1186 => to_unsigned(3646, 12), 1187 => to_unsigned(387, 12), 1188 => to_unsigned(919, 12), 1189 => to_unsigned(3098, 12), 1190 => to_unsigned(817, 12), 1191 => to_unsigned(1815, 12), 1192 => to_unsigned(650, 12), 1193 => to_unsigned(783, 12), 1194 => to_unsigned(1985, 12), 1195 => to_unsigned(1532, 12), 1196 => to_unsigned(212, 12), 1197 => to_unsigned(1239, 12), 1198 => to_unsigned(3606, 12), 1199 => to_unsigned(1003, 12), 1200 => to_unsigned(1012, 12), 1201 => to_unsigned(142, 12), 1202 => to_unsigned(1425, 12), 1203 => to_unsigned(4014, 12), 1204 => to_unsigned(3567, 12), 1205 => to_unsigned(3661, 12), 1206 => to_unsigned(944, 12), 1207 => to_unsigned(3773, 12), 1208 => to_unsigned(465, 12), 1209 => to_unsigned(3505, 12), 1210 => to_unsigned(1437, 12), 1211 => to_unsigned(124, 12), 1212 => to_unsigned(1347, 12), 1213 => to_unsigned(140, 12), 1214 => to_unsigned(3992, 12), 1215 => to_unsigned(3608, 12), 1216 => to_unsigned(702, 12), 1217 => to_unsigned(2981, 12), 1218 => to_unsigned(1611, 12), 1219 => to_unsigned(3429, 12), 1220 => to_unsigned(2058, 12), 1221 => to_unsigned(2246, 12), 1222 => to_unsigned(428, 12), 1223 => to_unsigned(3970, 12), 1224 => to_unsigned(1435, 12), 1225 => to_unsigned(1593, 12), 1226 => to_unsigned(726, 12), 1227 => to_unsigned(3197, 12), 1228 => to_unsigned(4081, 12), 1229 => to_unsigned(1100, 12), 1230 => to_unsigned(1151, 12), 1231 => to_unsigned(1797, 12), 1232 => to_unsigned(2703, 12), 1233 => to_unsigned(2454, 12), 1234 => to_unsigned(2109, 12), 1235 => to_unsigned(1585, 12), 1236 => to_unsigned(690, 12), 1237 => to_unsigned(1184, 12), 1238 => to_unsigned(1362, 12), 1239 => to_unsigned(1359, 12), 1240 => to_unsigned(2226, 12), 1241 => to_unsigned(152, 12), 1242 => to_unsigned(57, 12), 1243 => to_unsigned(2946, 12), 1244 => to_unsigned(3220, 12), 1245 => to_unsigned(3985, 12), 1246 => to_unsigned(3813, 12), 1247 => to_unsigned(2364, 12), 1248 => to_unsigned(2518, 12), 1249 => to_unsigned(3293, 12), 1250 => to_unsigned(1524, 12), 1251 => to_unsigned(1159, 12), 1252 => to_unsigned(1688, 12), 1253 => to_unsigned(3600, 12), 1254 => to_unsigned(707, 12), 1255 => to_unsigned(445, 12), 1256 => to_unsigned(3309, 12), 1257 => to_unsigned(1925, 12), 1258 => to_unsigned(497, 12), 1259 => to_unsigned(672, 12), 1260 => to_unsigned(2736, 12), 1261 => to_unsigned(2030, 12), 1262 => to_unsigned(3212, 12), 1263 => to_unsigned(1793, 12), 1264 => to_unsigned(1989, 12), 1265 => to_unsigned(3243, 12), 1266 => to_unsigned(2962, 12), 1267 => to_unsigned(2889, 12), 1268 => to_unsigned(2850, 12), 1269 => to_unsigned(1720, 12), 1270 => to_unsigned(240, 12), 1271 => to_unsigned(1770, 12), 1272 => to_unsigned(125, 12), 1273 => to_unsigned(3688, 12), 1274 => to_unsigned(3571, 12), 1275 => to_unsigned(1237, 12), 1276 => to_unsigned(1580, 12), 1277 => to_unsigned(3961, 12), 1278 => to_unsigned(1984, 12), 1279 => to_unsigned(3833, 12), 1280 => to_unsigned(2744, 12), 1281 => to_unsigned(970, 12), 1282 => to_unsigned(3764, 12), 1283 => to_unsigned(2169, 12), 1284 => to_unsigned(3082, 12), 1285 => to_unsigned(3164, 12), 1286 => to_unsigned(3092, 12), 1287 => to_unsigned(3990, 12), 1288 => to_unsigned(2741, 12), 1289 => to_unsigned(2146, 12), 1290 => to_unsigned(193, 12), 1291 => to_unsigned(2950, 12), 1292 => to_unsigned(2565, 12), 1293 => to_unsigned(2400, 12), 1294 => to_unsigned(2094, 12), 1295 => to_unsigned(3785, 12), 1296 => to_unsigned(1321, 12), 1297 => to_unsigned(3288, 12), 1298 => to_unsigned(1904, 12), 1299 => to_unsigned(1139, 12), 1300 => to_unsigned(2721, 12), 1301 => to_unsigned(804, 12), 1302 => to_unsigned(1838, 12), 1303 => to_unsigned(363, 12), 1304 => to_unsigned(4084, 12), 1305 => to_unsigned(3147, 12), 1306 => to_unsigned(2412, 12), 1307 => to_unsigned(1393, 12), 1308 => to_unsigned(2496, 12), 1309 => to_unsigned(290, 12), 1310 => to_unsigned(188, 12), 1311 => to_unsigned(780, 12), 1312 => to_unsigned(1721, 12), 1313 => to_unsigned(2469, 12), 1314 => to_unsigned(2496, 12), 1315 => to_unsigned(2132, 12), 1316 => to_unsigned(555, 12), 1317 => to_unsigned(2751, 12), 1318 => to_unsigned(3269, 12), 1319 => to_unsigned(1777, 12), 1320 => to_unsigned(977, 12), 1321 => to_unsigned(3873, 12), 1322 => to_unsigned(2209, 12), 1323 => to_unsigned(2631, 12), 1324 => to_unsigned(1267, 12), 1325 => to_unsigned(2250, 12), 1326 => to_unsigned(3655, 12), 1327 => to_unsigned(3563, 12), 1328 => to_unsigned(1666, 12), 1329 => to_unsigned(3139, 12), 1330 => to_unsigned(3852, 12), 1331 => to_unsigned(682, 12), 1332 => to_unsigned(3598, 12), 1333 => to_unsigned(2082, 12), 1334 => to_unsigned(2403, 12), 1335 => to_unsigned(3221, 12), 1336 => to_unsigned(3991, 12), 1337 => to_unsigned(136, 12), 1338 => to_unsigned(2032, 12), 1339 => to_unsigned(1689, 12), 1340 => to_unsigned(1932, 12), 1341 => to_unsigned(809, 12), 1342 => to_unsigned(3753, 12), 1343 => to_unsigned(2022, 12), 1344 => to_unsigned(1318, 12), 1345 => to_unsigned(3710, 12), 1346 => to_unsigned(3193, 12), 1347 => to_unsigned(3759, 12), 1348 => to_unsigned(2443, 12), 1349 => to_unsigned(518, 12), 1350 => to_unsigned(971, 12), 1351 => to_unsigned(911, 12), 1352 => to_unsigned(337, 12), 1353 => to_unsigned(3060, 12), 1354 => to_unsigned(146, 12), 1355 => to_unsigned(2804, 12), 1356 => to_unsigned(1541, 12), 1357 => to_unsigned(2170, 12), 1358 => to_unsigned(3471, 12), 1359 => to_unsigned(2053, 12), 1360 => to_unsigned(2891, 12), 1361 => to_unsigned(2659, 12), 1362 => to_unsigned(3011, 12), 1363 => to_unsigned(929, 12), 1364 => to_unsigned(2089, 12), 1365 => to_unsigned(720, 12), 1366 => to_unsigned(2703, 12), 1367 => to_unsigned(3628, 12), 1368 => to_unsigned(254, 12), 1369 => to_unsigned(1261, 12), 1370 => to_unsigned(792, 12), 1371 => to_unsigned(674, 12), 1372 => to_unsigned(1470, 12), 1373 => to_unsigned(3780, 12), 1374 => to_unsigned(2440, 12), 1375 => to_unsigned(2224, 12), 1376 => to_unsigned(2227, 12), 1377 => to_unsigned(2852, 12), 1378 => to_unsigned(602, 12), 1379 => to_unsigned(2219, 12), 1380 => to_unsigned(1345, 12), 1381 => to_unsigned(273, 12), 1382 => to_unsigned(2744, 12), 1383 => to_unsigned(650, 12), 1384 => to_unsigned(1287, 12), 1385 => to_unsigned(1733, 12), 1386 => to_unsigned(922, 12), 1387 => to_unsigned(1467, 12), 1388 => to_unsigned(2058, 12), 1389 => to_unsigned(409, 12), 1390 => to_unsigned(1190, 12), 1391 => to_unsigned(2382, 12), 1392 => to_unsigned(2990, 12), 1393 => to_unsigned(251, 12), 1394 => to_unsigned(4057, 12), 1395 => to_unsigned(2101, 12), 1396 => to_unsigned(2284, 12), 1397 => to_unsigned(2496, 12), 1398 => to_unsigned(630, 12), 1399 => to_unsigned(3293, 12), 1400 => to_unsigned(3579, 12), 1401 => to_unsigned(3978, 12), 1402 => to_unsigned(1749, 12), 1403 => to_unsigned(547, 12), 1404 => to_unsigned(3509, 12), 1405 => to_unsigned(2613, 12), 1406 => to_unsigned(956, 12), 1407 => to_unsigned(725, 12), 1408 => to_unsigned(4060, 12), 1409 => to_unsigned(638, 12), 1410 => to_unsigned(2073, 12), 1411 => to_unsigned(191, 12), 1412 => to_unsigned(1668, 12), 1413 => to_unsigned(1869, 12), 1414 => to_unsigned(1743, 12), 1415 => to_unsigned(2058, 12), 1416 => to_unsigned(1303, 12), 1417 => to_unsigned(3045, 12), 1418 => to_unsigned(2920, 12), 1419 => to_unsigned(3713, 12), 1420 => to_unsigned(954, 12), 1421 => to_unsigned(2883, 12), 1422 => to_unsigned(3612, 12), 1423 => to_unsigned(3213, 12), 1424 => to_unsigned(717, 12), 1425 => to_unsigned(2560, 12), 1426 => to_unsigned(318, 12), 1427 => to_unsigned(66, 12), 1428 => to_unsigned(3255, 12), 1429 => to_unsigned(378, 12), 1430 => to_unsigned(3390, 12), 1431 => to_unsigned(733, 12), 1432 => to_unsigned(1896, 12), 1433 => to_unsigned(2874, 12), 1434 => to_unsigned(1740, 12), 1435 => to_unsigned(2301, 12), 1436 => to_unsigned(3550, 12), 1437 => to_unsigned(2333, 12), 1438 => to_unsigned(2712, 12), 1439 => to_unsigned(1718, 12), 1440 => to_unsigned(1277, 12), 1441 => to_unsigned(1525, 12), 1442 => to_unsigned(2294, 12), 1443 => to_unsigned(2253, 12), 1444 => to_unsigned(3070, 12), 1445 => to_unsigned(778, 12), 1446 => to_unsigned(157, 12), 1447 => to_unsigned(2498, 12), 1448 => to_unsigned(2813, 12), 1449 => to_unsigned(3271, 12), 1450 => to_unsigned(3836, 12), 1451 => to_unsigned(1091, 12), 1452 => to_unsigned(2864, 12), 1453 => to_unsigned(860, 12), 1454 => to_unsigned(228, 12), 1455 => to_unsigned(623, 12), 1456 => to_unsigned(509, 12), 1457 => to_unsigned(2208, 12), 1458 => to_unsigned(894, 12), 1459 => to_unsigned(2666, 12), 1460 => to_unsigned(1965, 12), 1461 => to_unsigned(4023, 12), 1462 => to_unsigned(2029, 12), 1463 => to_unsigned(399, 12), 1464 => to_unsigned(1654, 12), 1465 => to_unsigned(3448, 12), 1466 => to_unsigned(1472, 12), 1467 => to_unsigned(682, 12), 1468 => to_unsigned(3231, 12), 1469 => to_unsigned(2197, 12), 1470 => to_unsigned(3209, 12), 1471 => to_unsigned(436, 12), 1472 => to_unsigned(1456, 12), 1473 => to_unsigned(1293, 12), 1474 => to_unsigned(2423, 12), 1475 => to_unsigned(599, 12), 1476 => to_unsigned(3380, 12), 1477 => to_unsigned(2451, 12), 1478 => to_unsigned(2009, 12), 1479 => to_unsigned(3084, 12), 1480 => to_unsigned(2917, 12), 1481 => to_unsigned(2071, 12), 1482 => to_unsigned(2805, 12), 1483 => to_unsigned(2946, 12), 1484 => to_unsigned(2118, 12), 1485 => to_unsigned(3543, 12), 1486 => to_unsigned(1116, 12), 1487 => to_unsigned(962, 12), 1488 => to_unsigned(3831, 12), 1489 => to_unsigned(1968, 12), 1490 => to_unsigned(596, 12), 1491 => to_unsigned(1336, 12), 1492 => to_unsigned(2273, 12), 1493 => to_unsigned(2032, 12), 1494 => to_unsigned(1956, 12), 1495 => to_unsigned(290, 12), 1496 => to_unsigned(2725, 12), 1497 => to_unsigned(1131, 12), 1498 => to_unsigned(1690, 12), 1499 => to_unsigned(2978, 12), 1500 => to_unsigned(3445, 12), 1501 => to_unsigned(3941, 12), 1502 => to_unsigned(1107, 12), 1503 => to_unsigned(2167, 12), 1504 => to_unsigned(572, 12), 1505 => to_unsigned(1950, 12), 1506 => to_unsigned(2871, 12), 1507 => to_unsigned(401, 12), 1508 => to_unsigned(2062, 12), 1509 => to_unsigned(396, 12), 1510 => to_unsigned(1734, 12), 1511 => to_unsigned(3621, 12), 1512 => to_unsigned(592, 12), 1513 => to_unsigned(1688, 12), 1514 => to_unsigned(1856, 12), 1515 => to_unsigned(990, 12), 1516 => to_unsigned(3819, 12), 1517 => to_unsigned(3791, 12), 1518 => to_unsigned(3856, 12), 1519 => to_unsigned(1115, 12), 1520 => to_unsigned(3114, 12), 1521 => to_unsigned(3332, 12), 1522 => to_unsigned(1020, 12), 1523 => to_unsigned(1787, 12), 1524 => to_unsigned(1061, 12), 1525 => to_unsigned(329, 12), 1526 => to_unsigned(70, 12), 1527 => to_unsigned(2587, 12), 1528 => to_unsigned(3872, 12), 1529 => to_unsigned(3614, 12), 1530 => to_unsigned(3702, 12), 1531 => to_unsigned(3488, 12), 1532 => to_unsigned(3492, 12), 1533 => to_unsigned(2843, 12), 1534 => to_unsigned(1638, 12), 1535 => to_unsigned(1094, 12), 1536 => to_unsigned(583, 12), 1537 => to_unsigned(2428, 12), 1538 => to_unsigned(1569, 12), 1539 => to_unsigned(205, 12), 1540 => to_unsigned(692, 12), 1541 => to_unsigned(1924, 12), 1542 => to_unsigned(1094, 12), 1543 => to_unsigned(2777, 12), 1544 => to_unsigned(3689, 12), 1545 => to_unsigned(1398, 12), 1546 => to_unsigned(2008, 12), 1547 => to_unsigned(4014, 12), 1548 => to_unsigned(1343, 12), 1549 => to_unsigned(1140, 12), 1550 => to_unsigned(3250, 12), 1551 => to_unsigned(1774, 12), 1552 => to_unsigned(1681, 12), 1553 => to_unsigned(3019, 12), 1554 => to_unsigned(125, 12), 1555 => to_unsigned(1177, 12), 1556 => to_unsigned(3698, 12), 1557 => to_unsigned(2575, 12), 1558 => to_unsigned(1619, 12), 1559 => to_unsigned(136, 12), 1560 => to_unsigned(1167, 12), 1561 => to_unsigned(3740, 12), 1562 => to_unsigned(1307, 12), 1563 => to_unsigned(1892, 12), 1564 => to_unsigned(3837, 12), 1565 => to_unsigned(316, 12), 1566 => to_unsigned(3828, 12), 1567 => to_unsigned(896, 12), 1568 => to_unsigned(3476, 12), 1569 => to_unsigned(3186, 12), 1570 => to_unsigned(707, 12), 1571 => to_unsigned(3700, 12), 1572 => to_unsigned(1556, 12), 1573 => to_unsigned(821, 12), 1574 => to_unsigned(600, 12), 1575 => to_unsigned(257, 12), 1576 => to_unsigned(3902, 12), 1577 => to_unsigned(3452, 12), 1578 => to_unsigned(1506, 12), 1579 => to_unsigned(556, 12), 1580 => to_unsigned(1119, 12), 1581 => to_unsigned(342, 12), 1582 => to_unsigned(547, 12), 1583 => to_unsigned(994, 12), 1584 => to_unsigned(1470, 12), 1585 => to_unsigned(3527, 12), 1586 => to_unsigned(3474, 12), 1587 => to_unsigned(2512, 12), 1588 => to_unsigned(3615, 12), 1589 => to_unsigned(2044, 12), 1590 => to_unsigned(1046, 12), 1591 => to_unsigned(3021, 12), 1592 => to_unsigned(3268, 12), 1593 => to_unsigned(583, 12), 1594 => to_unsigned(334, 12), 1595 => to_unsigned(1282, 12), 1596 => to_unsigned(1241, 12), 1597 => to_unsigned(1626, 12), 1598 => to_unsigned(3323, 12), 1599 => to_unsigned(2221, 12), 1600 => to_unsigned(1390, 12), 1601 => to_unsigned(3911, 12), 1602 => to_unsigned(2485, 12), 1603 => to_unsigned(2702, 12), 1604 => to_unsigned(1998, 12), 1605 => to_unsigned(436, 12), 1606 => to_unsigned(2306, 12), 1607 => to_unsigned(4044, 12), 1608 => to_unsigned(1517, 12), 1609 => to_unsigned(1153, 12), 1610 => to_unsigned(3896, 12), 1611 => to_unsigned(1122, 12), 1612 => to_unsigned(2563, 12), 1613 => to_unsigned(1357, 12), 1614 => to_unsigned(3599, 12), 1615 => to_unsigned(2563, 12), 1616 => to_unsigned(730, 12), 1617 => to_unsigned(2206, 12), 1618 => to_unsigned(2145, 12), 1619 => to_unsigned(939, 12), 1620 => to_unsigned(677, 12), 1621 => to_unsigned(899, 12), 1622 => to_unsigned(3456, 12), 1623 => to_unsigned(1533, 12), 1624 => to_unsigned(1068, 12), 1625 => to_unsigned(2207, 12), 1626 => to_unsigned(3450, 12), 1627 => to_unsigned(1240, 12), 1628 => to_unsigned(2646, 12), 1629 => to_unsigned(1312, 12), 1630 => to_unsigned(497, 12), 1631 => to_unsigned(834, 12), 1632 => to_unsigned(2472, 12), 1633 => to_unsigned(1481, 12), 1634 => to_unsigned(3621, 12), 1635 => to_unsigned(1762, 12), 1636 => to_unsigned(1442, 12), 1637 => to_unsigned(4094, 12), 1638 => to_unsigned(3660, 12), 1639 => to_unsigned(545, 12), 1640 => to_unsigned(79, 12), 1641 => to_unsigned(939, 12), 1642 => to_unsigned(1880, 12), 1643 => to_unsigned(1291, 12), 1644 => to_unsigned(615, 12), 1645 => to_unsigned(3571, 12), 1646 => to_unsigned(3020, 12), 1647 => to_unsigned(3281, 12), 1648 => to_unsigned(2747, 12), 1649 => to_unsigned(2754, 12), 1650 => to_unsigned(1, 12), 1651 => to_unsigned(3975, 12), 1652 => to_unsigned(922, 12), 1653 => to_unsigned(58, 12), 1654 => to_unsigned(791, 12), 1655 => to_unsigned(258, 12), 1656 => to_unsigned(37, 12), 1657 => to_unsigned(606, 12), 1658 => to_unsigned(1503, 12), 1659 => to_unsigned(2357, 12), 1660 => to_unsigned(2701, 12), 1661 => to_unsigned(872, 12), 1662 => to_unsigned(3532, 12), 1663 => to_unsigned(133, 12), 1664 => to_unsigned(1079, 12), 1665 => to_unsigned(1756, 12), 1666 => to_unsigned(2059, 12), 1667 => to_unsigned(3046, 12), 1668 => to_unsigned(2704, 12), 1669 => to_unsigned(1670, 12), 1670 => to_unsigned(4035, 12), 1671 => to_unsigned(4048, 12), 1672 => to_unsigned(1790, 12), 1673 => to_unsigned(363, 12), 1674 => to_unsigned(1646, 12), 1675 => to_unsigned(800, 12), 1676 => to_unsigned(2519, 12), 1677 => to_unsigned(1110, 12), 1678 => to_unsigned(2241, 12), 1679 => to_unsigned(2588, 12), 1680 => to_unsigned(1283, 12), 1681 => to_unsigned(2622, 12), 1682 => to_unsigned(496, 12), 1683 => to_unsigned(2868, 12), 1684 => to_unsigned(368, 12), 1685 => to_unsigned(1629, 12), 1686 => to_unsigned(1971, 12), 1687 => to_unsigned(2131, 12), 1688 => to_unsigned(3093, 12), 1689 => to_unsigned(1177, 12), 1690 => to_unsigned(2863, 12), 1691 => to_unsigned(3092, 12), 1692 => to_unsigned(533, 12), 1693 => to_unsigned(334, 12), 1694 => to_unsigned(3826, 12), 1695 => to_unsigned(1266, 12), 1696 => to_unsigned(2863, 12), 1697 => to_unsigned(3404, 12), 1698 => to_unsigned(2177, 12), 1699 => to_unsigned(2148, 12), 1700 => to_unsigned(4022, 12), 1701 => to_unsigned(2123, 12), 1702 => to_unsigned(3355, 12), 1703 => to_unsigned(2853, 12), 1704 => to_unsigned(3941, 12), 1705 => to_unsigned(1099, 12), 1706 => to_unsigned(1980, 12), 1707 => to_unsigned(3242, 12), 1708 => to_unsigned(511, 12), 1709 => to_unsigned(318, 12), 1710 => to_unsigned(46, 12), 1711 => to_unsigned(833, 12), 1712 => to_unsigned(1508, 12), 1713 => to_unsigned(896, 12), 1714 => to_unsigned(1859, 12), 1715 => to_unsigned(3689, 12), 1716 => to_unsigned(2270, 12), 1717 => to_unsigned(483, 12), 1718 => to_unsigned(55, 12), 1719 => to_unsigned(2268, 12), 1720 => to_unsigned(842, 12), 1721 => to_unsigned(3009, 12), 1722 => to_unsigned(4093, 12), 1723 => to_unsigned(3746, 12), 1724 => to_unsigned(4029, 12), 1725 => to_unsigned(1046, 12), 1726 => to_unsigned(3774, 12), 1727 => to_unsigned(1155, 12), 1728 => to_unsigned(434, 12), 1729 => to_unsigned(3487, 12), 1730 => to_unsigned(692, 12), 1731 => to_unsigned(2317, 12), 1732 => to_unsigned(1096, 12), 1733 => to_unsigned(1103, 12), 1734 => to_unsigned(161, 12), 1735 => to_unsigned(286, 12), 1736 => to_unsigned(4058, 12), 1737 => to_unsigned(1396, 12), 1738 => to_unsigned(3063, 12), 1739 => to_unsigned(3097, 12), 1740 => to_unsigned(2887, 12), 1741 => to_unsigned(824, 12), 1742 => to_unsigned(1912, 12), 1743 => to_unsigned(3841, 12), 1744 => to_unsigned(660, 12), 1745 => to_unsigned(3538, 12), 1746 => to_unsigned(2948, 12), 1747 => to_unsigned(680, 12), 1748 => to_unsigned(2181, 12), 1749 => to_unsigned(697, 12), 1750 => to_unsigned(3665, 12), 1751 => to_unsigned(4042, 12), 1752 => to_unsigned(3616, 12), 1753 => to_unsigned(2174, 12), 1754 => to_unsigned(1610, 12), 1755 => to_unsigned(2939, 12), 1756 => to_unsigned(2559, 12), 1757 => to_unsigned(732, 12), 1758 => to_unsigned(2883, 12), 1759 => to_unsigned(3890, 12), 1760 => to_unsigned(3706, 12), 1761 => to_unsigned(2020, 12), 1762 => to_unsigned(2491, 12), 1763 => to_unsigned(1584, 12), 1764 => to_unsigned(826, 12), 1765 => to_unsigned(3629, 12), 1766 => to_unsigned(3249, 12), 1767 => to_unsigned(31, 12), 1768 => to_unsigned(3113, 12), 1769 => to_unsigned(3698, 12), 1770 => to_unsigned(1255, 12), 1771 => to_unsigned(1663, 12), 1772 => to_unsigned(2254, 12), 1773 => to_unsigned(977, 12), 1774 => to_unsigned(3663, 12), 1775 => to_unsigned(2406, 12), 1776 => to_unsigned(2621, 12), 1777 => to_unsigned(3085, 12), 1778 => to_unsigned(1616, 12), 1779 => to_unsigned(1324, 12), 1780 => to_unsigned(1771, 12), 1781 => to_unsigned(2501, 12), 1782 => to_unsigned(2015, 12), 1783 => to_unsigned(3640, 12), 1784 => to_unsigned(3025, 12), 1785 => to_unsigned(3619, 12), 1786 => to_unsigned(3549, 12), 1787 => to_unsigned(1749, 12), 1788 => to_unsigned(3875, 12), 1789 => to_unsigned(2419, 12), 1790 => to_unsigned(826, 12), 1791 => to_unsigned(2371, 12), 1792 => to_unsigned(791, 12), 1793 => to_unsigned(450, 12), 1794 => to_unsigned(2140, 12), 1795 => to_unsigned(3784, 12), 1796 => to_unsigned(518, 12), 1797 => to_unsigned(3332, 12), 1798 => to_unsigned(3066, 12), 1799 => to_unsigned(3302, 12), 1800 => to_unsigned(1835, 12), 1801 => to_unsigned(3770, 12), 1802 => to_unsigned(3774, 12), 1803 => to_unsigned(2972, 12), 1804 => to_unsigned(1878, 12), 1805 => to_unsigned(2026, 12), 1806 => to_unsigned(2304, 12), 1807 => to_unsigned(905, 12), 1808 => to_unsigned(1348, 12), 1809 => to_unsigned(3582, 12), 1810 => to_unsigned(884, 12), 1811 => to_unsigned(3068, 12), 1812 => to_unsigned(3377, 12), 1813 => to_unsigned(2337, 12), 1814 => to_unsigned(1314, 12), 1815 => to_unsigned(2397, 12), 1816 => to_unsigned(3550, 12), 1817 => to_unsigned(1673, 12), 1818 => to_unsigned(2815, 12), 1819 => to_unsigned(2364, 12), 1820 => to_unsigned(2982, 12), 1821 => to_unsigned(3741, 12), 1822 => to_unsigned(1696, 12), 1823 => to_unsigned(487, 12), 1824 => to_unsigned(3251, 12), 1825 => to_unsigned(2493, 12), 1826 => to_unsigned(2790, 12), 1827 => to_unsigned(2113, 12), 1828 => to_unsigned(592, 12), 1829 => to_unsigned(2899, 12), 1830 => to_unsigned(2791, 12), 1831 => to_unsigned(3101, 12), 1832 => to_unsigned(2782, 12), 1833 => to_unsigned(601, 12), 1834 => to_unsigned(2674, 12), 1835 => to_unsigned(2880, 12), 1836 => to_unsigned(144, 12), 1837 => to_unsigned(2656, 12), 1838 => to_unsigned(2355, 12), 1839 => to_unsigned(2690, 12), 1840 => to_unsigned(2517, 12), 1841 => to_unsigned(1018, 12), 1842 => to_unsigned(2653, 12), 1843 => to_unsigned(252, 12), 1844 => to_unsigned(985, 12), 1845 => to_unsigned(676, 12), 1846 => to_unsigned(2237, 12), 1847 => to_unsigned(3653, 12), 1848 => to_unsigned(2122, 12), 1849 => to_unsigned(3611, 12), 1850 => to_unsigned(2796, 12), 1851 => to_unsigned(4023, 12), 1852 => to_unsigned(2324, 12), 1853 => to_unsigned(1832, 12), 1854 => to_unsigned(433, 12), 1855 => to_unsigned(3713, 12), 1856 => to_unsigned(2132, 12), 1857 => to_unsigned(2063, 12), 1858 => to_unsigned(358, 12), 1859 => to_unsigned(3581, 12), 1860 => to_unsigned(138, 12), 1861 => to_unsigned(2676, 12), 1862 => to_unsigned(2910, 12), 1863 => to_unsigned(1040, 12), 1864 => to_unsigned(960, 12), 1865 => to_unsigned(1161, 12), 1866 => to_unsigned(3483, 12), 1867 => to_unsigned(2663, 12), 1868 => to_unsigned(275, 12), 1869 => to_unsigned(1227, 12), 1870 => to_unsigned(2453, 12), 1871 => to_unsigned(3593, 12), 1872 => to_unsigned(2417, 12), 1873 => to_unsigned(3084, 12), 1874 => to_unsigned(4089, 12), 1875 => to_unsigned(138, 12), 1876 => to_unsigned(763, 12), 1877 => to_unsigned(3277, 12), 1878 => to_unsigned(2109, 12), 1879 => to_unsigned(1579, 12), 1880 => to_unsigned(1225, 12), 1881 => to_unsigned(3592, 12), 1882 => to_unsigned(2761, 12), 1883 => to_unsigned(1266, 12), 1884 => to_unsigned(2389, 12), 1885 => to_unsigned(2057, 12), 1886 => to_unsigned(2790, 12), 1887 => to_unsigned(3487, 12), 1888 => to_unsigned(1028, 12), 1889 => to_unsigned(886, 12), 1890 => to_unsigned(2426, 12), 1891 => to_unsigned(960, 12), 1892 => to_unsigned(784, 12), 1893 => to_unsigned(3872, 12), 1894 => to_unsigned(1405, 12), 1895 => to_unsigned(1471, 12), 1896 => to_unsigned(3997, 12), 1897 => to_unsigned(804, 12), 1898 => to_unsigned(4014, 12), 1899 => to_unsigned(1673, 12), 1900 => to_unsigned(3681, 12), 1901 => to_unsigned(1759, 12), 1902 => to_unsigned(971, 12), 1903 => to_unsigned(2477, 12), 1904 => to_unsigned(1696, 12), 1905 => to_unsigned(2642, 12), 1906 => to_unsigned(3032, 12), 1907 => to_unsigned(152, 12), 1908 => to_unsigned(4016, 12), 1909 => to_unsigned(3899, 12), 1910 => to_unsigned(2981, 12), 1911 => to_unsigned(2899, 12), 1912 => to_unsigned(2086, 12), 1913 => to_unsigned(1680, 12), 1914 => to_unsigned(1213, 12), 1915 => to_unsigned(2322, 12), 1916 => to_unsigned(2275, 12), 1917 => to_unsigned(624, 12), 1918 => to_unsigned(335, 12), 1919 => to_unsigned(3274, 12), 1920 => to_unsigned(3041, 12), 1921 => to_unsigned(1115, 12), 1922 => to_unsigned(735, 12), 1923 => to_unsigned(347, 12), 1924 => to_unsigned(2713, 12), 1925 => to_unsigned(137, 12), 1926 => to_unsigned(3413, 12), 1927 => to_unsigned(1973, 12), 1928 => to_unsigned(2257, 12), 1929 => to_unsigned(2693, 12), 1930 => to_unsigned(2277, 12), 1931 => to_unsigned(2873, 12), 1932 => to_unsigned(69, 12), 1933 => to_unsigned(3269, 12), 1934 => to_unsigned(738, 12), 1935 => to_unsigned(1968, 12), 1936 => to_unsigned(2828, 12), 1937 => to_unsigned(3025, 12), 1938 => to_unsigned(2540, 12), 1939 => to_unsigned(598, 12), 1940 => to_unsigned(58, 12), 1941 => to_unsigned(3221, 12), 1942 => to_unsigned(2161, 12), 1943 => to_unsigned(1890, 12), 1944 => to_unsigned(2168, 12), 1945 => to_unsigned(546, 12), 1946 => to_unsigned(1764, 12), 1947 => to_unsigned(3441, 12), 1948 => to_unsigned(1468, 12), 1949 => to_unsigned(809, 12), 1950 => to_unsigned(3724, 12), 1951 => to_unsigned(155, 12), 1952 => to_unsigned(699, 12), 1953 => to_unsigned(27, 12), 1954 => to_unsigned(901, 12), 1955 => to_unsigned(1420, 12), 1956 => to_unsigned(2628, 12), 1957 => to_unsigned(3831, 12), 1958 => to_unsigned(63, 12), 1959 => to_unsigned(1524, 12), 1960 => to_unsigned(980, 12), 1961 => to_unsigned(1727, 12), 1962 => to_unsigned(2434, 12), 1963 => to_unsigned(2584, 12), 1964 => to_unsigned(1551, 12), 1965 => to_unsigned(1233, 12), 1966 => to_unsigned(1374, 12), 1967 => to_unsigned(525, 12), 1968 => to_unsigned(939, 12), 1969 => to_unsigned(1369, 12), 1970 => to_unsigned(1467, 12), 1971 => to_unsigned(3932, 12), 1972 => to_unsigned(3381, 12), 1973 => to_unsigned(3471, 12), 1974 => to_unsigned(1284, 12), 1975 => to_unsigned(2112, 12), 1976 => to_unsigned(3170, 12), 1977 => to_unsigned(505, 12), 1978 => to_unsigned(1744, 12), 1979 => to_unsigned(2210, 12), 1980 => to_unsigned(1161, 12), 1981 => to_unsigned(709, 12), 1982 => to_unsigned(329, 12), 1983 => to_unsigned(262, 12), 1984 => to_unsigned(2242, 12), 1985 => to_unsigned(2944, 12), 1986 => to_unsigned(3382, 12), 1987 => to_unsigned(801, 12), 1988 => to_unsigned(480, 12), 1989 => to_unsigned(1113, 12), 1990 => to_unsigned(2369, 12), 1991 => to_unsigned(2740, 12), 1992 => to_unsigned(2791, 12), 1993 => to_unsigned(3622, 12), 1994 => to_unsigned(3929, 12), 1995 => to_unsigned(1792, 12), 1996 => to_unsigned(3511, 12), 1997 => to_unsigned(3449, 12), 1998 => to_unsigned(3864, 12), 1999 => to_unsigned(732, 12), 2000 => to_unsigned(703, 12), 2001 => to_unsigned(2302, 12), 2002 => to_unsigned(3080, 12), 2003 => to_unsigned(1307, 12), 2004 => to_unsigned(2311, 12), 2005 => to_unsigned(188, 12), 2006 => to_unsigned(2983, 12), 2007 => to_unsigned(643, 12), 2008 => to_unsigned(1650, 12), 2009 => to_unsigned(1380, 12), 2010 => to_unsigned(1801, 12), 2011 => to_unsigned(3390, 12), 2012 => to_unsigned(1048, 12), 2013 => to_unsigned(1983, 12), 2014 => to_unsigned(1273, 12), 2015 => to_unsigned(3821, 12), 2016 => to_unsigned(1260, 12), 2017 => to_unsigned(2022, 12), 2018 => to_unsigned(2262, 12), 2019 => to_unsigned(2755, 12), 2020 => to_unsigned(3697, 12), 2021 => to_unsigned(3059, 12), 2022 => to_unsigned(584, 12), 2023 => to_unsigned(745, 12), 2024 => to_unsigned(1713, 12), 2025 => to_unsigned(1268, 12), 2026 => to_unsigned(3220, 12), 2027 => to_unsigned(668, 12), 2028 => to_unsigned(2764, 12), 2029 => to_unsigned(1331, 12), 2030 => to_unsigned(3246, 12), 2031 => to_unsigned(1231, 12), 2032 => to_unsigned(3801, 12), 2033 => to_unsigned(2820, 12), 2034 => to_unsigned(556, 12), 2035 => to_unsigned(3095, 12), 2036 => to_unsigned(2996, 12), 2037 => to_unsigned(2239, 12), 2038 => to_unsigned(27, 12), 2039 => to_unsigned(2290, 12), 2040 => to_unsigned(3768, 12), 2041 => to_unsigned(2192, 12), 2042 => to_unsigned(3199, 12), 2043 => to_unsigned(3557, 12), 2044 => to_unsigned(979, 12), 2045 => to_unsigned(3646, 12), 2046 => to_unsigned(2357, 12), 2047 => to_unsigned(17, 12)),
            9 => (0 => to_unsigned(1508, 12), 1 => to_unsigned(1628, 12), 2 => to_unsigned(1646, 12), 3 => to_unsigned(1189, 12), 4 => to_unsigned(3987, 12), 5 => to_unsigned(3406, 12), 6 => to_unsigned(868, 12), 7 => to_unsigned(2805, 12), 8 => to_unsigned(2164, 12), 9 => to_unsigned(25, 12), 10 => to_unsigned(472, 12), 11 => to_unsigned(2499, 12), 12 => to_unsigned(1660, 12), 13 => to_unsigned(1812, 12), 14 => to_unsigned(3888, 12), 15 => to_unsigned(1513, 12), 16 => to_unsigned(3755, 12), 17 => to_unsigned(2706, 12), 18 => to_unsigned(2092, 12), 19 => to_unsigned(1837, 12), 20 => to_unsigned(2140, 12), 21 => to_unsigned(3144, 12), 22 => to_unsigned(565, 12), 23 => to_unsigned(2343, 12), 24 => to_unsigned(2254, 12), 25 => to_unsigned(3617, 12), 26 => to_unsigned(3544, 12), 27 => to_unsigned(2137, 12), 28 => to_unsigned(2962, 12), 29 => to_unsigned(2926, 12), 30 => to_unsigned(1219, 12), 31 => to_unsigned(2583, 12), 32 => to_unsigned(50, 12), 33 => to_unsigned(3580, 12), 34 => to_unsigned(354, 12), 35 => to_unsigned(3732, 12), 36 => to_unsigned(1839, 12), 37 => to_unsigned(3304, 12), 38 => to_unsigned(350, 12), 39 => to_unsigned(89, 12), 40 => to_unsigned(2532, 12), 41 => to_unsigned(1706, 12), 42 => to_unsigned(1809, 12), 43 => to_unsigned(2133, 12), 44 => to_unsigned(1340, 12), 45 => to_unsigned(2244, 12), 46 => to_unsigned(3763, 12), 47 => to_unsigned(2657, 12), 48 => to_unsigned(199, 12), 49 => to_unsigned(35, 12), 50 => to_unsigned(264, 12), 51 => to_unsigned(1325, 12), 52 => to_unsigned(581, 12), 53 => to_unsigned(71, 12), 54 => to_unsigned(3746, 12), 55 => to_unsigned(3576, 12), 56 => to_unsigned(1048, 12), 57 => to_unsigned(321, 12), 58 => to_unsigned(2145, 12), 59 => to_unsigned(2971, 12), 60 => to_unsigned(3205, 12), 61 => to_unsigned(3089, 12), 62 => to_unsigned(56, 12), 63 => to_unsigned(2147, 12), 64 => to_unsigned(2331, 12), 65 => to_unsigned(1631, 12), 66 => to_unsigned(3022, 12), 67 => to_unsigned(1740, 12), 68 => to_unsigned(556, 12), 69 => to_unsigned(2219, 12), 70 => to_unsigned(3258, 12), 71 => to_unsigned(3865, 12), 72 => to_unsigned(1123, 12), 73 => to_unsigned(2312, 12), 74 => to_unsigned(2866, 12), 75 => to_unsigned(3257, 12), 76 => to_unsigned(2731, 12), 77 => to_unsigned(2637, 12), 78 => to_unsigned(1299, 12), 79 => to_unsigned(3128, 12), 80 => to_unsigned(1072, 12), 81 => to_unsigned(2541, 12), 82 => to_unsigned(1740, 12), 83 => to_unsigned(3515, 12), 84 => to_unsigned(2894, 12), 85 => to_unsigned(898, 12), 86 => to_unsigned(888, 12), 87 => to_unsigned(1834, 12), 88 => to_unsigned(423, 12), 89 => to_unsigned(1780, 12), 90 => to_unsigned(673, 12), 91 => to_unsigned(2672, 12), 92 => to_unsigned(3762, 12), 93 => to_unsigned(950, 12), 94 => to_unsigned(274, 12), 95 => to_unsigned(1267, 12), 96 => to_unsigned(798, 12), 97 => to_unsigned(1927, 12), 98 => to_unsigned(4044, 12), 99 => to_unsigned(1395, 12), 100 => to_unsigned(3661, 12), 101 => to_unsigned(1742, 12), 102 => to_unsigned(1492, 12), 103 => to_unsigned(315, 12), 104 => to_unsigned(3539, 12), 105 => to_unsigned(3182, 12), 106 => to_unsigned(3624, 12), 107 => to_unsigned(3817, 12), 108 => to_unsigned(845, 12), 109 => to_unsigned(1992, 12), 110 => to_unsigned(402, 12), 111 => to_unsigned(3009, 12), 112 => to_unsigned(3470, 12), 113 => to_unsigned(3817, 12), 114 => to_unsigned(3588, 12), 115 => to_unsigned(1546, 12), 116 => to_unsigned(354, 12), 117 => to_unsigned(1407, 12), 118 => to_unsigned(2744, 12), 119 => to_unsigned(2534, 12), 120 => to_unsigned(1398, 12), 121 => to_unsigned(3750, 12), 122 => to_unsigned(4023, 12), 123 => to_unsigned(3106, 12), 124 => to_unsigned(375, 12), 125 => to_unsigned(3925, 12), 126 => to_unsigned(1673, 12), 127 => to_unsigned(421, 12), 128 => to_unsigned(3388, 12), 129 => to_unsigned(2626, 12), 130 => to_unsigned(532, 12), 131 => to_unsigned(2130, 12), 132 => to_unsigned(453, 12), 133 => to_unsigned(1615, 12), 134 => to_unsigned(922, 12), 135 => to_unsigned(4078, 12), 136 => to_unsigned(210, 12), 137 => to_unsigned(1072, 12), 138 => to_unsigned(2047, 12), 139 => to_unsigned(884, 12), 140 => to_unsigned(3887, 12), 141 => to_unsigned(3202, 12), 142 => to_unsigned(2593, 12), 143 => to_unsigned(3005, 12), 144 => to_unsigned(1613, 12), 145 => to_unsigned(1174, 12), 146 => to_unsigned(1871, 12), 147 => to_unsigned(3037, 12), 148 => to_unsigned(1286, 12), 149 => to_unsigned(786, 12), 150 => to_unsigned(2718, 12), 151 => to_unsigned(983, 12), 152 => to_unsigned(2662, 12), 153 => to_unsigned(476, 12), 154 => to_unsigned(633, 12), 155 => to_unsigned(73, 12), 156 => to_unsigned(2443, 12), 157 => to_unsigned(3482, 12), 158 => to_unsigned(3892, 12), 159 => to_unsigned(3036, 12), 160 => to_unsigned(2361, 12), 161 => to_unsigned(2794, 12), 162 => to_unsigned(2211, 12), 163 => to_unsigned(265, 12), 164 => to_unsigned(61, 12), 165 => to_unsigned(2806, 12), 166 => to_unsigned(3979, 12), 167 => to_unsigned(3346, 12), 168 => to_unsigned(2588, 12), 169 => to_unsigned(229, 12), 170 => to_unsigned(2795, 12), 171 => to_unsigned(299, 12), 172 => to_unsigned(1291, 12), 173 => to_unsigned(1129, 12), 174 => to_unsigned(148, 12), 175 => to_unsigned(249, 12), 176 => to_unsigned(1194, 12), 177 => to_unsigned(1393, 12), 178 => to_unsigned(257, 12), 179 => to_unsigned(1554, 12), 180 => to_unsigned(783, 12), 181 => to_unsigned(2858, 12), 182 => to_unsigned(1823, 12), 183 => to_unsigned(2617, 12), 184 => to_unsigned(2157, 12), 185 => to_unsigned(2646, 12), 186 => to_unsigned(809, 12), 187 => to_unsigned(3132, 12), 188 => to_unsigned(110, 12), 189 => to_unsigned(2076, 12), 190 => to_unsigned(2268, 12), 191 => to_unsigned(3439, 12), 192 => to_unsigned(2983, 12), 193 => to_unsigned(2296, 12), 194 => to_unsigned(3498, 12), 195 => to_unsigned(1522, 12), 196 => to_unsigned(3321, 12), 197 => to_unsigned(2121, 12), 198 => to_unsigned(1175, 12), 199 => to_unsigned(1734, 12), 200 => to_unsigned(2151, 12), 201 => to_unsigned(1098, 12), 202 => to_unsigned(3657, 12), 203 => to_unsigned(514, 12), 204 => to_unsigned(1458, 12), 205 => to_unsigned(1377, 12), 206 => to_unsigned(2638, 12), 207 => to_unsigned(349, 12), 208 => to_unsigned(2378, 12), 209 => to_unsigned(3128, 12), 210 => to_unsigned(2496, 12), 211 => to_unsigned(2472, 12), 212 => to_unsigned(3168, 12), 213 => to_unsigned(470, 12), 214 => to_unsigned(1930, 12), 215 => to_unsigned(3271, 12), 216 => to_unsigned(3259, 12), 217 => to_unsigned(85, 12), 218 => to_unsigned(3304, 12), 219 => to_unsigned(2351, 12), 220 => to_unsigned(1469, 12), 221 => to_unsigned(106, 12), 222 => to_unsigned(1836, 12), 223 => to_unsigned(3092, 12), 224 => to_unsigned(3505, 12), 225 => to_unsigned(1702, 12), 226 => to_unsigned(144, 12), 227 => to_unsigned(2385, 12), 228 => to_unsigned(3543, 12), 229 => to_unsigned(2808, 12), 230 => to_unsigned(295, 12), 231 => to_unsigned(949, 12), 232 => to_unsigned(1248, 12), 233 => to_unsigned(2414, 12), 234 => to_unsigned(2535, 12), 235 => to_unsigned(3070, 12), 236 => to_unsigned(241, 12), 237 => to_unsigned(320, 12), 238 => to_unsigned(462, 12), 239 => to_unsigned(451, 12), 240 => to_unsigned(1349, 12), 241 => to_unsigned(1654, 12), 242 => to_unsigned(549, 12), 243 => to_unsigned(2059, 12), 244 => to_unsigned(2113, 12), 245 => to_unsigned(3, 12), 246 => to_unsigned(2299, 12), 247 => to_unsigned(3142, 12), 248 => to_unsigned(1314, 12), 249 => to_unsigned(699, 12), 250 => to_unsigned(1513, 12), 251 => to_unsigned(1371, 12), 252 => to_unsigned(3858, 12), 253 => to_unsigned(3081, 12), 254 => to_unsigned(3945, 12), 255 => to_unsigned(2043, 12), 256 => to_unsigned(2148, 12), 257 => to_unsigned(2317, 12), 258 => to_unsigned(2162, 12), 259 => to_unsigned(216, 12), 260 => to_unsigned(1255, 12), 261 => to_unsigned(4078, 12), 262 => to_unsigned(3655, 12), 263 => to_unsigned(1113, 12), 264 => to_unsigned(845, 12), 265 => to_unsigned(798, 12), 266 => to_unsigned(1862, 12), 267 => to_unsigned(4018, 12), 268 => to_unsigned(3208, 12), 269 => to_unsigned(3305, 12), 270 => to_unsigned(3891, 12), 271 => to_unsigned(3866, 12), 272 => to_unsigned(2698, 12), 273 => to_unsigned(2338, 12), 274 => to_unsigned(821, 12), 275 => to_unsigned(3609, 12), 276 => to_unsigned(68, 12), 277 => to_unsigned(1903, 12), 278 => to_unsigned(3466, 12), 279 => to_unsigned(1613, 12), 280 => to_unsigned(1118, 12), 281 => to_unsigned(830, 12), 282 => to_unsigned(2815, 12), 283 => to_unsigned(1119, 12), 284 => to_unsigned(1186, 12), 285 => to_unsigned(2150, 12), 286 => to_unsigned(1495, 12), 287 => to_unsigned(2865, 12), 288 => to_unsigned(318, 12), 289 => to_unsigned(492, 12), 290 => to_unsigned(226, 12), 291 => to_unsigned(2936, 12), 292 => to_unsigned(1360, 12), 293 => to_unsigned(2582, 12), 294 => to_unsigned(1177, 12), 295 => to_unsigned(1227, 12), 296 => to_unsigned(519, 12), 297 => to_unsigned(3065, 12), 298 => to_unsigned(2686, 12), 299 => to_unsigned(3252, 12), 300 => to_unsigned(2756, 12), 301 => to_unsigned(156, 12), 302 => to_unsigned(3801, 12), 303 => to_unsigned(2660, 12), 304 => to_unsigned(361, 12), 305 => to_unsigned(3018, 12), 306 => to_unsigned(3575, 12), 307 => to_unsigned(403, 12), 308 => to_unsigned(1274, 12), 309 => to_unsigned(1813, 12), 310 => to_unsigned(2038, 12), 311 => to_unsigned(3479, 12), 312 => to_unsigned(3103, 12), 313 => to_unsigned(93, 12), 314 => to_unsigned(237, 12), 315 => to_unsigned(2229, 12), 316 => to_unsigned(1888, 12), 317 => to_unsigned(2603, 12), 318 => to_unsigned(3092, 12), 319 => to_unsigned(1406, 12), 320 => to_unsigned(1872, 12), 321 => to_unsigned(1, 12), 322 => to_unsigned(1284, 12), 323 => to_unsigned(3701, 12), 324 => to_unsigned(158, 12), 325 => to_unsigned(3677, 12), 326 => to_unsigned(3566, 12), 327 => to_unsigned(2088, 12), 328 => to_unsigned(2953, 12), 329 => to_unsigned(1085, 12), 330 => to_unsigned(1889, 12), 331 => to_unsigned(1, 12), 332 => to_unsigned(281, 12), 333 => to_unsigned(976, 12), 334 => to_unsigned(1050, 12), 335 => to_unsigned(1633, 12), 336 => to_unsigned(329, 12), 337 => to_unsigned(3111, 12), 338 => to_unsigned(923, 12), 339 => to_unsigned(2364, 12), 340 => to_unsigned(4038, 12), 341 => to_unsigned(1512, 12), 342 => to_unsigned(2906, 12), 343 => to_unsigned(2972, 12), 344 => to_unsigned(3905, 12), 345 => to_unsigned(725, 12), 346 => to_unsigned(2384, 12), 347 => to_unsigned(2385, 12), 348 => to_unsigned(198, 12), 349 => to_unsigned(2089, 12), 350 => to_unsigned(61, 12), 351 => to_unsigned(941, 12), 352 => to_unsigned(81, 12), 353 => to_unsigned(489, 12), 354 => to_unsigned(2181, 12), 355 => to_unsigned(225, 12), 356 => to_unsigned(1860, 12), 357 => to_unsigned(492, 12), 358 => to_unsigned(1129, 12), 359 => to_unsigned(2591, 12), 360 => to_unsigned(1705, 12), 361 => to_unsigned(2231, 12), 362 => to_unsigned(229, 12), 363 => to_unsigned(2990, 12), 364 => to_unsigned(3438, 12), 365 => to_unsigned(3475, 12), 366 => to_unsigned(1956, 12), 367 => to_unsigned(487, 12), 368 => to_unsigned(1798, 12), 369 => to_unsigned(2942, 12), 370 => to_unsigned(2164, 12), 371 => to_unsigned(1577, 12), 372 => to_unsigned(3149, 12), 373 => to_unsigned(3009, 12), 374 => to_unsigned(1478, 12), 375 => to_unsigned(3738, 12), 376 => to_unsigned(1704, 12), 377 => to_unsigned(2690, 12), 378 => to_unsigned(2380, 12), 379 => to_unsigned(3415, 12), 380 => to_unsigned(3758, 12), 381 => to_unsigned(1108, 12), 382 => to_unsigned(1586, 12), 383 => to_unsigned(2537, 12), 384 => to_unsigned(241, 12), 385 => to_unsigned(195, 12), 386 => to_unsigned(1283, 12), 387 => to_unsigned(101, 12), 388 => to_unsigned(2322, 12), 389 => to_unsigned(1087, 12), 390 => to_unsigned(2692, 12), 391 => to_unsigned(3824, 12), 392 => to_unsigned(3308, 12), 393 => to_unsigned(1159, 12), 394 => to_unsigned(401, 12), 395 => to_unsigned(305, 12), 396 => to_unsigned(3739, 12), 397 => to_unsigned(3121, 12), 398 => to_unsigned(3168, 12), 399 => to_unsigned(2522, 12), 400 => to_unsigned(2254, 12), 401 => to_unsigned(1521, 12), 402 => to_unsigned(2637, 12), 403 => to_unsigned(1802, 12), 404 => to_unsigned(3239, 12), 405 => to_unsigned(985, 12), 406 => to_unsigned(863, 12), 407 => to_unsigned(1323, 12), 408 => to_unsigned(2837, 12), 409 => to_unsigned(2345, 12), 410 => to_unsigned(125, 12), 411 => to_unsigned(1674, 12), 412 => to_unsigned(1706, 12), 413 => to_unsigned(2537, 12), 414 => to_unsigned(1603, 12), 415 => to_unsigned(4038, 12), 416 => to_unsigned(4010, 12), 417 => to_unsigned(2512, 12), 418 => to_unsigned(3103, 12), 419 => to_unsigned(1214, 12), 420 => to_unsigned(2113, 12), 421 => to_unsigned(2262, 12), 422 => to_unsigned(938, 12), 423 => to_unsigned(225, 12), 424 => to_unsigned(135, 12), 425 => to_unsigned(3384, 12), 426 => to_unsigned(2050, 12), 427 => to_unsigned(3231, 12), 428 => to_unsigned(3737, 12), 429 => to_unsigned(3763, 12), 430 => to_unsigned(1097, 12), 431 => to_unsigned(1323, 12), 432 => to_unsigned(225, 12), 433 => to_unsigned(3621, 12), 434 => to_unsigned(3941, 12), 435 => to_unsigned(2178, 12), 436 => to_unsigned(3768, 12), 437 => to_unsigned(357, 12), 438 => to_unsigned(3435, 12), 439 => to_unsigned(1075, 12), 440 => to_unsigned(3571, 12), 441 => to_unsigned(3139, 12), 442 => to_unsigned(1508, 12), 443 => to_unsigned(2007, 12), 444 => to_unsigned(3110, 12), 445 => to_unsigned(3784, 12), 446 => to_unsigned(3507, 12), 447 => to_unsigned(1539, 12), 448 => to_unsigned(356, 12), 449 => to_unsigned(1819, 12), 450 => to_unsigned(1485, 12), 451 => to_unsigned(1486, 12), 452 => to_unsigned(1309, 12), 453 => to_unsigned(2163, 12), 454 => to_unsigned(823, 12), 455 => to_unsigned(1692, 12), 456 => to_unsigned(112, 12), 457 => to_unsigned(1342, 12), 458 => to_unsigned(3434, 12), 459 => to_unsigned(1602, 12), 460 => to_unsigned(412, 12), 461 => to_unsigned(2513, 12), 462 => to_unsigned(3366, 12), 463 => to_unsigned(513, 12), 464 => to_unsigned(1627, 12), 465 => to_unsigned(2406, 12), 466 => to_unsigned(287, 12), 467 => to_unsigned(2958, 12), 468 => to_unsigned(1191, 12), 469 => to_unsigned(3774, 12), 470 => to_unsigned(359, 12), 471 => to_unsigned(1402, 12), 472 => to_unsigned(1980, 12), 473 => to_unsigned(3957, 12), 474 => to_unsigned(1658, 12), 475 => to_unsigned(1635, 12), 476 => to_unsigned(2012, 12), 477 => to_unsigned(456, 12), 478 => to_unsigned(902, 12), 479 => to_unsigned(1221, 12), 480 => to_unsigned(4073, 12), 481 => to_unsigned(1463, 12), 482 => to_unsigned(2604, 12), 483 => to_unsigned(1945, 12), 484 => to_unsigned(3586, 12), 485 => to_unsigned(2778, 12), 486 => to_unsigned(2540, 12), 487 => to_unsigned(1402, 12), 488 => to_unsigned(1679, 12), 489 => to_unsigned(69, 12), 490 => to_unsigned(2390, 12), 491 => to_unsigned(778, 12), 492 => to_unsigned(3200, 12), 493 => to_unsigned(311, 12), 494 => to_unsigned(2197, 12), 495 => to_unsigned(2440, 12), 496 => to_unsigned(3936, 12), 497 => to_unsigned(529, 12), 498 => to_unsigned(2828, 12), 499 => to_unsigned(415, 12), 500 => to_unsigned(381, 12), 501 => to_unsigned(1526, 12), 502 => to_unsigned(3123, 12), 503 => to_unsigned(3302, 12), 504 => to_unsigned(961, 12), 505 => to_unsigned(2404, 12), 506 => to_unsigned(1460, 12), 507 => to_unsigned(1835, 12), 508 => to_unsigned(4051, 12), 509 => to_unsigned(1289, 12), 510 => to_unsigned(2862, 12), 511 => to_unsigned(2770, 12), 512 => to_unsigned(2295, 12), 513 => to_unsigned(1337, 12), 514 => to_unsigned(2246, 12), 515 => to_unsigned(995, 12), 516 => to_unsigned(102, 12), 517 => to_unsigned(3813, 12), 518 => to_unsigned(2662, 12), 519 => to_unsigned(2125, 12), 520 => to_unsigned(3587, 12), 521 => to_unsigned(547, 12), 522 => to_unsigned(449, 12), 523 => to_unsigned(2826, 12), 524 => to_unsigned(3478, 12), 525 => to_unsigned(1521, 12), 526 => to_unsigned(248, 12), 527 => to_unsigned(2446, 12), 528 => to_unsigned(1557, 12), 529 => to_unsigned(449, 12), 530 => to_unsigned(2916, 12), 531 => to_unsigned(1712, 12), 532 => to_unsigned(132, 12), 533 => to_unsigned(2158, 12), 534 => to_unsigned(2509, 12), 535 => to_unsigned(1538, 12), 536 => to_unsigned(3686, 12), 537 => to_unsigned(3298, 12), 538 => to_unsigned(1559, 12), 539 => to_unsigned(1518, 12), 540 => to_unsigned(2208, 12), 541 => to_unsigned(1228, 12), 542 => to_unsigned(237, 12), 543 => to_unsigned(3650, 12), 544 => to_unsigned(3178, 12), 545 => to_unsigned(2419, 12), 546 => to_unsigned(2248, 12), 547 => to_unsigned(354, 12), 548 => to_unsigned(1281, 12), 549 => to_unsigned(19, 12), 550 => to_unsigned(2520, 12), 551 => to_unsigned(1882, 12), 552 => to_unsigned(1074, 12), 553 => to_unsigned(3760, 12), 554 => to_unsigned(932, 12), 555 => to_unsigned(2769, 12), 556 => to_unsigned(863, 12), 557 => to_unsigned(3477, 12), 558 => to_unsigned(2722, 12), 559 => to_unsigned(2257, 12), 560 => to_unsigned(2980, 12), 561 => to_unsigned(3898, 12), 562 => to_unsigned(2913, 12), 563 => to_unsigned(2698, 12), 564 => to_unsigned(1284, 12), 565 => to_unsigned(410, 12), 566 => to_unsigned(1372, 12), 567 => to_unsigned(1776, 12), 568 => to_unsigned(114, 12), 569 => to_unsigned(2656, 12), 570 => to_unsigned(3291, 12), 571 => to_unsigned(2716, 12), 572 => to_unsigned(97, 12), 573 => to_unsigned(1291, 12), 574 => to_unsigned(759, 12), 575 => to_unsigned(1103, 12), 576 => to_unsigned(2676, 12), 577 => to_unsigned(1468, 12), 578 => to_unsigned(3182, 12), 579 => to_unsigned(935, 12), 580 => to_unsigned(99, 12), 581 => to_unsigned(295, 12), 582 => to_unsigned(372, 12), 583 => to_unsigned(2736, 12), 584 => to_unsigned(1208, 12), 585 => to_unsigned(1304, 12), 586 => to_unsigned(433, 12), 587 => to_unsigned(1091, 12), 588 => to_unsigned(2100, 12), 589 => to_unsigned(3181, 12), 590 => to_unsigned(2882, 12), 591 => to_unsigned(3934, 12), 592 => to_unsigned(3034, 12), 593 => to_unsigned(493, 12), 594 => to_unsigned(3936, 12), 595 => to_unsigned(1771, 12), 596 => to_unsigned(961, 12), 597 => to_unsigned(1800, 12), 598 => to_unsigned(3729, 12), 599 => to_unsigned(2638, 12), 600 => to_unsigned(466, 12), 601 => to_unsigned(2844, 12), 602 => to_unsigned(3537, 12), 603 => to_unsigned(417, 12), 604 => to_unsigned(2007, 12), 605 => to_unsigned(2004, 12), 606 => to_unsigned(1471, 12), 607 => to_unsigned(1649, 12), 608 => to_unsigned(458, 12), 609 => to_unsigned(2895, 12), 610 => to_unsigned(2942, 12), 611 => to_unsigned(2521, 12), 612 => to_unsigned(1735, 12), 613 => to_unsigned(436, 12), 614 => to_unsigned(3272, 12), 615 => to_unsigned(3636, 12), 616 => to_unsigned(246, 12), 617 => to_unsigned(1175, 12), 618 => to_unsigned(2431, 12), 619 => to_unsigned(2842, 12), 620 => to_unsigned(98, 12), 621 => to_unsigned(698, 12), 622 => to_unsigned(3908, 12), 623 => to_unsigned(2521, 12), 624 => to_unsigned(2784, 12), 625 => to_unsigned(1458, 12), 626 => to_unsigned(763, 12), 627 => to_unsigned(628, 12), 628 => to_unsigned(338, 12), 629 => to_unsigned(2014, 12), 630 => to_unsigned(685, 12), 631 => to_unsigned(1398, 12), 632 => to_unsigned(48, 12), 633 => to_unsigned(948, 12), 634 => to_unsigned(3135, 12), 635 => to_unsigned(2654, 12), 636 => to_unsigned(1037, 12), 637 => to_unsigned(3214, 12), 638 => to_unsigned(4027, 12), 639 => to_unsigned(1702, 12), 640 => to_unsigned(2168, 12), 641 => to_unsigned(630, 12), 642 => to_unsigned(1379, 12), 643 => to_unsigned(3760, 12), 644 => to_unsigned(1460, 12), 645 => to_unsigned(2564, 12), 646 => to_unsigned(768, 12), 647 => to_unsigned(1584, 12), 648 => to_unsigned(1995, 12), 649 => to_unsigned(2653, 12), 650 => to_unsigned(1398, 12), 651 => to_unsigned(3578, 12), 652 => to_unsigned(1739, 12), 653 => to_unsigned(3122, 12), 654 => to_unsigned(2094, 12), 655 => to_unsigned(246, 12), 656 => to_unsigned(3582, 12), 657 => to_unsigned(299, 12), 658 => to_unsigned(3416, 12), 659 => to_unsigned(2771, 12), 660 => to_unsigned(895, 12), 661 => to_unsigned(2939, 12), 662 => to_unsigned(168, 12), 663 => to_unsigned(3158, 12), 664 => to_unsigned(3104, 12), 665 => to_unsigned(3758, 12), 666 => to_unsigned(3196, 12), 667 => to_unsigned(2162, 12), 668 => to_unsigned(780, 12), 669 => to_unsigned(1691, 12), 670 => to_unsigned(2951, 12), 671 => to_unsigned(372, 12), 672 => to_unsigned(1293, 12), 673 => to_unsigned(843, 12), 674 => to_unsigned(1410, 12), 675 => to_unsigned(945, 12), 676 => to_unsigned(2051, 12), 677 => to_unsigned(3868, 12), 678 => to_unsigned(4024, 12), 679 => to_unsigned(2239, 12), 680 => to_unsigned(2101, 12), 681 => to_unsigned(1929, 12), 682 => to_unsigned(250, 12), 683 => to_unsigned(2733, 12), 684 => to_unsigned(444, 12), 685 => to_unsigned(1847, 12), 686 => to_unsigned(1436, 12), 687 => to_unsigned(1342, 12), 688 => to_unsigned(2835, 12), 689 => to_unsigned(2039, 12), 690 => to_unsigned(3508, 12), 691 => to_unsigned(727, 12), 692 => to_unsigned(1715, 12), 693 => to_unsigned(3547, 12), 694 => to_unsigned(2917, 12), 695 => to_unsigned(838, 12), 696 => to_unsigned(1684, 12), 697 => to_unsigned(3151, 12), 698 => to_unsigned(1754, 12), 699 => to_unsigned(213, 12), 700 => to_unsigned(2812, 12), 701 => to_unsigned(725, 12), 702 => to_unsigned(1424, 12), 703 => to_unsigned(515, 12), 704 => to_unsigned(2268, 12), 705 => to_unsigned(2547, 12), 706 => to_unsigned(1908, 12), 707 => to_unsigned(838, 12), 708 => to_unsigned(3158, 12), 709 => to_unsigned(27, 12), 710 => to_unsigned(658, 12), 711 => to_unsigned(3287, 12), 712 => to_unsigned(90, 12), 713 => to_unsigned(2956, 12), 714 => to_unsigned(3259, 12), 715 => to_unsigned(1148, 12), 716 => to_unsigned(135, 12), 717 => to_unsigned(1097, 12), 718 => to_unsigned(1795, 12), 719 => to_unsigned(2270, 12), 720 => to_unsigned(655, 12), 721 => to_unsigned(2311, 12), 722 => to_unsigned(3060, 12), 723 => to_unsigned(3289, 12), 724 => to_unsigned(2462, 12), 725 => to_unsigned(1048, 12), 726 => to_unsigned(1265, 12), 727 => to_unsigned(118, 12), 728 => to_unsigned(931, 12), 729 => to_unsigned(163, 12), 730 => to_unsigned(1088, 12), 731 => to_unsigned(3874, 12), 732 => to_unsigned(3654, 12), 733 => to_unsigned(1839, 12), 734 => to_unsigned(1325, 12), 735 => to_unsigned(3587, 12), 736 => to_unsigned(3782, 12), 737 => to_unsigned(3890, 12), 738 => to_unsigned(2296, 12), 739 => to_unsigned(1366, 12), 740 => to_unsigned(1383, 12), 741 => to_unsigned(1528, 12), 742 => to_unsigned(496, 12), 743 => to_unsigned(391, 12), 744 => to_unsigned(2845, 12), 745 => to_unsigned(670, 12), 746 => to_unsigned(3725, 12), 747 => to_unsigned(259, 12), 748 => to_unsigned(835, 12), 749 => to_unsigned(3884, 12), 750 => to_unsigned(3506, 12), 751 => to_unsigned(934, 12), 752 => to_unsigned(1089, 12), 753 => to_unsigned(994, 12), 754 => to_unsigned(3987, 12), 755 => to_unsigned(3023, 12), 756 => to_unsigned(1142, 12), 757 => to_unsigned(2064, 12), 758 => to_unsigned(4015, 12), 759 => to_unsigned(1879, 12), 760 => to_unsigned(1576, 12), 761 => to_unsigned(4087, 12), 762 => to_unsigned(3191, 12), 763 => to_unsigned(2146, 12), 764 => to_unsigned(15, 12), 765 => to_unsigned(2865, 12), 766 => to_unsigned(2621, 12), 767 => to_unsigned(1250, 12), 768 => to_unsigned(2103, 12), 769 => to_unsigned(1903, 12), 770 => to_unsigned(2763, 12), 771 => to_unsigned(2810, 12), 772 => to_unsigned(1092, 12), 773 => to_unsigned(2461, 12), 774 => to_unsigned(136, 12), 775 => to_unsigned(1995, 12), 776 => to_unsigned(3024, 12), 777 => to_unsigned(3393, 12), 778 => to_unsigned(47, 12), 779 => to_unsigned(209, 12), 780 => to_unsigned(2413, 12), 781 => to_unsigned(2911, 12), 782 => to_unsigned(2664, 12), 783 => to_unsigned(1773, 12), 784 => to_unsigned(1530, 12), 785 => to_unsigned(2165, 12), 786 => to_unsigned(509, 12), 787 => to_unsigned(1038, 12), 788 => to_unsigned(766, 12), 789 => to_unsigned(2734, 12), 790 => to_unsigned(824, 12), 791 => to_unsigned(2043, 12), 792 => to_unsigned(4026, 12), 793 => to_unsigned(2673, 12), 794 => to_unsigned(3144, 12), 795 => to_unsigned(65, 12), 796 => to_unsigned(1371, 12), 797 => to_unsigned(3051, 12), 798 => to_unsigned(2761, 12), 799 => to_unsigned(2625, 12), 800 => to_unsigned(3971, 12), 801 => to_unsigned(2736, 12), 802 => to_unsigned(1533, 12), 803 => to_unsigned(2623, 12), 804 => to_unsigned(3758, 12), 805 => to_unsigned(1953, 12), 806 => to_unsigned(1025, 12), 807 => to_unsigned(2339, 12), 808 => to_unsigned(3320, 12), 809 => to_unsigned(3521, 12), 810 => to_unsigned(2785, 12), 811 => to_unsigned(2500, 12), 812 => to_unsigned(1535, 12), 813 => to_unsigned(922, 12), 814 => to_unsigned(1714, 12), 815 => to_unsigned(1051, 12), 816 => to_unsigned(3442, 12), 817 => to_unsigned(943, 12), 818 => to_unsigned(778, 12), 819 => to_unsigned(3732, 12), 820 => to_unsigned(2421, 12), 821 => to_unsigned(2086, 12), 822 => to_unsigned(472, 12), 823 => to_unsigned(68, 12), 824 => to_unsigned(1997, 12), 825 => to_unsigned(2906, 12), 826 => to_unsigned(2283, 12), 827 => to_unsigned(3517, 12), 828 => to_unsigned(2213, 12), 829 => to_unsigned(255, 12), 830 => to_unsigned(178, 12), 831 => to_unsigned(586, 12), 832 => to_unsigned(2347, 12), 833 => to_unsigned(3100, 12), 834 => to_unsigned(427, 12), 835 => to_unsigned(1034, 12), 836 => to_unsigned(1751, 12), 837 => to_unsigned(1598, 12), 838 => to_unsigned(3044, 12), 839 => to_unsigned(519, 12), 840 => to_unsigned(2927, 12), 841 => to_unsigned(1649, 12), 842 => to_unsigned(3153, 12), 843 => to_unsigned(2740, 12), 844 => to_unsigned(3904, 12), 845 => to_unsigned(1024, 12), 846 => to_unsigned(2378, 12), 847 => to_unsigned(758, 12), 848 => to_unsigned(283, 12), 849 => to_unsigned(1793, 12), 850 => to_unsigned(1524, 12), 851 => to_unsigned(2507, 12), 852 => to_unsigned(2554, 12), 853 => to_unsigned(4062, 12), 854 => to_unsigned(1062, 12), 855 => to_unsigned(3195, 12), 856 => to_unsigned(2224, 12), 857 => to_unsigned(3138, 12), 858 => to_unsigned(799, 12), 859 => to_unsigned(318, 12), 860 => to_unsigned(3342, 12), 861 => to_unsigned(75, 12), 862 => to_unsigned(443, 12), 863 => to_unsigned(1749, 12), 864 => to_unsigned(2742, 12), 865 => to_unsigned(3837, 12), 866 => to_unsigned(3911, 12), 867 => to_unsigned(588, 12), 868 => to_unsigned(2804, 12), 869 => to_unsigned(2864, 12), 870 => to_unsigned(1707, 12), 871 => to_unsigned(1393, 12), 872 => to_unsigned(1776, 12), 873 => to_unsigned(1029, 12), 874 => to_unsigned(1213, 12), 875 => to_unsigned(961, 12), 876 => to_unsigned(2209, 12), 877 => to_unsigned(229, 12), 878 => to_unsigned(2752, 12), 879 => to_unsigned(1068, 12), 880 => to_unsigned(815, 12), 881 => to_unsigned(1217, 12), 882 => to_unsigned(1554, 12), 883 => to_unsigned(859, 12), 884 => to_unsigned(1919, 12), 885 => to_unsigned(2674, 12), 886 => to_unsigned(904, 12), 887 => to_unsigned(3629, 12), 888 => to_unsigned(1779, 12), 889 => to_unsigned(2382, 12), 890 => to_unsigned(2840, 12), 891 => to_unsigned(3064, 12), 892 => to_unsigned(1554, 12), 893 => to_unsigned(9, 12), 894 => to_unsigned(955, 12), 895 => to_unsigned(3993, 12), 896 => to_unsigned(3902, 12), 897 => to_unsigned(2043, 12), 898 => to_unsigned(1177, 12), 899 => to_unsigned(4007, 12), 900 => to_unsigned(1560, 12), 901 => to_unsigned(1780, 12), 902 => to_unsigned(488, 12), 903 => to_unsigned(2092, 12), 904 => to_unsigned(2561, 12), 905 => to_unsigned(3590, 12), 906 => to_unsigned(2350, 12), 907 => to_unsigned(299, 12), 908 => to_unsigned(3491, 12), 909 => to_unsigned(1630, 12), 910 => to_unsigned(497, 12), 911 => to_unsigned(4083, 12), 912 => to_unsigned(751, 12), 913 => to_unsigned(708, 12), 914 => to_unsigned(2028, 12), 915 => to_unsigned(209, 12), 916 => to_unsigned(648, 12), 917 => to_unsigned(1652, 12), 918 => to_unsigned(3752, 12), 919 => to_unsigned(1091, 12), 920 => to_unsigned(2918, 12), 921 => to_unsigned(2151, 12), 922 => to_unsigned(3957, 12), 923 => to_unsigned(2049, 12), 924 => to_unsigned(1024, 12), 925 => to_unsigned(732, 12), 926 => to_unsigned(3887, 12), 927 => to_unsigned(2164, 12), 928 => to_unsigned(2722, 12), 929 => to_unsigned(3217, 12), 930 => to_unsigned(3138, 12), 931 => to_unsigned(1178, 12), 932 => to_unsigned(1572, 12), 933 => to_unsigned(2071, 12), 934 => to_unsigned(1216, 12), 935 => to_unsigned(1246, 12), 936 => to_unsigned(3905, 12), 937 => to_unsigned(836, 12), 938 => to_unsigned(4054, 12), 939 => to_unsigned(731, 12), 940 => to_unsigned(2438, 12), 941 => to_unsigned(381, 12), 942 => to_unsigned(765, 12), 943 => to_unsigned(2264, 12), 944 => to_unsigned(2005, 12), 945 => to_unsigned(1834, 12), 946 => to_unsigned(1278, 12), 947 => to_unsigned(747, 12), 948 => to_unsigned(1146, 12), 949 => to_unsigned(2359, 12), 950 => to_unsigned(1780, 12), 951 => to_unsigned(1540, 12), 952 => to_unsigned(1443, 12), 953 => to_unsigned(935, 12), 954 => to_unsigned(1379, 12), 955 => to_unsigned(3969, 12), 956 => to_unsigned(4074, 12), 957 => to_unsigned(2216, 12), 958 => to_unsigned(1815, 12), 959 => to_unsigned(1705, 12), 960 => to_unsigned(2179, 12), 961 => to_unsigned(252, 12), 962 => to_unsigned(2076, 12), 963 => to_unsigned(2818, 12), 964 => to_unsigned(1455, 12), 965 => to_unsigned(3673, 12), 966 => to_unsigned(2775, 12), 967 => to_unsigned(1635, 12), 968 => to_unsigned(3800, 12), 969 => to_unsigned(1454, 12), 970 => to_unsigned(3831, 12), 971 => to_unsigned(2909, 12), 972 => to_unsigned(2430, 12), 973 => to_unsigned(312, 12), 974 => to_unsigned(3177, 12), 975 => to_unsigned(574, 12), 976 => to_unsigned(3749, 12), 977 => to_unsigned(319, 12), 978 => to_unsigned(2189, 12), 979 => to_unsigned(2196, 12), 980 => to_unsigned(505, 12), 981 => to_unsigned(3474, 12), 982 => to_unsigned(3365, 12), 983 => to_unsigned(134, 12), 984 => to_unsigned(1111, 12), 985 => to_unsigned(1546, 12), 986 => to_unsigned(3258, 12), 987 => to_unsigned(740, 12), 988 => to_unsigned(3649, 12), 989 => to_unsigned(1964, 12), 990 => to_unsigned(629, 12), 991 => to_unsigned(3432, 12), 992 => to_unsigned(595, 12), 993 => to_unsigned(1935, 12), 994 => to_unsigned(3275, 12), 995 => to_unsigned(639, 12), 996 => to_unsigned(3273, 12), 997 => to_unsigned(2028, 12), 998 => to_unsigned(1489, 12), 999 => to_unsigned(3626, 12), 1000 => to_unsigned(2985, 12), 1001 => to_unsigned(3865, 12), 1002 => to_unsigned(3652, 12), 1003 => to_unsigned(4047, 12), 1004 => to_unsigned(1922, 12), 1005 => to_unsigned(2303, 12), 1006 => to_unsigned(1113, 12), 1007 => to_unsigned(1543, 12), 1008 => to_unsigned(1655, 12), 1009 => to_unsigned(1599, 12), 1010 => to_unsigned(3690, 12), 1011 => to_unsigned(2065, 12), 1012 => to_unsigned(1904, 12), 1013 => to_unsigned(3452, 12), 1014 => to_unsigned(1546, 12), 1015 => to_unsigned(1699, 12), 1016 => to_unsigned(1957, 12), 1017 => to_unsigned(1790, 12), 1018 => to_unsigned(2903, 12), 1019 => to_unsigned(1833, 12), 1020 => to_unsigned(1391, 12), 1021 => to_unsigned(2525, 12), 1022 => to_unsigned(2938, 12), 1023 => to_unsigned(1839, 12), 1024 => to_unsigned(252, 12), 1025 => to_unsigned(1198, 12), 1026 => to_unsigned(1573, 12), 1027 => to_unsigned(2729, 12), 1028 => to_unsigned(1191, 12), 1029 => to_unsigned(2982, 12), 1030 => to_unsigned(2415, 12), 1031 => to_unsigned(889, 12), 1032 => to_unsigned(464, 12), 1033 => to_unsigned(1460, 12), 1034 => to_unsigned(2013, 12), 1035 => to_unsigned(1042, 12), 1036 => to_unsigned(1259, 12), 1037 => to_unsigned(3120, 12), 1038 => to_unsigned(1367, 12), 1039 => to_unsigned(3717, 12), 1040 => to_unsigned(3447, 12), 1041 => to_unsigned(504, 12), 1042 => to_unsigned(571, 12), 1043 => to_unsigned(182, 12), 1044 => to_unsigned(2038, 12), 1045 => to_unsigned(555, 12), 1046 => to_unsigned(3949, 12), 1047 => to_unsigned(524, 12), 1048 => to_unsigned(27, 12), 1049 => to_unsigned(911, 12), 1050 => to_unsigned(2459, 12), 1051 => to_unsigned(3181, 12), 1052 => to_unsigned(2960, 12), 1053 => to_unsigned(1722, 12), 1054 => to_unsigned(1841, 12), 1055 => to_unsigned(1510, 12), 1056 => to_unsigned(1466, 12), 1057 => to_unsigned(2335, 12), 1058 => to_unsigned(1458, 12), 1059 => to_unsigned(3460, 12), 1060 => to_unsigned(408, 12), 1061 => to_unsigned(664, 12), 1062 => to_unsigned(4044, 12), 1063 => to_unsigned(2742, 12), 1064 => to_unsigned(3182, 12), 1065 => to_unsigned(3873, 12), 1066 => to_unsigned(3451, 12), 1067 => to_unsigned(2689, 12), 1068 => to_unsigned(1100, 12), 1069 => to_unsigned(1859, 12), 1070 => to_unsigned(3161, 12), 1071 => to_unsigned(3631, 12), 1072 => to_unsigned(1426, 12), 1073 => to_unsigned(2228, 12), 1074 => to_unsigned(3219, 12), 1075 => to_unsigned(347, 12), 1076 => to_unsigned(3665, 12), 1077 => to_unsigned(2911, 12), 1078 => to_unsigned(2843, 12), 1079 => to_unsigned(20, 12), 1080 => to_unsigned(2933, 12), 1081 => to_unsigned(670, 12), 1082 => to_unsigned(2034, 12), 1083 => to_unsigned(429, 12), 1084 => to_unsigned(1874, 12), 1085 => to_unsigned(1522, 12), 1086 => to_unsigned(137, 12), 1087 => to_unsigned(1233, 12), 1088 => to_unsigned(3288, 12), 1089 => to_unsigned(96, 12), 1090 => to_unsigned(2619, 12), 1091 => to_unsigned(2575, 12), 1092 => to_unsigned(1141, 12), 1093 => to_unsigned(3798, 12), 1094 => to_unsigned(382, 12), 1095 => to_unsigned(1676, 12), 1096 => to_unsigned(2557, 12), 1097 => to_unsigned(2342, 12), 1098 => to_unsigned(3693, 12), 1099 => to_unsigned(2145, 12), 1100 => to_unsigned(135, 12), 1101 => to_unsigned(3331, 12), 1102 => to_unsigned(2643, 12), 1103 => to_unsigned(1840, 12), 1104 => to_unsigned(2764, 12), 1105 => to_unsigned(2725, 12), 1106 => to_unsigned(2105, 12), 1107 => to_unsigned(747, 12), 1108 => to_unsigned(2265, 12), 1109 => to_unsigned(2488, 12), 1110 => to_unsigned(313, 12), 1111 => to_unsigned(3980, 12), 1112 => to_unsigned(1918, 12), 1113 => to_unsigned(1336, 12), 1114 => to_unsigned(181, 12), 1115 => to_unsigned(1263, 12), 1116 => to_unsigned(2965, 12), 1117 => to_unsigned(496, 12), 1118 => to_unsigned(3833, 12), 1119 => to_unsigned(3379, 12), 1120 => to_unsigned(3843, 12), 1121 => to_unsigned(1629, 12), 1122 => to_unsigned(3535, 12), 1123 => to_unsigned(969, 12), 1124 => to_unsigned(600, 12), 1125 => to_unsigned(508, 12), 1126 => to_unsigned(2871, 12), 1127 => to_unsigned(1410, 12), 1128 => to_unsigned(3437, 12), 1129 => to_unsigned(3411, 12), 1130 => to_unsigned(2583, 12), 1131 => to_unsigned(3349, 12), 1132 => to_unsigned(571, 12), 1133 => to_unsigned(2650, 12), 1134 => to_unsigned(2154, 12), 1135 => to_unsigned(49, 12), 1136 => to_unsigned(1238, 12), 1137 => to_unsigned(2538, 12), 1138 => to_unsigned(3043, 12), 1139 => to_unsigned(1867, 12), 1140 => to_unsigned(2306, 12), 1141 => to_unsigned(945, 12), 1142 => to_unsigned(3948, 12), 1143 => to_unsigned(3796, 12), 1144 => to_unsigned(907, 12), 1145 => to_unsigned(2867, 12), 1146 => to_unsigned(3051, 12), 1147 => to_unsigned(3702, 12), 1148 => to_unsigned(3237, 12), 1149 => to_unsigned(1035, 12), 1150 => to_unsigned(1435, 12), 1151 => to_unsigned(2928, 12), 1152 => to_unsigned(500, 12), 1153 => to_unsigned(3776, 12), 1154 => to_unsigned(754, 12), 1155 => to_unsigned(1699, 12), 1156 => to_unsigned(3264, 12), 1157 => to_unsigned(2220, 12), 1158 => to_unsigned(995, 12), 1159 => to_unsigned(26, 12), 1160 => to_unsigned(3819, 12), 1161 => to_unsigned(3040, 12), 1162 => to_unsigned(3564, 12), 1163 => to_unsigned(1869, 12), 1164 => to_unsigned(1277, 12), 1165 => to_unsigned(761, 12), 1166 => to_unsigned(200, 12), 1167 => to_unsigned(2483, 12), 1168 => to_unsigned(3251, 12), 1169 => to_unsigned(59, 12), 1170 => to_unsigned(1168, 12), 1171 => to_unsigned(3518, 12), 1172 => to_unsigned(135, 12), 1173 => to_unsigned(3903, 12), 1174 => to_unsigned(1715, 12), 1175 => to_unsigned(3656, 12), 1176 => to_unsigned(384, 12), 1177 => to_unsigned(3342, 12), 1178 => to_unsigned(953, 12), 1179 => to_unsigned(3336, 12), 1180 => to_unsigned(426, 12), 1181 => to_unsigned(4059, 12), 1182 => to_unsigned(871, 12), 1183 => to_unsigned(116, 12), 1184 => to_unsigned(3092, 12), 1185 => to_unsigned(3746, 12), 1186 => to_unsigned(2200, 12), 1187 => to_unsigned(2, 12), 1188 => to_unsigned(1217, 12), 1189 => to_unsigned(535, 12), 1190 => to_unsigned(95, 12), 1191 => to_unsigned(1194, 12), 1192 => to_unsigned(3100, 12), 1193 => to_unsigned(1704, 12), 1194 => to_unsigned(1879, 12), 1195 => to_unsigned(1825, 12), 1196 => to_unsigned(500, 12), 1197 => to_unsigned(2778, 12), 1198 => to_unsigned(2764, 12), 1199 => to_unsigned(463, 12), 1200 => to_unsigned(1044, 12), 1201 => to_unsigned(1710, 12), 1202 => to_unsigned(4063, 12), 1203 => to_unsigned(3902, 12), 1204 => to_unsigned(2810, 12), 1205 => to_unsigned(139, 12), 1206 => to_unsigned(1379, 12), 1207 => to_unsigned(292, 12), 1208 => to_unsigned(3532, 12), 1209 => to_unsigned(3993, 12), 1210 => to_unsigned(3092, 12), 1211 => to_unsigned(3598, 12), 1212 => to_unsigned(2941, 12), 1213 => to_unsigned(1071, 12), 1214 => to_unsigned(1437, 12), 1215 => to_unsigned(718, 12), 1216 => to_unsigned(2783, 12), 1217 => to_unsigned(4043, 12), 1218 => to_unsigned(2671, 12), 1219 => to_unsigned(409, 12), 1220 => to_unsigned(1371, 12), 1221 => to_unsigned(2631, 12), 1222 => to_unsigned(204, 12), 1223 => to_unsigned(1280, 12), 1224 => to_unsigned(1757, 12), 1225 => to_unsigned(2197, 12), 1226 => to_unsigned(3718, 12), 1227 => to_unsigned(438, 12), 1228 => to_unsigned(1785, 12), 1229 => to_unsigned(1696, 12), 1230 => to_unsigned(559, 12), 1231 => to_unsigned(1495, 12), 1232 => to_unsigned(326, 12), 1233 => to_unsigned(994, 12), 1234 => to_unsigned(1876, 12), 1235 => to_unsigned(1923, 12), 1236 => to_unsigned(2977, 12), 1237 => to_unsigned(3906, 12), 1238 => to_unsigned(1705, 12), 1239 => to_unsigned(3781, 12), 1240 => to_unsigned(3012, 12), 1241 => to_unsigned(1179, 12), 1242 => to_unsigned(1932, 12), 1243 => to_unsigned(2769, 12), 1244 => to_unsigned(1815, 12), 1245 => to_unsigned(502, 12), 1246 => to_unsigned(714, 12), 1247 => to_unsigned(1786, 12), 1248 => to_unsigned(2743, 12), 1249 => to_unsigned(1361, 12), 1250 => to_unsigned(762, 12), 1251 => to_unsigned(726, 12), 1252 => to_unsigned(1188, 12), 1253 => to_unsigned(1258, 12), 1254 => to_unsigned(1056, 12), 1255 => to_unsigned(2325, 12), 1256 => to_unsigned(760, 12), 1257 => to_unsigned(1752, 12), 1258 => to_unsigned(804, 12), 1259 => to_unsigned(2561, 12), 1260 => to_unsigned(3191, 12), 1261 => to_unsigned(1557, 12), 1262 => to_unsigned(1358, 12), 1263 => to_unsigned(1968, 12), 1264 => to_unsigned(1900, 12), 1265 => to_unsigned(3587, 12), 1266 => to_unsigned(2451, 12), 1267 => to_unsigned(3377, 12), 1268 => to_unsigned(1422, 12), 1269 => to_unsigned(2602, 12), 1270 => to_unsigned(2618, 12), 1271 => to_unsigned(1649, 12), 1272 => to_unsigned(3831, 12), 1273 => to_unsigned(2534, 12), 1274 => to_unsigned(910, 12), 1275 => to_unsigned(2981, 12), 1276 => to_unsigned(3783, 12), 1277 => to_unsigned(1726, 12), 1278 => to_unsigned(3637, 12), 1279 => to_unsigned(2901, 12), 1280 => to_unsigned(2852, 12), 1281 => to_unsigned(1982, 12), 1282 => to_unsigned(1158, 12), 1283 => to_unsigned(1830, 12), 1284 => to_unsigned(1298, 12), 1285 => to_unsigned(1865, 12), 1286 => to_unsigned(1381, 12), 1287 => to_unsigned(2278, 12), 1288 => to_unsigned(3131, 12), 1289 => to_unsigned(2777, 12), 1290 => to_unsigned(4023, 12), 1291 => to_unsigned(2247, 12), 1292 => to_unsigned(3674, 12), 1293 => to_unsigned(1495, 12), 1294 => to_unsigned(1171, 12), 1295 => to_unsigned(979, 12), 1296 => to_unsigned(2821, 12), 1297 => to_unsigned(1847, 12), 1298 => to_unsigned(3380, 12), 1299 => to_unsigned(3387, 12), 1300 => to_unsigned(2556, 12), 1301 => to_unsigned(3110, 12), 1302 => to_unsigned(2475, 12), 1303 => to_unsigned(2551, 12), 1304 => to_unsigned(2329, 12), 1305 => to_unsigned(2406, 12), 1306 => to_unsigned(1077, 12), 1307 => to_unsigned(1659, 12), 1308 => to_unsigned(2690, 12), 1309 => to_unsigned(3603, 12), 1310 => to_unsigned(2095, 12), 1311 => to_unsigned(394, 12), 1312 => to_unsigned(1262, 12), 1313 => to_unsigned(4032, 12), 1314 => to_unsigned(3035, 12), 1315 => to_unsigned(578, 12), 1316 => to_unsigned(3253, 12), 1317 => to_unsigned(148, 12), 1318 => to_unsigned(764, 12), 1319 => to_unsigned(3270, 12), 1320 => to_unsigned(3500, 12), 1321 => to_unsigned(1151, 12), 1322 => to_unsigned(1835, 12), 1323 => to_unsigned(432, 12), 1324 => to_unsigned(3819, 12), 1325 => to_unsigned(2016, 12), 1326 => to_unsigned(2413, 12), 1327 => to_unsigned(1168, 12), 1328 => to_unsigned(383, 12), 1329 => to_unsigned(871, 12), 1330 => to_unsigned(617, 12), 1331 => to_unsigned(189, 12), 1332 => to_unsigned(3268, 12), 1333 => to_unsigned(3447, 12), 1334 => to_unsigned(3475, 12), 1335 => to_unsigned(2544, 12), 1336 => to_unsigned(2952, 12), 1337 => to_unsigned(498, 12), 1338 => to_unsigned(3024, 12), 1339 => to_unsigned(4065, 12), 1340 => to_unsigned(437, 12), 1341 => to_unsigned(441, 12), 1342 => to_unsigned(2704, 12), 1343 => to_unsigned(3616, 12), 1344 => to_unsigned(3426, 12), 1345 => to_unsigned(850, 12), 1346 => to_unsigned(3741, 12), 1347 => to_unsigned(1004, 12), 1348 => to_unsigned(3699, 12), 1349 => to_unsigned(279, 12), 1350 => to_unsigned(1526, 12), 1351 => to_unsigned(702, 12), 1352 => to_unsigned(2255, 12), 1353 => to_unsigned(3302, 12), 1354 => to_unsigned(2388, 12), 1355 => to_unsigned(798, 12), 1356 => to_unsigned(2798, 12), 1357 => to_unsigned(2490, 12), 1358 => to_unsigned(3670, 12), 1359 => to_unsigned(3066, 12), 1360 => to_unsigned(1756, 12), 1361 => to_unsigned(1735, 12), 1362 => to_unsigned(3813, 12), 1363 => to_unsigned(2482, 12), 1364 => to_unsigned(1141, 12), 1365 => to_unsigned(701, 12), 1366 => to_unsigned(813, 12), 1367 => to_unsigned(150, 12), 1368 => to_unsigned(2616, 12), 1369 => to_unsigned(1792, 12), 1370 => to_unsigned(512, 12), 1371 => to_unsigned(4008, 12), 1372 => to_unsigned(3752, 12), 1373 => to_unsigned(1877, 12), 1374 => to_unsigned(220, 12), 1375 => to_unsigned(3145, 12), 1376 => to_unsigned(2315, 12), 1377 => to_unsigned(825, 12), 1378 => to_unsigned(4062, 12), 1379 => to_unsigned(1360, 12), 1380 => to_unsigned(1472, 12), 1381 => to_unsigned(2718, 12), 1382 => to_unsigned(3245, 12), 1383 => to_unsigned(1353, 12), 1384 => to_unsigned(1474, 12), 1385 => to_unsigned(1806, 12), 1386 => to_unsigned(3212, 12), 1387 => to_unsigned(169, 12), 1388 => to_unsigned(1038, 12), 1389 => to_unsigned(3684, 12), 1390 => to_unsigned(2859, 12), 1391 => to_unsigned(870, 12), 1392 => to_unsigned(1225, 12), 1393 => to_unsigned(2187, 12), 1394 => to_unsigned(3454, 12), 1395 => to_unsigned(508, 12), 1396 => to_unsigned(858, 12), 1397 => to_unsigned(2515, 12), 1398 => to_unsigned(54, 12), 1399 => to_unsigned(303, 12), 1400 => to_unsigned(1579, 12), 1401 => to_unsigned(4042, 12), 1402 => to_unsigned(148, 12), 1403 => to_unsigned(2281, 12), 1404 => to_unsigned(3056, 12), 1405 => to_unsigned(52, 12), 1406 => to_unsigned(544, 12), 1407 => to_unsigned(3987, 12), 1408 => to_unsigned(2540, 12), 1409 => to_unsigned(1897, 12), 1410 => to_unsigned(1897, 12), 1411 => to_unsigned(1374, 12), 1412 => to_unsigned(2640, 12), 1413 => to_unsigned(2458, 12), 1414 => to_unsigned(1577, 12), 1415 => to_unsigned(4082, 12), 1416 => to_unsigned(1846, 12), 1417 => to_unsigned(3428, 12), 1418 => to_unsigned(1616, 12), 1419 => to_unsigned(2568, 12), 1420 => to_unsigned(3958, 12), 1421 => to_unsigned(1350, 12), 1422 => to_unsigned(2069, 12), 1423 => to_unsigned(3963, 12), 1424 => to_unsigned(727, 12), 1425 => to_unsigned(1636, 12), 1426 => to_unsigned(2204, 12), 1427 => to_unsigned(1840, 12), 1428 => to_unsigned(3401, 12), 1429 => to_unsigned(2979, 12), 1430 => to_unsigned(2430, 12), 1431 => to_unsigned(2679, 12), 1432 => to_unsigned(285, 12), 1433 => to_unsigned(122, 12), 1434 => to_unsigned(3758, 12), 1435 => to_unsigned(3502, 12), 1436 => to_unsigned(2863, 12), 1437 => to_unsigned(2419, 12), 1438 => to_unsigned(991, 12), 1439 => to_unsigned(1522, 12), 1440 => to_unsigned(712, 12), 1441 => to_unsigned(1329, 12), 1442 => to_unsigned(481, 12), 1443 => to_unsigned(2236, 12), 1444 => to_unsigned(2822, 12), 1445 => to_unsigned(2089, 12), 1446 => to_unsigned(4071, 12), 1447 => to_unsigned(227, 12), 1448 => to_unsigned(1762, 12), 1449 => to_unsigned(1750, 12), 1450 => to_unsigned(3950, 12), 1451 => to_unsigned(3998, 12), 1452 => to_unsigned(2816, 12), 1453 => to_unsigned(3367, 12), 1454 => to_unsigned(3193, 12), 1455 => to_unsigned(966, 12), 1456 => to_unsigned(3150, 12), 1457 => to_unsigned(1199, 12), 1458 => to_unsigned(727, 12), 1459 => to_unsigned(342, 12), 1460 => to_unsigned(1639, 12), 1461 => to_unsigned(2119, 12), 1462 => to_unsigned(3755, 12), 1463 => to_unsigned(1719, 12), 1464 => to_unsigned(2074, 12), 1465 => to_unsigned(1351, 12), 1466 => to_unsigned(632, 12), 1467 => to_unsigned(3247, 12), 1468 => to_unsigned(2054, 12), 1469 => to_unsigned(2749, 12), 1470 => to_unsigned(552, 12), 1471 => to_unsigned(798, 12), 1472 => to_unsigned(1764, 12), 1473 => to_unsigned(2695, 12), 1474 => to_unsigned(2187, 12), 1475 => to_unsigned(2996, 12), 1476 => to_unsigned(539, 12), 1477 => to_unsigned(18, 12), 1478 => to_unsigned(2897, 12), 1479 => to_unsigned(1418, 12), 1480 => to_unsigned(404, 12), 1481 => to_unsigned(2225, 12), 1482 => to_unsigned(705, 12), 1483 => to_unsigned(917, 12), 1484 => to_unsigned(2366, 12), 1485 => to_unsigned(3164, 12), 1486 => to_unsigned(3305, 12), 1487 => to_unsigned(1222, 12), 1488 => to_unsigned(3004, 12), 1489 => to_unsigned(3890, 12), 1490 => to_unsigned(1436, 12), 1491 => to_unsigned(3138, 12), 1492 => to_unsigned(3071, 12), 1493 => to_unsigned(842, 12), 1494 => to_unsigned(2665, 12), 1495 => to_unsigned(886, 12), 1496 => to_unsigned(2076, 12), 1497 => to_unsigned(1616, 12), 1498 => to_unsigned(164, 12), 1499 => to_unsigned(638, 12), 1500 => to_unsigned(2921, 12), 1501 => to_unsigned(3504, 12), 1502 => to_unsigned(375, 12), 1503 => to_unsigned(1373, 12), 1504 => to_unsigned(2706, 12), 1505 => to_unsigned(2689, 12), 1506 => to_unsigned(1134, 12), 1507 => to_unsigned(210, 12), 1508 => to_unsigned(3886, 12), 1509 => to_unsigned(826, 12), 1510 => to_unsigned(1449, 12), 1511 => to_unsigned(976, 12), 1512 => to_unsigned(339, 12), 1513 => to_unsigned(966, 12), 1514 => to_unsigned(1375, 12), 1515 => to_unsigned(10, 12), 1516 => to_unsigned(1054, 12), 1517 => to_unsigned(1524, 12), 1518 => to_unsigned(2015, 12), 1519 => to_unsigned(1251, 12), 1520 => to_unsigned(1942, 12), 1521 => to_unsigned(3210, 12), 1522 => to_unsigned(2923, 12), 1523 => to_unsigned(2189, 12), 1524 => to_unsigned(2784, 12), 1525 => to_unsigned(3726, 12), 1526 => to_unsigned(3384, 12), 1527 => to_unsigned(269, 12), 1528 => to_unsigned(2534, 12), 1529 => to_unsigned(3232, 12), 1530 => to_unsigned(2984, 12), 1531 => to_unsigned(3875, 12), 1532 => to_unsigned(4017, 12), 1533 => to_unsigned(2459, 12), 1534 => to_unsigned(2652, 12), 1535 => to_unsigned(3052, 12), 1536 => to_unsigned(2010, 12), 1537 => to_unsigned(2956, 12), 1538 => to_unsigned(223, 12), 1539 => to_unsigned(563, 12), 1540 => to_unsigned(33, 12), 1541 => to_unsigned(3384, 12), 1542 => to_unsigned(3886, 12), 1543 => to_unsigned(3397, 12), 1544 => to_unsigned(1005, 12), 1545 => to_unsigned(2683, 12), 1546 => to_unsigned(1339, 12), 1547 => to_unsigned(2772, 12), 1548 => to_unsigned(1168, 12), 1549 => to_unsigned(295, 12), 1550 => to_unsigned(1827, 12), 1551 => to_unsigned(2456, 12), 1552 => to_unsigned(3994, 12), 1553 => to_unsigned(2823, 12), 1554 => to_unsigned(164, 12), 1555 => to_unsigned(1637, 12), 1556 => to_unsigned(3864, 12), 1557 => to_unsigned(1490, 12), 1558 => to_unsigned(2205, 12), 1559 => to_unsigned(3226, 12), 1560 => to_unsigned(1879, 12), 1561 => to_unsigned(1966, 12), 1562 => to_unsigned(2091, 12), 1563 => to_unsigned(2198, 12), 1564 => to_unsigned(301, 12), 1565 => to_unsigned(2475, 12), 1566 => to_unsigned(3202, 12), 1567 => to_unsigned(1233, 12), 1568 => to_unsigned(61, 12), 1569 => to_unsigned(1472, 12), 1570 => to_unsigned(3424, 12), 1571 => to_unsigned(3627, 12), 1572 => to_unsigned(516, 12), 1573 => to_unsigned(422, 12), 1574 => to_unsigned(1692, 12), 1575 => to_unsigned(2106, 12), 1576 => to_unsigned(3618, 12), 1577 => to_unsigned(2205, 12), 1578 => to_unsigned(3880, 12), 1579 => to_unsigned(2540, 12), 1580 => to_unsigned(2425, 12), 1581 => to_unsigned(144, 12), 1582 => to_unsigned(158, 12), 1583 => to_unsigned(2303, 12), 1584 => to_unsigned(3080, 12), 1585 => to_unsigned(1836, 12), 1586 => to_unsigned(1378, 12), 1587 => to_unsigned(2881, 12), 1588 => to_unsigned(1175, 12), 1589 => to_unsigned(3707, 12), 1590 => to_unsigned(3933, 12), 1591 => to_unsigned(3924, 12), 1592 => to_unsigned(965, 12), 1593 => to_unsigned(2973, 12), 1594 => to_unsigned(169, 12), 1595 => to_unsigned(957, 12), 1596 => to_unsigned(3520, 12), 1597 => to_unsigned(1831, 12), 1598 => to_unsigned(593, 12), 1599 => to_unsigned(3095, 12), 1600 => to_unsigned(219, 12), 1601 => to_unsigned(3980, 12), 1602 => to_unsigned(2739, 12), 1603 => to_unsigned(3799, 12), 1604 => to_unsigned(2513, 12), 1605 => to_unsigned(2395, 12), 1606 => to_unsigned(987, 12), 1607 => to_unsigned(2924, 12), 1608 => to_unsigned(2246, 12), 1609 => to_unsigned(820, 12), 1610 => to_unsigned(4019, 12), 1611 => to_unsigned(202, 12), 1612 => to_unsigned(175, 12), 1613 => to_unsigned(2057, 12), 1614 => to_unsigned(609, 12), 1615 => to_unsigned(3121, 12), 1616 => to_unsigned(956, 12), 1617 => to_unsigned(3403, 12), 1618 => to_unsigned(3957, 12), 1619 => to_unsigned(1820, 12), 1620 => to_unsigned(2370, 12), 1621 => to_unsigned(2745, 12), 1622 => to_unsigned(885, 12), 1623 => to_unsigned(1158, 12), 1624 => to_unsigned(2977, 12), 1625 => to_unsigned(2187, 12), 1626 => to_unsigned(3379, 12), 1627 => to_unsigned(1499, 12), 1628 => to_unsigned(3479, 12), 1629 => to_unsigned(1743, 12), 1630 => to_unsigned(2208, 12), 1631 => to_unsigned(1220, 12), 1632 => to_unsigned(601, 12), 1633 => to_unsigned(2791, 12), 1634 => to_unsigned(3182, 12), 1635 => to_unsigned(3000, 12), 1636 => to_unsigned(1295, 12), 1637 => to_unsigned(472, 12), 1638 => to_unsigned(3234, 12), 1639 => to_unsigned(2722, 12), 1640 => to_unsigned(42, 12), 1641 => to_unsigned(3096, 12), 1642 => to_unsigned(752, 12), 1643 => to_unsigned(539, 12), 1644 => to_unsigned(1314, 12), 1645 => to_unsigned(1946, 12), 1646 => to_unsigned(2660, 12), 1647 => to_unsigned(3674, 12), 1648 => to_unsigned(2042, 12), 1649 => to_unsigned(1525, 12), 1650 => to_unsigned(3710, 12), 1651 => to_unsigned(493, 12), 1652 => to_unsigned(1451, 12), 1653 => to_unsigned(2085, 12), 1654 => to_unsigned(3192, 12), 1655 => to_unsigned(2786, 12), 1656 => to_unsigned(2660, 12), 1657 => to_unsigned(51, 12), 1658 => to_unsigned(1079, 12), 1659 => to_unsigned(1779, 12), 1660 => to_unsigned(3307, 12), 1661 => to_unsigned(972, 12), 1662 => to_unsigned(2344, 12), 1663 => to_unsigned(941, 12), 1664 => to_unsigned(275, 12), 1665 => to_unsigned(2708, 12), 1666 => to_unsigned(970, 12), 1667 => to_unsigned(791, 12), 1668 => to_unsigned(470, 12), 1669 => to_unsigned(2998, 12), 1670 => to_unsigned(450, 12), 1671 => to_unsigned(1339, 12), 1672 => to_unsigned(3199, 12), 1673 => to_unsigned(1568, 12), 1674 => to_unsigned(1715, 12), 1675 => to_unsigned(946, 12), 1676 => to_unsigned(992, 12), 1677 => to_unsigned(3496, 12), 1678 => to_unsigned(2410, 12), 1679 => to_unsigned(3442, 12), 1680 => to_unsigned(888, 12), 1681 => to_unsigned(1282, 12), 1682 => to_unsigned(82, 12), 1683 => to_unsigned(1341, 12), 1684 => to_unsigned(3156, 12), 1685 => to_unsigned(1327, 12), 1686 => to_unsigned(250, 12), 1687 => to_unsigned(718, 12), 1688 => to_unsigned(2775, 12), 1689 => to_unsigned(1230, 12), 1690 => to_unsigned(3061, 12), 1691 => to_unsigned(823, 12), 1692 => to_unsigned(1331, 12), 1693 => to_unsigned(821, 12), 1694 => to_unsigned(3354, 12), 1695 => to_unsigned(2879, 12), 1696 => to_unsigned(967, 12), 1697 => to_unsigned(3391, 12), 1698 => to_unsigned(2450, 12), 1699 => to_unsigned(2281, 12), 1700 => to_unsigned(1343, 12), 1701 => to_unsigned(150, 12), 1702 => to_unsigned(3868, 12), 1703 => to_unsigned(2491, 12), 1704 => to_unsigned(734, 12), 1705 => to_unsigned(1540, 12), 1706 => to_unsigned(3439, 12), 1707 => to_unsigned(632, 12), 1708 => to_unsigned(3051, 12), 1709 => to_unsigned(319, 12), 1710 => to_unsigned(364, 12), 1711 => to_unsigned(1695, 12), 1712 => to_unsigned(1129, 12), 1713 => to_unsigned(660, 12), 1714 => to_unsigned(1713, 12), 1715 => to_unsigned(1318, 12), 1716 => to_unsigned(731, 12), 1717 => to_unsigned(3270, 12), 1718 => to_unsigned(105, 12), 1719 => to_unsigned(1022, 12), 1720 => to_unsigned(1542, 12), 1721 => to_unsigned(1442, 12), 1722 => to_unsigned(2252, 12), 1723 => to_unsigned(4043, 12), 1724 => to_unsigned(2913, 12), 1725 => to_unsigned(2358, 12), 1726 => to_unsigned(2729, 12), 1727 => to_unsigned(324, 12), 1728 => to_unsigned(1841, 12), 1729 => to_unsigned(791, 12), 1730 => to_unsigned(1172, 12), 1731 => to_unsigned(897, 12), 1732 => to_unsigned(2284, 12), 1733 => to_unsigned(2702, 12), 1734 => to_unsigned(1022, 12), 1735 => to_unsigned(694, 12), 1736 => to_unsigned(136, 12), 1737 => to_unsigned(88, 12), 1738 => to_unsigned(252, 12), 1739 => to_unsigned(309, 12), 1740 => to_unsigned(2512, 12), 1741 => to_unsigned(3560, 12), 1742 => to_unsigned(4066, 12), 1743 => to_unsigned(746, 12), 1744 => to_unsigned(537, 12), 1745 => to_unsigned(2795, 12), 1746 => to_unsigned(699, 12), 1747 => to_unsigned(1334, 12), 1748 => to_unsigned(2548, 12), 1749 => to_unsigned(535, 12), 1750 => to_unsigned(3072, 12), 1751 => to_unsigned(2682, 12), 1752 => to_unsigned(1204, 12), 1753 => to_unsigned(3162, 12), 1754 => to_unsigned(8, 12), 1755 => to_unsigned(413, 12), 1756 => to_unsigned(2842, 12), 1757 => to_unsigned(925, 12), 1758 => to_unsigned(2600, 12), 1759 => to_unsigned(2319, 12), 1760 => to_unsigned(2305, 12), 1761 => to_unsigned(3262, 12), 1762 => to_unsigned(2633, 12), 1763 => to_unsigned(1049, 12), 1764 => to_unsigned(2427, 12), 1765 => to_unsigned(2092, 12), 1766 => to_unsigned(3355, 12), 1767 => to_unsigned(1102, 12), 1768 => to_unsigned(2929, 12), 1769 => to_unsigned(2591, 12), 1770 => to_unsigned(1265, 12), 1771 => to_unsigned(1952, 12), 1772 => to_unsigned(2815, 12), 1773 => to_unsigned(967, 12), 1774 => to_unsigned(2087, 12), 1775 => to_unsigned(2683, 12), 1776 => to_unsigned(10, 12), 1777 => to_unsigned(3822, 12), 1778 => to_unsigned(4009, 12), 1779 => to_unsigned(3201, 12), 1780 => to_unsigned(542, 12), 1781 => to_unsigned(3999, 12), 1782 => to_unsigned(3114, 12), 1783 => to_unsigned(2995, 12), 1784 => to_unsigned(375, 12), 1785 => to_unsigned(1484, 12), 1786 => to_unsigned(709, 12), 1787 => to_unsigned(3744, 12), 1788 => to_unsigned(1505, 12), 1789 => to_unsigned(2319, 12), 1790 => to_unsigned(2862, 12), 1791 => to_unsigned(1571, 12), 1792 => to_unsigned(1337, 12), 1793 => to_unsigned(2548, 12), 1794 => to_unsigned(2278, 12), 1795 => to_unsigned(862, 12), 1796 => to_unsigned(581, 12), 1797 => to_unsigned(857, 12), 1798 => to_unsigned(677, 12), 1799 => to_unsigned(1815, 12), 1800 => to_unsigned(4021, 12), 1801 => to_unsigned(3389, 12), 1802 => to_unsigned(3992, 12), 1803 => to_unsigned(179, 12), 1804 => to_unsigned(662, 12), 1805 => to_unsigned(2550, 12), 1806 => to_unsigned(2886, 12), 1807 => to_unsigned(916, 12), 1808 => to_unsigned(209, 12), 1809 => to_unsigned(2238, 12), 1810 => to_unsigned(1112, 12), 1811 => to_unsigned(3554, 12), 1812 => to_unsigned(65, 12), 1813 => to_unsigned(1063, 12), 1814 => to_unsigned(171, 12), 1815 => to_unsigned(2199, 12), 1816 => to_unsigned(1819, 12), 1817 => to_unsigned(928, 12), 1818 => to_unsigned(4057, 12), 1819 => to_unsigned(2368, 12), 1820 => to_unsigned(2547, 12), 1821 => to_unsigned(3608, 12), 1822 => to_unsigned(1893, 12), 1823 => to_unsigned(3415, 12), 1824 => to_unsigned(3313, 12), 1825 => to_unsigned(849, 12), 1826 => to_unsigned(1278, 12), 1827 => to_unsigned(2909, 12), 1828 => to_unsigned(1460, 12), 1829 => to_unsigned(1795, 12), 1830 => to_unsigned(3829, 12), 1831 => to_unsigned(3058, 12), 1832 => to_unsigned(1996, 12), 1833 => to_unsigned(483, 12), 1834 => to_unsigned(3747, 12), 1835 => to_unsigned(3882, 12), 1836 => to_unsigned(1622, 12), 1837 => to_unsigned(1148, 12), 1838 => to_unsigned(222, 12), 1839 => to_unsigned(1606, 12), 1840 => to_unsigned(2622, 12), 1841 => to_unsigned(2105, 12), 1842 => to_unsigned(173, 12), 1843 => to_unsigned(200, 12), 1844 => to_unsigned(2489, 12), 1845 => to_unsigned(2287, 12), 1846 => to_unsigned(2192, 12), 1847 => to_unsigned(198, 12), 1848 => to_unsigned(3210, 12), 1849 => to_unsigned(1356, 12), 1850 => to_unsigned(2042, 12), 1851 => to_unsigned(3655, 12), 1852 => to_unsigned(4040, 12), 1853 => to_unsigned(445, 12), 1854 => to_unsigned(1117, 12), 1855 => to_unsigned(4038, 12), 1856 => to_unsigned(1799, 12), 1857 => to_unsigned(1938, 12), 1858 => to_unsigned(1856, 12), 1859 => to_unsigned(61, 12), 1860 => to_unsigned(2298, 12), 1861 => to_unsigned(1323, 12), 1862 => to_unsigned(143, 12), 1863 => to_unsigned(3818, 12), 1864 => to_unsigned(3546, 12), 1865 => to_unsigned(1716, 12), 1866 => to_unsigned(2278, 12), 1867 => to_unsigned(3464, 12), 1868 => to_unsigned(274, 12), 1869 => to_unsigned(1004, 12), 1870 => to_unsigned(594, 12), 1871 => to_unsigned(334, 12), 1872 => to_unsigned(3276, 12), 1873 => to_unsigned(1116, 12), 1874 => to_unsigned(425, 12), 1875 => to_unsigned(1744, 12), 1876 => to_unsigned(1206, 12), 1877 => to_unsigned(3326, 12), 1878 => to_unsigned(1637, 12), 1879 => to_unsigned(2274, 12), 1880 => to_unsigned(1531, 12), 1881 => to_unsigned(1709, 12), 1882 => to_unsigned(2743, 12), 1883 => to_unsigned(2395, 12), 1884 => to_unsigned(3480, 12), 1885 => to_unsigned(320, 12), 1886 => to_unsigned(3830, 12), 1887 => to_unsigned(9, 12), 1888 => to_unsigned(2636, 12), 1889 => to_unsigned(3426, 12), 1890 => to_unsigned(3925, 12), 1891 => to_unsigned(3086, 12), 1892 => to_unsigned(3972, 12), 1893 => to_unsigned(393, 12), 1894 => to_unsigned(1429, 12), 1895 => to_unsigned(2707, 12), 1896 => to_unsigned(855, 12), 1897 => to_unsigned(1307, 12), 1898 => to_unsigned(3710, 12), 1899 => to_unsigned(4083, 12), 1900 => to_unsigned(593, 12), 1901 => to_unsigned(1162, 12), 1902 => to_unsigned(798, 12), 1903 => to_unsigned(427, 12), 1904 => to_unsigned(928, 12), 1905 => to_unsigned(1287, 12), 1906 => to_unsigned(1060, 12), 1907 => to_unsigned(3440, 12), 1908 => to_unsigned(1467, 12), 1909 => to_unsigned(183, 12), 1910 => to_unsigned(3662, 12), 1911 => to_unsigned(3046, 12), 1912 => to_unsigned(640, 12), 1913 => to_unsigned(387, 12), 1914 => to_unsigned(2523, 12), 1915 => to_unsigned(1707, 12), 1916 => to_unsigned(26, 12), 1917 => to_unsigned(3869, 12), 1918 => to_unsigned(839, 12), 1919 => to_unsigned(3262, 12), 1920 => to_unsigned(1880, 12), 1921 => to_unsigned(1584, 12), 1922 => to_unsigned(853, 12), 1923 => to_unsigned(4000, 12), 1924 => to_unsigned(3975, 12), 1925 => to_unsigned(1502, 12), 1926 => to_unsigned(199, 12), 1927 => to_unsigned(2885, 12), 1928 => to_unsigned(2512, 12), 1929 => to_unsigned(1544, 12), 1930 => to_unsigned(4024, 12), 1931 => to_unsigned(2045, 12), 1932 => to_unsigned(231, 12), 1933 => to_unsigned(3544, 12), 1934 => to_unsigned(3515, 12), 1935 => to_unsigned(2123, 12), 1936 => to_unsigned(2170, 12), 1937 => to_unsigned(982, 12), 1938 => to_unsigned(2850, 12), 1939 => to_unsigned(3384, 12), 1940 => to_unsigned(873, 12), 1941 => to_unsigned(2723, 12), 1942 => to_unsigned(2662, 12), 1943 => to_unsigned(2474, 12), 1944 => to_unsigned(3301, 12), 1945 => to_unsigned(3973, 12), 1946 => to_unsigned(3119, 12), 1947 => to_unsigned(2010, 12), 1948 => to_unsigned(2738, 12), 1949 => to_unsigned(2797, 12), 1950 => to_unsigned(2179, 12), 1951 => to_unsigned(409, 12), 1952 => to_unsigned(2795, 12), 1953 => to_unsigned(2241, 12), 1954 => to_unsigned(1958, 12), 1955 => to_unsigned(242, 12), 1956 => to_unsigned(1963, 12), 1957 => to_unsigned(3671, 12), 1958 => to_unsigned(1174, 12), 1959 => to_unsigned(3693, 12), 1960 => to_unsigned(3741, 12), 1961 => to_unsigned(1315, 12), 1962 => to_unsigned(3331, 12), 1963 => to_unsigned(979, 12), 1964 => to_unsigned(3687, 12), 1965 => to_unsigned(1725, 12), 1966 => to_unsigned(1474, 12), 1967 => to_unsigned(276, 12), 1968 => to_unsigned(19, 12), 1969 => to_unsigned(1008, 12), 1970 => to_unsigned(2885, 12), 1971 => to_unsigned(2864, 12), 1972 => to_unsigned(3964, 12), 1973 => to_unsigned(3589, 12), 1974 => to_unsigned(559, 12), 1975 => to_unsigned(1234, 12), 1976 => to_unsigned(420, 12), 1977 => to_unsigned(1499, 12), 1978 => to_unsigned(3146, 12), 1979 => to_unsigned(2369, 12), 1980 => to_unsigned(2687, 12), 1981 => to_unsigned(3878, 12), 1982 => to_unsigned(129, 12), 1983 => to_unsigned(2763, 12), 1984 => to_unsigned(3759, 12), 1985 => to_unsigned(438, 12), 1986 => to_unsigned(79, 12), 1987 => to_unsigned(1203, 12), 1988 => to_unsigned(3113, 12), 1989 => to_unsigned(1419, 12), 1990 => to_unsigned(1799, 12), 1991 => to_unsigned(4031, 12), 1992 => to_unsigned(3195, 12), 1993 => to_unsigned(2019, 12), 1994 => to_unsigned(918, 12), 1995 => to_unsigned(1533, 12), 1996 => to_unsigned(3366, 12), 1997 => to_unsigned(142, 12), 1998 => to_unsigned(718, 12), 1999 => to_unsigned(3024, 12), 2000 => to_unsigned(2543, 12), 2001 => to_unsigned(3616, 12), 2002 => to_unsigned(361, 12), 2003 => to_unsigned(886, 12), 2004 => to_unsigned(2537, 12), 2005 => to_unsigned(362, 12), 2006 => to_unsigned(651, 12), 2007 => to_unsigned(625, 12), 2008 => to_unsigned(4087, 12), 2009 => to_unsigned(2849, 12), 2010 => to_unsigned(923, 12), 2011 => to_unsigned(2276, 12), 2012 => to_unsigned(1910, 12), 2013 => to_unsigned(1758, 12), 2014 => to_unsigned(52, 12), 2015 => to_unsigned(3169, 12), 2016 => to_unsigned(3519, 12), 2017 => to_unsigned(3990, 12), 2018 => to_unsigned(2422, 12), 2019 => to_unsigned(2688, 12), 2020 => to_unsigned(416, 12), 2021 => to_unsigned(1184, 12), 2022 => to_unsigned(3615, 12), 2023 => to_unsigned(191, 12), 2024 => to_unsigned(533, 12), 2025 => to_unsigned(738, 12), 2026 => to_unsigned(2534, 12), 2027 => to_unsigned(441, 12), 2028 => to_unsigned(1547, 12), 2029 => to_unsigned(3036, 12), 2030 => to_unsigned(626, 12), 2031 => to_unsigned(3797, 12), 2032 => to_unsigned(3118, 12), 2033 => to_unsigned(166, 12), 2034 => to_unsigned(2838, 12), 2035 => to_unsigned(2447, 12), 2036 => to_unsigned(1754, 12), 2037 => to_unsigned(3883, 12), 2038 => to_unsigned(2302, 12), 2039 => to_unsigned(1188, 12), 2040 => to_unsigned(60, 12), 2041 => to_unsigned(2420, 12), 2042 => to_unsigned(2501, 12), 2043 => to_unsigned(677, 12), 2044 => to_unsigned(579, 12), 2045 => to_unsigned(3542, 12), 2046 => to_unsigned(3682, 12), 2047 => to_unsigned(2487, 12))
        )
    );

    type averages_t is array(0 to 2) of vnir_row_t;
    constant averages : averages_t := (
        0 => (0 => to_unsigned(2627, 12), 1 => to_unsigned(1494, 12), 2 => to_unsigned(1808, 12), 3 => to_unsigned(2243, 12), 4 => to_unsigned(1698, 12), 5 => to_unsigned(2068, 12), 6 => to_unsigned(2295, 12), 7 => to_unsigned(1841, 12), 8 => to_unsigned(1596, 12), 9 => to_unsigned(2170, 12), 10 => to_unsigned(1996, 12), 11 => to_unsigned(2465, 12), 12 => to_unsigned(2247, 12), 13 => to_unsigned(2454, 12), 14 => to_unsigned(2362, 12), 15 => to_unsigned(1718, 12), 16 => to_unsigned(1196, 12), 17 => to_unsigned(1932, 12), 18 => to_unsigned(2288, 12), 19 => to_unsigned(1443, 12), 20 => to_unsigned(2273, 12), 21 => to_unsigned(2790, 12), 22 => to_unsigned(1954, 12), 23 => to_unsigned(2041, 12), 24 => to_unsigned(2662, 12), 25 => to_unsigned(2126, 12), 26 => to_unsigned(2011, 12), 27 => to_unsigned(1933, 12), 28 => to_unsigned(1402, 12), 29 => to_unsigned(2082, 12), 30 => to_unsigned(2129, 12), 31 => to_unsigned(1875, 12), 32 => to_unsigned(1550, 12), 33 => to_unsigned(2127, 12), 34 => to_unsigned(2086, 12), 35 => to_unsigned(1903, 12), 36 => to_unsigned(1677, 12), 37 => to_unsigned(1793, 12), 38 => to_unsigned(1911, 12), 39 => to_unsigned(2231, 12), 40 => to_unsigned(1374, 12), 41 => to_unsigned(2256, 12), 42 => to_unsigned(1933, 12), 43 => to_unsigned(1663, 12), 44 => to_unsigned(1676, 12), 45 => to_unsigned(1799, 12), 46 => to_unsigned(1544, 12), 47 => to_unsigned(1712, 12), 48 => to_unsigned(1834, 12), 49 => to_unsigned(1474, 12), 50 => to_unsigned(1690, 12), 51 => to_unsigned(2256, 12), 52 => to_unsigned(2639, 12), 53 => to_unsigned(2044, 12), 54 => to_unsigned(2199, 12), 55 => to_unsigned(1750, 12), 56 => to_unsigned(1807, 12), 57 => to_unsigned(1541, 12), 58 => to_unsigned(2040, 12), 59 => to_unsigned(2622, 12), 60 => to_unsigned(2275, 12), 61 => to_unsigned(2893, 12), 62 => to_unsigned(2483, 12), 63 => to_unsigned(1633, 12), 64 => to_unsigned(1669, 12), 65 => to_unsigned(2163, 12), 66 => to_unsigned(1408, 12), 67 => to_unsigned(1882, 12), 68 => to_unsigned(1784, 12), 69 => to_unsigned(1725, 12), 70 => to_unsigned(1856, 12), 71 => to_unsigned(2163, 12), 72 => to_unsigned(2538, 12), 73 => to_unsigned(2312, 12), 74 => to_unsigned(2359, 12), 75 => to_unsigned(1758, 12), 76 => to_unsigned(2413, 12), 77 => to_unsigned(1850, 12), 78 => to_unsigned(1507, 12), 79 => to_unsigned(2742, 12), 80 => to_unsigned(2515, 12), 81 => to_unsigned(1991, 12), 82 => to_unsigned(2110, 12), 83 => to_unsigned(1641, 12), 84 => to_unsigned(2093, 12), 85 => to_unsigned(2306, 12), 86 => to_unsigned(2296, 12), 87 => to_unsigned(2041, 12), 88 => to_unsigned(2683, 12), 89 => to_unsigned(2116, 12), 90 => to_unsigned(1691, 12), 91 => to_unsigned(2057, 12), 92 => to_unsigned(1730, 12), 93 => to_unsigned(1929, 12), 94 => to_unsigned(2142, 12), 95 => to_unsigned(1723, 12), 96 => to_unsigned(2150, 12), 97 => to_unsigned(2057, 12), 98 => to_unsigned(2208, 12), 99 => to_unsigned(2378, 12), 100 => to_unsigned(2198, 12), 101 => to_unsigned(1801, 12), 102 => to_unsigned(2297, 12), 103 => to_unsigned(2167, 12), 104 => to_unsigned(1970, 12), 105 => to_unsigned(2199, 12), 106 => to_unsigned(2486, 12), 107 => to_unsigned(2229, 12), 108 => to_unsigned(2478, 12), 109 => to_unsigned(2014, 12), 110 => to_unsigned(1315, 12), 111 => to_unsigned(1053, 12), 112 => to_unsigned(2162, 12), 113 => to_unsigned(1920, 12), 114 => to_unsigned(2131, 12), 115 => to_unsigned(2409, 12), 116 => to_unsigned(2116, 12), 117 => to_unsigned(2038, 12), 118 => to_unsigned(2427, 12), 119 => to_unsigned(2038, 12), 120 => to_unsigned(2818, 12), 121 => to_unsigned(2321, 12), 122 => to_unsigned(1641, 12), 123 => to_unsigned(1276, 12), 124 => to_unsigned(1870, 12), 125 => to_unsigned(1926, 12), 126 => to_unsigned(1886, 12), 127 => to_unsigned(2530, 12), 128 => to_unsigned(2049, 12), 129 => to_unsigned(2040, 12), 130 => to_unsigned(2128, 12), 131 => to_unsigned(2220, 12), 132 => to_unsigned(1940, 12), 133 => to_unsigned(2369, 12), 134 => to_unsigned(2097, 12), 135 => to_unsigned(1550, 12), 136 => to_unsigned(2358, 12), 137 => to_unsigned(2015, 12), 138 => to_unsigned(2457, 12), 139 => to_unsigned(2222, 12), 140 => to_unsigned(2550, 12), 141 => to_unsigned(1611, 12), 142 => to_unsigned(1960, 12), 143 => to_unsigned(2579, 12), 144 => to_unsigned(1921, 12), 145 => to_unsigned(2036, 12), 146 => to_unsigned(1673, 12), 147 => to_unsigned(2618, 12), 148 => to_unsigned(1814, 12), 149 => to_unsigned(2425, 12), 150 => to_unsigned(1848, 12), 151 => to_unsigned(1717, 12), 152 => to_unsigned(2037, 12), 153 => to_unsigned(1963, 12), 154 => to_unsigned(2454, 12), 155 => to_unsigned(1973, 12), 156 => to_unsigned(1958, 12), 157 => to_unsigned(2350, 12), 158 => to_unsigned(2018, 12), 159 => to_unsigned(2521, 12), 160 => to_unsigned(1663, 12), 161 => to_unsigned(2410, 12), 162 => to_unsigned(1983, 12), 163 => to_unsigned(1740, 12), 164 => to_unsigned(2133, 12), 165 => to_unsigned(1733, 12), 166 => to_unsigned(2279, 12), 167 => to_unsigned(1656, 12), 168 => to_unsigned(2839, 12), 169 => to_unsigned(1613, 12), 170 => to_unsigned(2022, 12), 171 => to_unsigned(1911, 12), 172 => to_unsigned(1519, 12), 173 => to_unsigned(2115, 12), 174 => to_unsigned(2596, 12), 175 => to_unsigned(1188, 12), 176 => to_unsigned(1231, 12), 177 => to_unsigned(1600, 12), 178 => to_unsigned(2548, 12), 179 => to_unsigned(2103, 12), 180 => to_unsigned(1557, 12), 181 => to_unsigned(2406, 12), 182 => to_unsigned(2518, 12), 183 => to_unsigned(2022, 12), 184 => to_unsigned(1913, 12), 185 => to_unsigned(2567, 12), 186 => to_unsigned(2488, 12), 187 => to_unsigned(2348, 12), 188 => to_unsigned(1225, 12), 189 => to_unsigned(2043, 12), 190 => to_unsigned(1648, 12), 191 => to_unsigned(1565, 12), 192 => to_unsigned(1814, 12), 193 => to_unsigned(2166, 12), 194 => to_unsigned(2065, 12), 195 => to_unsigned(2123, 12), 196 => to_unsigned(2221, 12), 197 => to_unsigned(2475, 12), 198 => to_unsigned(1498, 12), 199 => to_unsigned(1330, 12), 200 => to_unsigned(1333, 12), 201 => to_unsigned(1877, 12), 202 => to_unsigned(1878, 12), 203 => to_unsigned(1943, 12), 204 => to_unsigned(2455, 12), 205 => to_unsigned(1936, 12), 206 => to_unsigned(1695, 12), 207 => to_unsigned(2688, 12), 208 => to_unsigned(2505, 12), 209 => to_unsigned(2246, 12), 210 => to_unsigned(1934, 12), 211 => to_unsigned(2211, 12), 212 => to_unsigned(2202, 12), 213 => to_unsigned(1465, 12), 214 => to_unsigned(2120, 12), 215 => to_unsigned(2251, 12), 216 => to_unsigned(1844, 12), 217 => to_unsigned(2486, 12), 218 => to_unsigned(1656, 12), 219 => to_unsigned(2329, 12), 220 => to_unsigned(3148, 12), 221 => to_unsigned(2202, 12), 222 => to_unsigned(1758, 12), 223 => to_unsigned(2200, 12), 224 => to_unsigned(1882, 12), 225 => to_unsigned(2427, 12), 226 => to_unsigned(1295, 12), 227 => to_unsigned(2312, 12), 228 => to_unsigned(1965, 12), 229 => to_unsigned(2105, 12), 230 => to_unsigned(2508, 12), 231 => to_unsigned(1629, 12), 232 => to_unsigned(1723, 12), 233 => to_unsigned(2349, 12), 234 => to_unsigned(2303, 12), 235 => to_unsigned(1680, 12), 236 => to_unsigned(2442, 12), 237 => to_unsigned(1911, 12), 238 => to_unsigned(1869, 12), 239 => to_unsigned(2205, 12), 240 => to_unsigned(2324, 12), 241 => to_unsigned(2365, 12), 242 => to_unsigned(1774, 12), 243 => to_unsigned(1129, 12), 244 => to_unsigned(2058, 12), 245 => to_unsigned(1316, 12), 246 => to_unsigned(1718, 12), 247 => to_unsigned(1875, 12), 248 => to_unsigned(1458, 12), 249 => to_unsigned(2440, 12), 250 => to_unsigned(1975, 12), 251 => to_unsigned(1945, 12), 252 => to_unsigned(2557, 12), 253 => to_unsigned(1370, 12), 254 => to_unsigned(1792, 12), 255 => to_unsigned(1328, 12), 256 => to_unsigned(2337, 12), 257 => to_unsigned(2016, 12), 258 => to_unsigned(1580, 12), 259 => to_unsigned(1238, 12), 260 => to_unsigned(1883, 12), 261 => to_unsigned(1445, 12), 262 => to_unsigned(1785, 12), 263 => to_unsigned(2223, 12), 264 => to_unsigned(2449, 12), 265 => to_unsigned(2448, 12), 266 => to_unsigned(1548, 12), 267 => to_unsigned(1882, 12), 268 => to_unsigned(1871, 12), 269 => to_unsigned(1908, 12), 270 => to_unsigned(1821, 12), 271 => to_unsigned(1988, 12), 272 => to_unsigned(1799, 12), 273 => to_unsigned(2312, 12), 274 => to_unsigned(2730, 12), 275 => to_unsigned(2453, 12), 276 => to_unsigned(2496, 12), 277 => to_unsigned(1610, 12), 278 => to_unsigned(1917, 12), 279 => to_unsigned(2858, 12), 280 => to_unsigned(1842, 12), 281 => to_unsigned(1766, 12), 282 => to_unsigned(2041, 12), 283 => to_unsigned(2247, 12), 284 => to_unsigned(2404, 12), 285 => to_unsigned(1996, 12), 286 => to_unsigned(1595, 12), 287 => to_unsigned(1200, 12), 288 => to_unsigned(1765, 12), 289 => to_unsigned(1870, 12), 290 => to_unsigned(1922, 12), 291 => to_unsigned(2323, 12), 292 => to_unsigned(2057, 12), 293 => to_unsigned(1816, 12), 294 => to_unsigned(2659, 12), 295 => to_unsigned(2533, 12), 296 => to_unsigned(1614, 12), 297 => to_unsigned(1837, 12), 298 => to_unsigned(2591, 12), 299 => to_unsigned(1614, 12), 300 => to_unsigned(1761, 12), 301 => to_unsigned(2517, 12), 302 => to_unsigned(2239, 12), 303 => to_unsigned(2561, 12), 304 => to_unsigned(2244, 12), 305 => to_unsigned(1454, 12), 306 => to_unsigned(2204, 12), 307 => to_unsigned(1906, 12), 308 => to_unsigned(2046, 12), 309 => to_unsigned(1733, 12), 310 => to_unsigned(1983, 12), 311 => to_unsigned(2111, 12), 312 => to_unsigned(1556, 12), 313 => to_unsigned(2550, 12), 314 => to_unsigned(1999, 12), 315 => to_unsigned(2413, 12), 316 => to_unsigned(1957, 12), 317 => to_unsigned(2795, 12), 318 => to_unsigned(2663, 12), 319 => to_unsigned(1879, 12), 320 => to_unsigned(1997, 12), 321 => to_unsigned(2099, 12), 322 => to_unsigned(1814, 12), 323 => to_unsigned(1965, 12), 324 => to_unsigned(2176, 12), 325 => to_unsigned(1905, 12), 326 => to_unsigned(2172, 12), 327 => to_unsigned(2050, 12), 328 => to_unsigned(2166, 12), 329 => to_unsigned(2534, 12), 330 => to_unsigned(2063, 12), 331 => to_unsigned(2341, 12), 332 => to_unsigned(1510, 12), 333 => to_unsigned(2083, 12), 334 => to_unsigned(1558, 12), 335 => to_unsigned(2103, 12), 336 => to_unsigned(2479, 12), 337 => to_unsigned(2299, 12), 338 => to_unsigned(2480, 12), 339 => to_unsigned(2645, 12), 340 => to_unsigned(1230, 12), 341 => to_unsigned(2823, 12), 342 => to_unsigned(1948, 12), 343 => to_unsigned(1487, 12), 344 => to_unsigned(2335, 12), 345 => to_unsigned(2172, 12), 346 => to_unsigned(1465, 12), 347 => to_unsigned(2542, 12), 348 => to_unsigned(1990, 12), 349 => to_unsigned(2332, 12), 350 => to_unsigned(1639, 12), 351 => to_unsigned(1369, 12), 352 => to_unsigned(1480, 12), 353 => to_unsigned(2330, 12), 354 => to_unsigned(1834, 12), 355 => to_unsigned(2556, 12), 356 => to_unsigned(1323, 12), 357 => to_unsigned(1708, 12), 358 => to_unsigned(2056, 12), 359 => to_unsigned(1828, 12), 360 => to_unsigned(2523, 12), 361 => to_unsigned(2398, 12), 362 => to_unsigned(1867, 12), 363 => to_unsigned(2229, 12), 364 => to_unsigned(1670, 12), 365 => to_unsigned(2449, 12), 366 => to_unsigned(1690, 12), 367 => to_unsigned(1072, 12), 368 => to_unsigned(1552, 12), 369 => to_unsigned(1532, 12), 370 => to_unsigned(2397, 12), 371 => to_unsigned(1598, 12), 372 => to_unsigned(2051, 12), 373 => to_unsigned(2122, 12), 374 => to_unsigned(2039, 12), 375 => to_unsigned(1607, 12), 376 => to_unsigned(2080, 12), 377 => to_unsigned(2132, 12), 378 => to_unsigned(2023, 12), 379 => to_unsigned(1855, 12), 380 => to_unsigned(1592, 12), 381 => to_unsigned(2100, 12), 382 => to_unsigned(1764, 12), 383 => to_unsigned(2186, 12), 384 => to_unsigned(2073, 12), 385 => to_unsigned(1667, 12), 386 => to_unsigned(1941, 12), 387 => to_unsigned(2027, 12), 388 => to_unsigned(2576, 12), 389 => to_unsigned(2761, 12), 390 => to_unsigned(2530, 12), 391 => to_unsigned(1916, 12), 392 => to_unsigned(2126, 12), 393 => to_unsigned(2775, 12), 394 => to_unsigned(1585, 12), 395 => to_unsigned(2428, 12), 396 => to_unsigned(2403, 12), 397 => to_unsigned(2188, 12), 398 => to_unsigned(2582, 12), 399 => to_unsigned(2349, 12), 400 => to_unsigned(2009, 12), 401 => to_unsigned(2639, 12), 402 => to_unsigned(1796, 12), 403 => to_unsigned(1787, 12), 404 => to_unsigned(2605, 12), 405 => to_unsigned(2290, 12), 406 => to_unsigned(1710, 12), 407 => to_unsigned(2136, 12), 408 => to_unsigned(2061, 12), 409 => to_unsigned(2350, 12), 410 => to_unsigned(1545, 12), 411 => to_unsigned(1432, 12), 412 => to_unsigned(2452, 12), 413 => to_unsigned(1849, 12), 414 => to_unsigned(1566, 12), 415 => to_unsigned(2104, 12), 416 => to_unsigned(1412, 12), 417 => to_unsigned(2352, 12), 418 => to_unsigned(2367, 12), 419 => to_unsigned(1412, 12), 420 => to_unsigned(2076, 12), 421 => to_unsigned(2038, 12), 422 => to_unsigned(2555, 12), 423 => to_unsigned(2188, 12), 424 => to_unsigned(2475, 12), 425 => to_unsigned(1238, 12), 426 => to_unsigned(2181, 12), 427 => to_unsigned(2173, 12), 428 => to_unsigned(1487, 12), 429 => to_unsigned(2502, 12), 430 => to_unsigned(1844, 12), 431 => to_unsigned(2174, 12), 432 => to_unsigned(1639, 12), 433 => to_unsigned(1944, 12), 434 => to_unsigned(908, 12), 435 => to_unsigned(1766, 12), 436 => to_unsigned(2062, 12), 437 => to_unsigned(2034, 12), 438 => to_unsigned(1698, 12), 439 => to_unsigned(2230, 12), 440 => to_unsigned(1622, 12), 441 => to_unsigned(2365, 12), 442 => to_unsigned(1966, 12), 443 => to_unsigned(2125, 12), 444 => to_unsigned(2265, 12), 445 => to_unsigned(1847, 12), 446 => to_unsigned(2711, 12), 447 => to_unsigned(1873, 12), 448 => to_unsigned(2594, 12), 449 => to_unsigned(1710, 12), 450 => to_unsigned(2534, 12), 451 => to_unsigned(2581, 12), 452 => to_unsigned(1617, 12), 453 => to_unsigned(1561, 12), 454 => to_unsigned(1603, 12), 455 => to_unsigned(1719, 12), 456 => to_unsigned(2500, 12), 457 => to_unsigned(1917, 12), 458 => to_unsigned(2075, 12), 459 => to_unsigned(2622, 12), 460 => to_unsigned(1729, 12), 461 => to_unsigned(1966, 12), 462 => to_unsigned(1714, 12), 463 => to_unsigned(2229, 12), 464 => to_unsigned(2618, 12), 465 => to_unsigned(2045, 12), 466 => to_unsigned(1707, 12), 467 => to_unsigned(2490, 12), 468 => to_unsigned(1703, 12), 469 => to_unsigned(2173, 12), 470 => to_unsigned(2090, 12), 471 => to_unsigned(1792, 12), 472 => to_unsigned(2186, 12), 473 => to_unsigned(1837, 12), 474 => to_unsigned(1662, 12), 475 => to_unsigned(1861, 12), 476 => to_unsigned(1606, 12), 477 => to_unsigned(1924, 12), 478 => to_unsigned(1355, 12), 479 => to_unsigned(2262, 12), 480 => to_unsigned(1851, 12), 481 => to_unsigned(2367, 12), 482 => to_unsigned(1827, 12), 483 => to_unsigned(2383, 12), 484 => to_unsigned(2392, 12), 485 => to_unsigned(2331, 12), 486 => to_unsigned(2461, 12), 487 => to_unsigned(1776, 12), 488 => to_unsigned(2476, 12), 489 => to_unsigned(1863, 12), 490 => to_unsigned(2053, 12), 491 => to_unsigned(1653, 12), 492 => to_unsigned(1213, 12), 493 => to_unsigned(1198, 12), 494 => to_unsigned(1809, 12), 495 => to_unsigned(1255, 12), 496 => to_unsigned(2252, 12), 497 => to_unsigned(2260, 12), 498 => to_unsigned(2329, 12), 499 => to_unsigned(1418, 12), 500 => to_unsigned(2002, 12), 501 => to_unsigned(2361, 12), 502 => to_unsigned(2577, 12), 503 => to_unsigned(1796, 12), 504 => to_unsigned(1719, 12), 505 => to_unsigned(2087, 12), 506 => to_unsigned(2251, 12), 507 => to_unsigned(2164, 12), 508 => to_unsigned(2465, 12), 509 => to_unsigned(2466, 12), 510 => to_unsigned(1948, 12), 511 => to_unsigned(1417, 12), 512 => to_unsigned(2333, 12), 513 => to_unsigned(2192, 12), 514 => to_unsigned(1853, 12), 515 => to_unsigned(1932, 12), 516 => to_unsigned(1845, 12), 517 => to_unsigned(1601, 12), 518 => to_unsigned(2281, 12), 519 => to_unsigned(1236, 12), 520 => to_unsigned(1612, 12), 521 => to_unsigned(2096, 12), 522 => to_unsigned(1773, 12), 523 => to_unsigned(2038, 12), 524 => to_unsigned(2011, 12), 525 => to_unsigned(2581, 12), 526 => to_unsigned(2108, 12), 527 => to_unsigned(2348, 12), 528 => to_unsigned(1330, 12), 529 => to_unsigned(1889, 12), 530 => to_unsigned(1973, 12), 531 => to_unsigned(1564, 12), 532 => to_unsigned(2490, 12), 533 => to_unsigned(1750, 12), 534 => to_unsigned(2117, 12), 535 => to_unsigned(2117, 12), 536 => to_unsigned(2211, 12), 537 => to_unsigned(1220, 12), 538 => to_unsigned(2330, 12), 539 => to_unsigned(3107, 12), 540 => to_unsigned(1641, 12), 541 => to_unsigned(2197, 12), 542 => to_unsigned(1597, 12), 543 => to_unsigned(2086, 12), 544 => to_unsigned(2029, 12), 545 => to_unsigned(2713, 12), 546 => to_unsigned(2101, 12), 547 => to_unsigned(1702, 12), 548 => to_unsigned(2189, 12), 549 => to_unsigned(2430, 12), 550 => to_unsigned(2306, 12), 551 => to_unsigned(1426, 12), 552 => to_unsigned(1641, 12), 553 => to_unsigned(2456, 12), 554 => to_unsigned(2139, 12), 555 => to_unsigned(1004, 12), 556 => to_unsigned(2797, 12), 557 => to_unsigned(2112, 12), 558 => to_unsigned(1868, 12), 559 => to_unsigned(1976, 12), 560 => to_unsigned(1435, 12), 561 => to_unsigned(2652, 12), 562 => to_unsigned(1886, 12), 563 => to_unsigned(2398, 12), 564 => to_unsigned(2144, 12), 565 => to_unsigned(2487, 12), 566 => to_unsigned(1522, 12), 567 => to_unsigned(2191, 12), 568 => to_unsigned(1548, 12), 569 => to_unsigned(2314, 12), 570 => to_unsigned(1742, 12), 571 => to_unsigned(2068, 12), 572 => to_unsigned(1980, 12), 573 => to_unsigned(958, 12), 574 => to_unsigned(2167, 12), 575 => to_unsigned(1612, 12), 576 => to_unsigned(1503, 12), 577 => to_unsigned(2378, 12), 578 => to_unsigned(2274, 12), 579 => to_unsigned(1989, 12), 580 => to_unsigned(1574, 12), 581 => to_unsigned(1387, 12), 582 => to_unsigned(1992, 12), 583 => to_unsigned(2095, 12), 584 => to_unsigned(2279, 12), 585 => to_unsigned(2572, 12), 586 => to_unsigned(2621, 12), 587 => to_unsigned(1448, 12), 588 => to_unsigned(2598, 12), 589 => to_unsigned(2203, 12), 590 => to_unsigned(2580, 12), 591 => to_unsigned(1591, 12), 592 => to_unsigned(2490, 12), 593 => to_unsigned(1954, 12), 594 => to_unsigned(2101, 12), 595 => to_unsigned(2465, 12), 596 => to_unsigned(2102, 12), 597 => to_unsigned(1492, 12), 598 => to_unsigned(2599, 12), 599 => to_unsigned(1647, 12), 600 => to_unsigned(2317, 12), 601 => to_unsigned(2098, 12), 602 => to_unsigned(1516, 12), 603 => to_unsigned(2223, 12), 604 => to_unsigned(2429, 12), 605 => to_unsigned(2065, 12), 606 => to_unsigned(1940, 12), 607 => to_unsigned(2246, 12), 608 => to_unsigned(1784, 12), 609 => to_unsigned(2050, 12), 610 => to_unsigned(1850, 12), 611 => to_unsigned(1440, 12), 612 => to_unsigned(1861, 12), 613 => to_unsigned(2038, 12), 614 => to_unsigned(2176, 12), 615 => to_unsigned(1948, 12), 616 => to_unsigned(1739, 12), 617 => to_unsigned(2835, 12), 618 => to_unsigned(2001, 12), 619 => to_unsigned(1043, 12), 620 => to_unsigned(1855, 12), 621 => to_unsigned(2367, 12), 622 => to_unsigned(2648, 12), 623 => to_unsigned(2654, 12), 624 => to_unsigned(2138, 12), 625 => to_unsigned(2497, 12), 626 => to_unsigned(2598, 12), 627 => to_unsigned(2345, 12), 628 => to_unsigned(1914, 12), 629 => to_unsigned(2161, 12), 630 => to_unsigned(1770, 12), 631 => to_unsigned(2163, 12), 632 => to_unsigned(2259, 12), 633 => to_unsigned(1959, 12), 634 => to_unsigned(2150, 12), 635 => to_unsigned(1332, 12), 636 => to_unsigned(1401, 12), 637 => to_unsigned(1780, 12), 638 => to_unsigned(1839, 12), 639 => to_unsigned(2399, 12), 640 => to_unsigned(2965, 12), 641 => to_unsigned(1649, 12), 642 => to_unsigned(1951, 12), 643 => to_unsigned(2186, 12), 644 => to_unsigned(1815, 12), 645 => to_unsigned(1668, 12), 646 => to_unsigned(1718, 12), 647 => to_unsigned(1977, 12), 648 => to_unsigned(2345, 12), 649 => to_unsigned(1649, 12), 650 => to_unsigned(2256, 12), 651 => to_unsigned(1488, 12), 652 => to_unsigned(2292, 12), 653 => to_unsigned(2581, 12), 654 => to_unsigned(2904, 12), 655 => to_unsigned(2099, 12), 656 => to_unsigned(2004, 12), 657 => to_unsigned(2392, 12), 658 => to_unsigned(2222, 12), 659 => to_unsigned(1925, 12), 660 => to_unsigned(2395, 12), 661 => to_unsigned(1770, 12), 662 => to_unsigned(2328, 12), 663 => to_unsigned(2189, 12), 664 => to_unsigned(2349, 12), 665 => to_unsigned(1989, 12), 666 => to_unsigned(2165, 12), 667 => to_unsigned(1736, 12), 668 => to_unsigned(2525, 12), 669 => to_unsigned(2410, 12), 670 => to_unsigned(2862, 12), 671 => to_unsigned(2258, 12), 672 => to_unsigned(2096, 12), 673 => to_unsigned(1924, 12), 674 => to_unsigned(1364, 12), 675 => to_unsigned(1939, 12), 676 => to_unsigned(2091, 12), 677 => to_unsigned(2398, 12), 678 => to_unsigned(1836, 12), 679 => to_unsigned(1921, 12), 680 => to_unsigned(1711, 12), 681 => to_unsigned(2284, 12), 682 => to_unsigned(2564, 12), 683 => to_unsigned(2042, 12), 684 => to_unsigned(2127, 12), 685 => to_unsigned(1571, 12), 686 => to_unsigned(1402, 12), 687 => to_unsigned(1132, 12), 688 => to_unsigned(1257, 12), 689 => to_unsigned(2369, 12), 690 => to_unsigned(1888, 12), 691 => to_unsigned(2046, 12), 692 => to_unsigned(1851, 12), 693 => to_unsigned(2558, 12), 694 => to_unsigned(1700, 12), 695 => to_unsigned(998, 12), 696 => to_unsigned(2189, 12), 697 => to_unsigned(1690, 12), 698 => to_unsigned(2297, 12), 699 => to_unsigned(1646, 12), 700 => to_unsigned(2383, 12), 701 => to_unsigned(2366, 12), 702 => to_unsigned(2167, 12), 703 => to_unsigned(2831, 12), 704 => to_unsigned(2140, 12), 705 => to_unsigned(1819, 12), 706 => to_unsigned(2099, 12), 707 => to_unsigned(1551, 12), 708 => to_unsigned(2419, 12), 709 => to_unsigned(2077, 12), 710 => to_unsigned(2100, 12), 711 => to_unsigned(2356, 12), 712 => to_unsigned(2200, 12), 713 => to_unsigned(1915, 12), 714 => to_unsigned(1314, 12), 715 => to_unsigned(1767, 12), 716 => to_unsigned(1617, 12), 717 => to_unsigned(1975, 12), 718 => to_unsigned(2075, 12), 719 => to_unsigned(1808, 12), 720 => to_unsigned(2395, 12), 721 => to_unsigned(2022, 12), 722 => to_unsigned(2924, 12), 723 => to_unsigned(2592, 12), 724 => to_unsigned(2301, 12), 725 => to_unsigned(2447, 12), 726 => to_unsigned(961, 12), 727 => to_unsigned(1941, 12), 728 => to_unsigned(2148, 12), 729 => to_unsigned(2414, 12), 730 => to_unsigned(1999, 12), 731 => to_unsigned(2472, 12), 732 => to_unsigned(1894, 12), 733 => to_unsigned(2568, 12), 734 => to_unsigned(2420, 12), 735 => to_unsigned(1714, 12), 736 => to_unsigned(1801, 12), 737 => to_unsigned(1836, 12), 738 => to_unsigned(1834, 12), 739 => to_unsigned(1906, 12), 740 => to_unsigned(2327, 12), 741 => to_unsigned(2118, 12), 742 => to_unsigned(1234, 12), 743 => to_unsigned(2082, 12), 744 => to_unsigned(3155, 12), 745 => to_unsigned(1761, 12), 746 => to_unsigned(2173, 12), 747 => to_unsigned(2217, 12), 748 => to_unsigned(2525, 12), 749 => to_unsigned(2083, 12), 750 => to_unsigned(2168, 12), 751 => to_unsigned(2423, 12), 752 => to_unsigned(2707, 12), 753 => to_unsigned(1829, 12), 754 => to_unsigned(2237, 12), 755 => to_unsigned(1615, 12), 756 => to_unsigned(2099, 12), 757 => to_unsigned(2239, 12), 758 => to_unsigned(2639, 12), 759 => to_unsigned(2159, 12), 760 => to_unsigned(2047, 12), 761 => to_unsigned(2429, 12), 762 => to_unsigned(2439, 12), 763 => to_unsigned(1967, 12), 764 => to_unsigned(1837, 12), 765 => to_unsigned(2312, 12), 766 => to_unsigned(2380, 12), 767 => to_unsigned(2601, 12), 768 => to_unsigned(2307, 12), 769 => to_unsigned(2115, 12), 770 => to_unsigned(2068, 12), 771 => to_unsigned(2264, 12), 772 => to_unsigned(2558, 12), 773 => to_unsigned(1870, 12), 774 => to_unsigned(1750, 12), 775 => to_unsigned(1788, 12), 776 => to_unsigned(2684, 12), 777 => to_unsigned(1571, 12), 778 => to_unsigned(1898, 12), 779 => to_unsigned(2019, 12), 780 => to_unsigned(1736, 12), 781 => to_unsigned(2426, 12), 782 => to_unsigned(2628, 12), 783 => to_unsigned(2369, 12), 784 => to_unsigned(2200, 12), 785 => to_unsigned(2015, 12), 786 => to_unsigned(1674, 12), 787 => to_unsigned(2695, 12), 788 => to_unsigned(1834, 12), 789 => to_unsigned(2188, 12), 790 => to_unsigned(1658, 12), 791 => to_unsigned(1789, 12), 792 => to_unsigned(2054, 12), 793 => to_unsigned(2449, 12), 794 => to_unsigned(1297, 12), 795 => to_unsigned(2114, 12), 796 => to_unsigned(2608, 12), 797 => to_unsigned(2023, 12), 798 => to_unsigned(1935, 12), 799 => to_unsigned(3038, 12), 800 => to_unsigned(1839, 12), 801 => to_unsigned(2108, 12), 802 => to_unsigned(2547, 12), 803 => to_unsigned(1777, 12), 804 => to_unsigned(1844, 12), 805 => to_unsigned(1986, 12), 806 => to_unsigned(1703, 12), 807 => to_unsigned(2060, 12), 808 => to_unsigned(2488, 12), 809 => to_unsigned(2374, 12), 810 => to_unsigned(2478, 12), 811 => to_unsigned(1842, 12), 812 => to_unsigned(2276, 12), 813 => to_unsigned(2340, 12), 814 => to_unsigned(2819, 12), 815 => to_unsigned(2492, 12), 816 => to_unsigned(2029, 12), 817 => to_unsigned(1747, 12), 818 => to_unsigned(2312, 12), 819 => to_unsigned(2137, 12), 820 => to_unsigned(1906, 12), 821 => to_unsigned(2719, 12), 822 => to_unsigned(1650, 12), 823 => to_unsigned(1947, 12), 824 => to_unsigned(1625, 12), 825 => to_unsigned(2648, 12), 826 => to_unsigned(2472, 12), 827 => to_unsigned(1809, 12), 828 => to_unsigned(1406, 12), 829 => to_unsigned(2408, 12), 830 => to_unsigned(2096, 12), 831 => to_unsigned(2066, 12), 832 => to_unsigned(2494, 12), 833 => to_unsigned(1596, 12), 834 => to_unsigned(2018, 12), 835 => to_unsigned(2357, 12), 836 => to_unsigned(1841, 12), 837 => to_unsigned(1768, 12), 838 => to_unsigned(2157, 12), 839 => to_unsigned(1842, 12), 840 => to_unsigned(2157, 12), 841 => to_unsigned(2096, 12), 842 => to_unsigned(2160, 12), 843 => to_unsigned(1828, 12), 844 => to_unsigned(1662, 12), 845 => to_unsigned(1832, 12), 846 => to_unsigned(1872, 12), 847 => to_unsigned(1557, 12), 848 => to_unsigned(2290, 12), 849 => to_unsigned(2038, 12), 850 => to_unsigned(1926, 12), 851 => to_unsigned(1678, 12), 852 => to_unsigned(1935, 12), 853 => to_unsigned(2220, 12), 854 => to_unsigned(1618, 12), 855 => to_unsigned(2026, 12), 856 => to_unsigned(2578, 12), 857 => to_unsigned(2601, 12), 858 => to_unsigned(2858, 12), 859 => to_unsigned(1946, 12), 860 => to_unsigned(2290, 12), 861 => to_unsigned(1960, 12), 862 => to_unsigned(2332, 12), 863 => to_unsigned(1972, 12), 864 => to_unsigned(2430, 12), 865 => to_unsigned(2149, 12), 866 => to_unsigned(2108, 12), 867 => to_unsigned(2009, 12), 868 => to_unsigned(1631, 12), 869 => to_unsigned(2031, 12), 870 => to_unsigned(1459, 12), 871 => to_unsigned(2180, 12), 872 => to_unsigned(1622, 12), 873 => to_unsigned(1908, 12), 874 => to_unsigned(2059, 12), 875 => to_unsigned(1568, 12), 876 => to_unsigned(1994, 12), 877 => to_unsigned(1902, 12), 878 => to_unsigned(1964, 12), 879 => to_unsigned(1265, 12), 880 => to_unsigned(1106, 12), 881 => to_unsigned(2330, 12), 882 => to_unsigned(1990, 12), 883 => to_unsigned(1545, 12), 884 => to_unsigned(1850, 12), 885 => to_unsigned(2221, 12), 886 => to_unsigned(1887, 12), 887 => to_unsigned(2070, 12), 888 => to_unsigned(1746, 12), 889 => to_unsigned(1685, 12), 890 => to_unsigned(920, 12), 891 => to_unsigned(2346, 12), 892 => to_unsigned(1632, 12), 893 => to_unsigned(2078, 12), 894 => to_unsigned(1362, 12), 895 => to_unsigned(2020, 12), 896 => to_unsigned(1669, 12), 897 => to_unsigned(2173, 12), 898 => to_unsigned(1265, 12), 899 => to_unsigned(2600, 12), 900 => to_unsigned(2237, 12), 901 => to_unsigned(2033, 12), 902 => to_unsigned(1807, 12), 903 => to_unsigned(2129, 12), 904 => to_unsigned(2054, 12), 905 => to_unsigned(2171, 12), 906 => to_unsigned(2231, 12), 907 => to_unsigned(1665, 12), 908 => to_unsigned(2119, 12), 909 => to_unsigned(2120, 12), 910 => to_unsigned(2559, 12), 911 => to_unsigned(2099, 12), 912 => to_unsigned(1886, 12), 913 => to_unsigned(2000, 12), 914 => to_unsigned(2321, 12), 915 => to_unsigned(1891, 12), 916 => to_unsigned(2051, 12), 917 => to_unsigned(1453, 12), 918 => to_unsigned(1964, 12), 919 => to_unsigned(1585, 12), 920 => to_unsigned(1426, 12), 921 => to_unsigned(1583, 12), 922 => to_unsigned(2577, 12), 923 => to_unsigned(2174, 12), 924 => to_unsigned(2384, 12), 925 => to_unsigned(2071, 12), 926 => to_unsigned(2003, 12), 927 => to_unsigned(2113, 12), 928 => to_unsigned(2068, 12), 929 => to_unsigned(2075, 12), 930 => to_unsigned(1958, 12), 931 => to_unsigned(1637, 12), 932 => to_unsigned(1741, 12), 933 => to_unsigned(2472, 12), 934 => to_unsigned(1595, 12), 935 => to_unsigned(2107, 12), 936 => to_unsigned(2632, 12), 937 => to_unsigned(1694, 12), 938 => to_unsigned(1983, 12), 939 => to_unsigned(1313, 12), 940 => to_unsigned(1717, 12), 941 => to_unsigned(1774, 12), 942 => to_unsigned(1985, 12), 943 => to_unsigned(2149, 12), 944 => to_unsigned(2182, 12), 945 => to_unsigned(2356, 12), 946 => to_unsigned(2192, 12), 947 => to_unsigned(2938, 12), 948 => to_unsigned(1971, 12), 949 => to_unsigned(2262, 12), 950 => to_unsigned(2231, 12), 951 => to_unsigned(2582, 12), 952 => to_unsigned(2479, 12), 953 => to_unsigned(2472, 12), 954 => to_unsigned(1121, 12), 955 => to_unsigned(2510, 12), 956 => to_unsigned(1962, 12), 957 => to_unsigned(1667, 12), 958 => to_unsigned(2218, 12), 959 => to_unsigned(1658, 12), 960 => to_unsigned(2379, 12), 961 => to_unsigned(2645, 12), 962 => to_unsigned(1915, 12), 963 => to_unsigned(1746, 12), 964 => to_unsigned(2095, 12), 965 => to_unsigned(2165, 12), 966 => to_unsigned(1708, 12), 967 => to_unsigned(2437, 12), 968 => to_unsigned(2208, 12), 969 => to_unsigned(2463, 12), 970 => to_unsigned(1193, 12), 971 => to_unsigned(2181, 12), 972 => to_unsigned(1598, 12), 973 => to_unsigned(2007, 12), 974 => to_unsigned(2267, 12), 975 => to_unsigned(1903, 12), 976 => to_unsigned(2076, 12), 977 => to_unsigned(2695, 12), 978 => to_unsigned(1044, 12), 979 => to_unsigned(2121, 12), 980 => to_unsigned(1958, 12), 981 => to_unsigned(1735, 12), 982 => to_unsigned(1758, 12), 983 => to_unsigned(1927, 12), 984 => to_unsigned(1912, 12), 985 => to_unsigned(2371, 12), 986 => to_unsigned(2730, 12), 987 => to_unsigned(1954, 12), 988 => to_unsigned(1924, 12), 989 => to_unsigned(2450, 12), 990 => to_unsigned(2118, 12), 991 => to_unsigned(2284, 12), 992 => to_unsigned(1968, 12), 993 => to_unsigned(2218, 12), 994 => to_unsigned(1503, 12), 995 => to_unsigned(2068, 12), 996 => to_unsigned(2328, 12), 997 => to_unsigned(1943, 12), 998 => to_unsigned(2089, 12), 999 => to_unsigned(1841, 12), 1000 => to_unsigned(2532, 12), 1001 => to_unsigned(1590, 12), 1002 => to_unsigned(2424, 12), 1003 => to_unsigned(1789, 12), 1004 => to_unsigned(1504, 12), 1005 => to_unsigned(2428, 12), 1006 => to_unsigned(2279, 12), 1007 => to_unsigned(1818, 12), 1008 => to_unsigned(2239, 12), 1009 => to_unsigned(1589, 12), 1010 => to_unsigned(1737, 12), 1011 => to_unsigned(1427, 12), 1012 => to_unsigned(2083, 12), 1013 => to_unsigned(1743, 12), 1014 => to_unsigned(1370, 12), 1015 => to_unsigned(1724, 12), 1016 => to_unsigned(2193, 12), 1017 => to_unsigned(2388, 12), 1018 => to_unsigned(2100, 12), 1019 => to_unsigned(2735, 12), 1020 => to_unsigned(2038, 12), 1021 => to_unsigned(1793, 12), 1022 => to_unsigned(2279, 12), 1023 => to_unsigned(1929, 12), 1024 => to_unsigned(2549, 12), 1025 => to_unsigned(2148, 12), 1026 => to_unsigned(1894, 12), 1027 => to_unsigned(1682, 12), 1028 => to_unsigned(2058, 12), 1029 => to_unsigned(2478, 12), 1030 => to_unsigned(1709, 12), 1031 => to_unsigned(1870, 12), 1032 => to_unsigned(2354, 12), 1033 => to_unsigned(1847, 12), 1034 => to_unsigned(2241, 12), 1035 => to_unsigned(2511, 12), 1036 => to_unsigned(2044, 12), 1037 => to_unsigned(1926, 12), 1038 => to_unsigned(1841, 12), 1039 => to_unsigned(2658, 12), 1040 => to_unsigned(2587, 12), 1041 => to_unsigned(1836, 12), 1042 => to_unsigned(2197, 12), 1043 => to_unsigned(2462, 12), 1044 => to_unsigned(3149, 12), 1045 => to_unsigned(2306, 12), 1046 => to_unsigned(1765, 12), 1047 => to_unsigned(2162, 12), 1048 => to_unsigned(2144, 12), 1049 => to_unsigned(2286, 12), 1050 => to_unsigned(1779, 12), 1051 => to_unsigned(1670, 12), 1052 => to_unsigned(1665, 12), 1053 => to_unsigned(2289, 12), 1054 => to_unsigned(2643, 12), 1055 => to_unsigned(2363, 12), 1056 => to_unsigned(2194, 12), 1057 => to_unsigned(2345, 12), 1058 => to_unsigned(1799, 12), 1059 => to_unsigned(1579, 12), 1060 => to_unsigned(1965, 12), 1061 => to_unsigned(1345, 12), 1062 => to_unsigned(2556, 12), 1063 => to_unsigned(1699, 12), 1064 => to_unsigned(2235, 12), 1065 => to_unsigned(2068, 12), 1066 => to_unsigned(2825, 12), 1067 => to_unsigned(2207, 12), 1068 => to_unsigned(2396, 12), 1069 => to_unsigned(2358, 12), 1070 => to_unsigned(2192, 12), 1071 => to_unsigned(2483, 12), 1072 => to_unsigned(1712, 12), 1073 => to_unsigned(1477, 12), 1074 => to_unsigned(1103, 12), 1075 => to_unsigned(2690, 12), 1076 => to_unsigned(1653, 12), 1077 => to_unsigned(1840, 12), 1078 => to_unsigned(2563, 12), 1079 => to_unsigned(2138, 12), 1080 => to_unsigned(2705, 12), 1081 => to_unsigned(1985, 12), 1082 => to_unsigned(2190, 12), 1083 => to_unsigned(2004, 12), 1084 => to_unsigned(2219, 12), 1085 => to_unsigned(2134, 12), 1086 => to_unsigned(1658, 12), 1087 => to_unsigned(2345, 12), 1088 => to_unsigned(1933, 12), 1089 => to_unsigned(2584, 12), 1090 => to_unsigned(1818, 12), 1091 => to_unsigned(2458, 12), 1092 => to_unsigned(2571, 12), 1093 => to_unsigned(2091, 12), 1094 => to_unsigned(2205, 12), 1095 => to_unsigned(2102, 12), 1096 => to_unsigned(2189, 12), 1097 => to_unsigned(1664, 12), 1098 => to_unsigned(1784, 12), 1099 => to_unsigned(1688, 12), 1100 => to_unsigned(1440, 12), 1101 => to_unsigned(2160, 12), 1102 => to_unsigned(2685, 12), 1103 => to_unsigned(1995, 12), 1104 => to_unsigned(2405, 12), 1105 => to_unsigned(2235, 12), 1106 => to_unsigned(2435, 12), 1107 => to_unsigned(2115, 12), 1108 => to_unsigned(2029, 12), 1109 => to_unsigned(1311, 12), 1110 => to_unsigned(2102, 12), 1111 => to_unsigned(1865, 12), 1112 => to_unsigned(1073, 12), 1113 => to_unsigned(1807, 12), 1114 => to_unsigned(2222, 12), 1115 => to_unsigned(1650, 12), 1116 => to_unsigned(2259, 12), 1117 => to_unsigned(2396, 12), 1118 => to_unsigned(2037, 12), 1119 => to_unsigned(2378, 12), 1120 => to_unsigned(1578, 12), 1121 => to_unsigned(2199, 12), 1122 => to_unsigned(1915, 12), 1123 => to_unsigned(933, 12), 1124 => to_unsigned(1976, 12), 1125 => to_unsigned(1712, 12), 1126 => to_unsigned(2423, 12), 1127 => to_unsigned(2221, 12), 1128 => to_unsigned(2156, 12), 1129 => to_unsigned(1613, 12), 1130 => to_unsigned(1765, 12), 1131 => to_unsigned(1436, 12), 1132 => to_unsigned(2111, 12), 1133 => to_unsigned(1390, 12), 1134 => to_unsigned(1892, 12), 1135 => to_unsigned(2339, 12), 1136 => to_unsigned(1381, 12), 1137 => to_unsigned(2167, 12), 1138 => to_unsigned(1901, 12), 1139 => to_unsigned(1481, 12), 1140 => to_unsigned(1989, 12), 1141 => to_unsigned(1994, 12), 1142 => to_unsigned(2339, 12), 1143 => to_unsigned(1536, 12), 1144 => to_unsigned(2241, 12), 1145 => to_unsigned(1995, 12), 1146 => to_unsigned(2331, 12), 1147 => to_unsigned(1840, 12), 1148 => to_unsigned(2092, 12), 1149 => to_unsigned(2307, 12), 1150 => to_unsigned(2072, 12), 1151 => to_unsigned(2119, 12), 1152 => to_unsigned(2499, 12), 1153 => to_unsigned(1960, 12), 1154 => to_unsigned(2416, 12), 1155 => to_unsigned(2449, 12), 1156 => to_unsigned(1533, 12), 1157 => to_unsigned(1787, 12), 1158 => to_unsigned(2147, 12), 1159 => to_unsigned(2949, 12), 1160 => to_unsigned(2403, 12), 1161 => to_unsigned(1872, 12), 1162 => to_unsigned(2563, 12), 1163 => to_unsigned(1944, 12), 1164 => to_unsigned(1519, 12), 1165 => to_unsigned(2267, 12), 1166 => to_unsigned(2498, 12), 1167 => to_unsigned(1595, 12), 1168 => to_unsigned(2716, 12), 1169 => to_unsigned(1863, 12), 1170 => to_unsigned(2026, 12), 1171 => to_unsigned(1748, 12), 1172 => to_unsigned(3040, 12), 1173 => to_unsigned(1869, 12), 1174 => to_unsigned(1788, 12), 1175 => to_unsigned(2050, 12), 1176 => to_unsigned(2347, 12), 1177 => to_unsigned(2337, 12), 1178 => to_unsigned(2452, 12), 1179 => to_unsigned(1418, 12), 1180 => to_unsigned(1837, 12), 1181 => to_unsigned(1993, 12), 1182 => to_unsigned(1580, 12), 1183 => to_unsigned(2092, 12), 1184 => to_unsigned(2110, 12), 1185 => to_unsigned(2200, 12), 1186 => to_unsigned(3132, 12), 1187 => to_unsigned(2639, 12), 1188 => to_unsigned(2052, 12), 1189 => to_unsigned(1428, 12), 1190 => to_unsigned(2148, 12), 1191 => to_unsigned(1507, 12), 1192 => to_unsigned(1193, 12), 1193 => to_unsigned(2113, 12), 1194 => to_unsigned(1922, 12), 1195 => to_unsigned(2332, 12), 1196 => to_unsigned(2682, 12), 1197 => to_unsigned(2237, 12), 1198 => to_unsigned(2296, 12), 1199 => to_unsigned(2133, 12), 1200 => to_unsigned(2158, 12), 1201 => to_unsigned(2638, 12), 1202 => to_unsigned(2720, 12), 1203 => to_unsigned(1829, 12), 1204 => to_unsigned(1613, 12), 1205 => to_unsigned(2210, 12), 1206 => to_unsigned(1688, 12), 1207 => to_unsigned(2122, 12), 1208 => to_unsigned(1633, 12), 1209 => to_unsigned(1861, 12), 1210 => to_unsigned(2774, 12), 1211 => to_unsigned(2951, 12), 1212 => to_unsigned(1900, 12), 1213 => to_unsigned(2512, 12), 1214 => to_unsigned(2585, 12), 1215 => to_unsigned(1809, 12), 1216 => to_unsigned(2351, 12), 1217 => to_unsigned(1608, 12), 1218 => to_unsigned(1490, 12), 1219 => to_unsigned(1879, 12), 1220 => to_unsigned(1770, 12), 1221 => to_unsigned(1692, 12), 1222 => to_unsigned(1822, 12), 1223 => to_unsigned(1995, 12), 1224 => to_unsigned(1781, 12), 1225 => to_unsigned(2292, 12), 1226 => to_unsigned(1941, 12), 1227 => to_unsigned(2207, 12), 1228 => to_unsigned(1863, 12), 1229 => to_unsigned(2186, 12), 1230 => to_unsigned(1949, 12), 1231 => to_unsigned(2339, 12), 1232 => to_unsigned(2143, 12), 1233 => to_unsigned(2708, 12), 1234 => to_unsigned(2306, 12), 1235 => to_unsigned(1721, 12), 1236 => to_unsigned(2272, 12), 1237 => to_unsigned(1903, 12), 1238 => to_unsigned(2354, 12), 1239 => to_unsigned(1742, 12), 1240 => to_unsigned(1684, 12), 1241 => to_unsigned(2517, 12), 1242 => to_unsigned(1663, 12), 1243 => to_unsigned(1821, 12), 1244 => to_unsigned(1932, 12), 1245 => to_unsigned(2089, 12), 1246 => to_unsigned(2595, 12), 1247 => to_unsigned(2026, 12), 1248 => to_unsigned(1521, 12), 1249 => to_unsigned(1192, 12), 1250 => to_unsigned(2282, 12), 1251 => to_unsigned(2605, 12), 1252 => to_unsigned(2207, 12), 1253 => to_unsigned(1832, 12), 1254 => to_unsigned(1876, 12), 1255 => to_unsigned(2039, 12), 1256 => to_unsigned(2406, 12), 1257 => to_unsigned(2370, 12), 1258 => to_unsigned(1901, 12), 1259 => to_unsigned(2319, 12), 1260 => to_unsigned(2505, 12), 1261 => to_unsigned(2023, 12), 1262 => to_unsigned(1935, 12), 1263 => to_unsigned(1991, 12), 1264 => to_unsigned(2570, 12), 1265 => to_unsigned(1511, 12), 1266 => to_unsigned(3294, 12), 1267 => to_unsigned(2312, 12), 1268 => to_unsigned(2491, 12), 1269 => to_unsigned(1964, 12), 1270 => to_unsigned(1997, 12), 1271 => to_unsigned(1911, 12), 1272 => to_unsigned(1615, 12), 1273 => to_unsigned(2408, 12), 1274 => to_unsigned(2725, 12), 1275 => to_unsigned(2417, 12), 1276 => to_unsigned(2287, 12), 1277 => to_unsigned(2778, 12), 1278 => to_unsigned(2258, 12), 1279 => to_unsigned(1619, 12), 1280 => to_unsigned(1983, 12), 1281 => to_unsigned(2664, 12), 1282 => to_unsigned(2248, 12), 1283 => to_unsigned(1440, 12), 1284 => to_unsigned(2440, 12), 1285 => to_unsigned(2050, 12), 1286 => to_unsigned(1608, 12), 1287 => to_unsigned(2261, 12), 1288 => to_unsigned(2481, 12), 1289 => to_unsigned(1486, 12), 1290 => to_unsigned(1847, 12), 1291 => to_unsigned(2644, 12), 1292 => to_unsigned(1635, 12), 1293 => to_unsigned(1865, 12), 1294 => to_unsigned(1783, 12), 1295 => to_unsigned(2158, 12), 1296 => to_unsigned(1802, 12), 1297 => to_unsigned(1392, 12), 1298 => to_unsigned(2124, 12), 1299 => to_unsigned(1869, 12), 1300 => to_unsigned(2290, 12), 1301 => to_unsigned(1536, 12), 1302 => to_unsigned(1851, 12), 1303 => to_unsigned(2083, 12), 1304 => to_unsigned(2363, 12), 1305 => to_unsigned(1929, 12), 1306 => to_unsigned(1879, 12), 1307 => to_unsigned(2729, 12), 1308 => to_unsigned(1682, 12), 1309 => to_unsigned(1888, 12), 1310 => to_unsigned(2350, 12), 1311 => to_unsigned(2484, 12), 1312 => to_unsigned(2015, 12), 1313 => to_unsigned(2808, 12), 1314 => to_unsigned(2292, 12), 1315 => to_unsigned(2373, 12), 1316 => to_unsigned(1742, 12), 1317 => to_unsigned(2007, 12), 1318 => to_unsigned(1780, 12), 1319 => to_unsigned(1827, 12), 1320 => to_unsigned(1967, 12), 1321 => to_unsigned(1630, 12), 1322 => to_unsigned(2259, 12), 1323 => to_unsigned(1572, 12), 1324 => to_unsigned(2020, 12), 1325 => to_unsigned(2485, 12), 1326 => to_unsigned(1869, 12), 1327 => to_unsigned(2370, 12), 1328 => to_unsigned(2189, 12), 1329 => to_unsigned(2547, 12), 1330 => to_unsigned(2011, 12), 1331 => to_unsigned(2803, 12), 1332 => to_unsigned(1763, 12), 1333 => to_unsigned(2128, 12), 1334 => to_unsigned(2018, 12), 1335 => to_unsigned(2587, 12), 1336 => to_unsigned(1922, 12), 1337 => to_unsigned(1811, 12), 1338 => to_unsigned(2245, 12), 1339 => to_unsigned(2242, 12), 1340 => to_unsigned(1946, 12), 1341 => to_unsigned(1842, 12), 1342 => to_unsigned(1648, 12), 1343 => to_unsigned(2177, 12), 1344 => to_unsigned(1887, 12), 1345 => to_unsigned(2160, 12), 1346 => to_unsigned(2149, 12), 1347 => to_unsigned(1917, 12), 1348 => to_unsigned(2890, 12), 1349 => to_unsigned(2638, 12), 1350 => to_unsigned(1665, 12), 1351 => to_unsigned(1717, 12), 1352 => to_unsigned(2053, 12), 1353 => to_unsigned(1974, 12), 1354 => to_unsigned(2326, 12), 1355 => to_unsigned(1941, 12), 1356 => to_unsigned(1588, 12), 1357 => to_unsigned(1374, 12), 1358 => to_unsigned(2144, 12), 1359 => to_unsigned(1937, 12), 1360 => to_unsigned(2135, 12), 1361 => to_unsigned(1902, 12), 1362 => to_unsigned(2144, 12), 1363 => to_unsigned(2284, 12), 1364 => to_unsigned(2026, 12), 1365 => to_unsigned(2175, 12), 1366 => to_unsigned(2334, 12), 1367 => to_unsigned(1957, 12), 1368 => to_unsigned(1885, 12), 1369 => to_unsigned(2187, 12), 1370 => to_unsigned(1618, 12), 1371 => to_unsigned(2591, 12), 1372 => to_unsigned(1989, 12), 1373 => to_unsigned(2296, 12), 1374 => to_unsigned(2178, 12), 1375 => to_unsigned(1768, 12), 1376 => to_unsigned(2591, 12), 1377 => to_unsigned(1796, 12), 1378 => to_unsigned(1864, 12), 1379 => to_unsigned(1537, 12), 1380 => to_unsigned(1921, 12), 1381 => to_unsigned(2167, 12), 1382 => to_unsigned(1489, 12), 1383 => to_unsigned(1994, 12), 1384 => to_unsigned(2048, 12), 1385 => to_unsigned(2546, 12), 1386 => to_unsigned(1516, 12), 1387 => to_unsigned(2179, 12), 1388 => to_unsigned(2619, 12), 1389 => to_unsigned(1969, 12), 1390 => to_unsigned(1787, 12), 1391 => to_unsigned(2062, 12), 1392 => to_unsigned(2792, 12), 1393 => to_unsigned(2069, 12), 1394 => to_unsigned(2449, 12), 1395 => to_unsigned(2123, 12), 1396 => to_unsigned(1199, 12), 1397 => to_unsigned(2082, 12), 1398 => to_unsigned(1881, 12), 1399 => to_unsigned(2141, 12), 1400 => to_unsigned(1942, 12), 1401 => to_unsigned(1994, 12), 1402 => to_unsigned(1824, 12), 1403 => to_unsigned(2257, 12), 1404 => to_unsigned(1910, 12), 1405 => to_unsigned(2281, 12), 1406 => to_unsigned(2460, 12), 1407 => to_unsigned(2298, 12), 1408 => to_unsigned(1935, 12), 1409 => to_unsigned(2120, 12), 1410 => to_unsigned(1887, 12), 1411 => to_unsigned(1713, 12), 1412 => to_unsigned(1684, 12), 1413 => to_unsigned(1623, 12), 1414 => to_unsigned(2239, 12), 1415 => to_unsigned(1901, 12), 1416 => to_unsigned(1544, 12), 1417 => to_unsigned(1839, 12), 1418 => to_unsigned(1932, 12), 1419 => to_unsigned(1296, 12), 1420 => to_unsigned(1834, 12), 1421 => to_unsigned(1739, 12), 1422 => to_unsigned(2117, 12), 1423 => to_unsigned(2599, 12), 1424 => to_unsigned(2463, 12), 1425 => to_unsigned(1726, 12), 1426 => to_unsigned(2142, 12), 1427 => to_unsigned(1827, 12), 1428 => to_unsigned(2418, 12), 1429 => to_unsigned(1790, 12), 1430 => to_unsigned(2197, 12), 1431 => to_unsigned(2109, 12), 1432 => to_unsigned(2186, 12), 1433 => to_unsigned(2346, 12), 1434 => to_unsigned(2636, 12), 1435 => to_unsigned(1698, 12), 1436 => to_unsigned(2147, 12), 1437 => to_unsigned(1938, 12), 1438 => to_unsigned(2103, 12), 1439 => to_unsigned(1464, 12), 1440 => to_unsigned(1341, 12), 1441 => to_unsigned(2147, 12), 1442 => to_unsigned(1572, 12), 1443 => to_unsigned(1849, 12), 1444 => to_unsigned(2713, 12), 1445 => to_unsigned(2414, 12), 1446 => to_unsigned(1433, 12), 1447 => to_unsigned(2304, 12), 1448 => to_unsigned(2689, 12), 1449 => to_unsigned(2157, 12), 1450 => to_unsigned(1449, 12), 1451 => to_unsigned(2205, 12), 1452 => to_unsigned(1799, 12), 1453 => to_unsigned(2377, 12), 1454 => to_unsigned(1958, 12), 1455 => to_unsigned(2257, 12), 1456 => to_unsigned(1593, 12), 1457 => to_unsigned(2534, 12), 1458 => to_unsigned(2693, 12), 1459 => to_unsigned(2193, 12), 1460 => to_unsigned(1960, 12), 1461 => to_unsigned(2068, 12), 1462 => to_unsigned(1851, 12), 1463 => to_unsigned(1919, 12), 1464 => to_unsigned(1829, 12), 1465 => to_unsigned(1899, 12), 1466 => to_unsigned(1667, 12), 1467 => to_unsigned(1857, 12), 1468 => to_unsigned(2332, 12), 1469 => to_unsigned(1972, 12), 1470 => to_unsigned(1158, 12), 1471 => to_unsigned(1731, 12), 1472 => to_unsigned(2477, 12), 1473 => to_unsigned(1709, 12), 1474 => to_unsigned(2375, 12), 1475 => to_unsigned(2229, 12), 1476 => to_unsigned(1993, 12), 1477 => to_unsigned(2375, 12), 1478 => to_unsigned(2554, 12), 1479 => to_unsigned(1753, 12), 1480 => to_unsigned(2036, 12), 1481 => to_unsigned(1660, 12), 1482 => to_unsigned(1507, 12), 1483 => to_unsigned(2502, 12), 1484 => to_unsigned(2080, 12), 1485 => to_unsigned(2507, 12), 1486 => to_unsigned(2655, 12), 1487 => to_unsigned(1605, 12), 1488 => to_unsigned(1932, 12), 1489 => to_unsigned(2261, 12), 1490 => to_unsigned(2596, 12), 1491 => to_unsigned(2345, 12), 1492 => to_unsigned(2549, 12), 1493 => to_unsigned(2952, 12), 1494 => to_unsigned(2367, 12), 1495 => to_unsigned(1613, 12), 1496 => to_unsigned(2189, 12), 1497 => to_unsigned(2262, 12), 1498 => to_unsigned(1717, 12), 1499 => to_unsigned(2629, 12), 1500 => to_unsigned(1974, 12), 1501 => to_unsigned(2039, 12), 1502 => to_unsigned(2109, 12), 1503 => to_unsigned(2438, 12), 1504 => to_unsigned(2423, 12), 1505 => to_unsigned(1611, 12), 1506 => to_unsigned(2133, 12), 1507 => to_unsigned(2954, 12), 1508 => to_unsigned(2148, 12), 1509 => to_unsigned(1836, 12), 1510 => to_unsigned(1637, 12), 1511 => to_unsigned(1709, 12), 1512 => to_unsigned(2410, 12), 1513 => to_unsigned(1943, 12), 1514 => to_unsigned(1509, 12), 1515 => to_unsigned(1877, 12), 1516 => to_unsigned(2191, 12), 1517 => to_unsigned(1884, 12), 1518 => to_unsigned(2181, 12), 1519 => to_unsigned(2745, 12), 1520 => to_unsigned(2196, 12), 1521 => to_unsigned(1723, 12), 1522 => to_unsigned(2326, 12), 1523 => to_unsigned(2602, 12), 1524 => to_unsigned(2020, 12), 1525 => to_unsigned(2175, 12), 1526 => to_unsigned(1986, 12), 1527 => to_unsigned(1357, 12), 1528 => to_unsigned(1779, 12), 1529 => to_unsigned(2626, 12), 1530 => to_unsigned(2465, 12), 1531 => to_unsigned(2214, 12), 1532 => to_unsigned(2125, 12), 1533 => to_unsigned(1483, 12), 1534 => to_unsigned(2841, 12), 1535 => to_unsigned(2433, 12), 1536 => to_unsigned(1812, 12), 1537 => to_unsigned(2512, 12), 1538 => to_unsigned(1860, 12), 1539 => to_unsigned(1493, 12), 1540 => to_unsigned(1647, 12), 1541 => to_unsigned(1732, 12), 1542 => to_unsigned(1568, 12), 1543 => to_unsigned(1740, 12), 1544 => to_unsigned(2021, 12), 1545 => to_unsigned(1621, 12), 1546 => to_unsigned(1964, 12), 1547 => to_unsigned(2448, 12), 1548 => to_unsigned(2137, 12), 1549 => to_unsigned(2239, 12), 1550 => to_unsigned(1895, 12), 1551 => to_unsigned(2588, 12), 1552 => to_unsigned(2253, 12), 1553 => to_unsigned(2460, 12), 1554 => to_unsigned(1691, 12), 1555 => to_unsigned(1900, 12), 1556 => to_unsigned(1902, 12), 1557 => to_unsigned(1793, 12), 1558 => to_unsigned(1829, 12), 1559 => to_unsigned(2187, 12), 1560 => to_unsigned(1920, 12), 1561 => to_unsigned(1819, 12), 1562 => to_unsigned(2514, 12), 1563 => to_unsigned(2043, 12), 1564 => to_unsigned(2114, 12), 1565 => to_unsigned(2617, 12), 1566 => to_unsigned(1451, 12), 1567 => to_unsigned(1938, 12), 1568 => to_unsigned(2468, 12), 1569 => to_unsigned(2341, 12), 1570 => to_unsigned(2502, 12), 1571 => to_unsigned(1797, 12), 1572 => to_unsigned(1830, 12), 1573 => to_unsigned(2468, 12), 1574 => to_unsigned(2048, 12), 1575 => to_unsigned(2448, 12), 1576 => to_unsigned(2323, 12), 1577 => to_unsigned(1792, 12), 1578 => to_unsigned(2673, 12), 1579 => to_unsigned(2146, 12), 1580 => to_unsigned(1740, 12), 1581 => to_unsigned(2113, 12), 1582 => to_unsigned(1389, 12), 1583 => to_unsigned(2610, 12), 1584 => to_unsigned(1507, 12), 1585 => to_unsigned(1316, 12), 1586 => to_unsigned(2833, 12), 1587 => to_unsigned(1848, 12), 1588 => to_unsigned(1947, 12), 1589 => to_unsigned(1870, 12), 1590 => to_unsigned(2132, 12), 1591 => to_unsigned(1424, 12), 1592 => to_unsigned(2795, 12), 1593 => to_unsigned(2046, 12), 1594 => to_unsigned(1988, 12), 1595 => to_unsigned(2149, 12), 1596 => to_unsigned(1991, 12), 1597 => to_unsigned(1760, 12), 1598 => to_unsigned(1769, 12), 1599 => to_unsigned(1913, 12), 1600 => to_unsigned(2288, 12), 1601 => to_unsigned(1724, 12), 1602 => to_unsigned(2455, 12), 1603 => to_unsigned(1745, 12), 1604 => to_unsigned(1931, 12), 1605 => to_unsigned(2146, 12), 1606 => to_unsigned(2385, 12), 1607 => to_unsigned(1813, 12), 1608 => to_unsigned(1974, 12), 1609 => to_unsigned(2196, 12), 1610 => to_unsigned(1729, 12), 1611 => to_unsigned(2715, 12), 1612 => to_unsigned(1534, 12), 1613 => to_unsigned(2579, 12), 1614 => to_unsigned(1839, 12), 1615 => to_unsigned(2017, 12), 1616 => to_unsigned(1911, 12), 1617 => to_unsigned(2572, 12), 1618 => to_unsigned(2024, 12), 1619 => to_unsigned(2201, 12), 1620 => to_unsigned(1866, 12), 1621 => to_unsigned(1623, 12), 1622 => to_unsigned(1677, 12), 1623 => to_unsigned(1016, 12), 1624 => to_unsigned(1821, 12), 1625 => to_unsigned(1611, 12), 1626 => to_unsigned(2084, 12), 1627 => to_unsigned(2220, 12), 1628 => to_unsigned(2512, 12), 1629 => to_unsigned(1850, 12), 1630 => to_unsigned(2517, 12), 1631 => to_unsigned(2209, 12), 1632 => to_unsigned(2067, 12), 1633 => to_unsigned(1963, 12), 1634 => to_unsigned(1641, 12), 1635 => to_unsigned(2560, 12), 1636 => to_unsigned(1714, 12), 1637 => to_unsigned(2063, 12), 1638 => to_unsigned(1357, 12), 1639 => to_unsigned(2298, 12), 1640 => to_unsigned(2477, 12), 1641 => to_unsigned(2274, 12), 1642 => to_unsigned(1224, 12), 1643 => to_unsigned(2050, 12), 1644 => to_unsigned(1627, 12), 1645 => to_unsigned(2004, 12), 1646 => to_unsigned(2320, 12), 1647 => to_unsigned(1824, 12), 1648 => to_unsigned(1845, 12), 1649 => to_unsigned(2052, 12), 1650 => to_unsigned(2312, 12), 1651 => to_unsigned(2226, 12), 1652 => to_unsigned(1739, 12), 1653 => to_unsigned(2084, 12), 1654 => to_unsigned(1957, 12), 1655 => to_unsigned(1353, 12), 1656 => to_unsigned(2275, 12), 1657 => to_unsigned(1905, 12), 1658 => to_unsigned(2285, 12), 1659 => to_unsigned(2162, 12), 1660 => to_unsigned(1826, 12), 1661 => to_unsigned(2974, 12), 1662 => to_unsigned(2469, 12), 1663 => to_unsigned(1845, 12), 1664 => to_unsigned(1709, 12), 1665 => to_unsigned(1592, 12), 1666 => to_unsigned(2101, 12), 1667 => to_unsigned(2913, 12), 1668 => to_unsigned(1872, 12), 1669 => to_unsigned(1297, 12), 1670 => to_unsigned(2518, 12), 1671 => to_unsigned(1218, 12), 1672 => to_unsigned(2324, 12), 1673 => to_unsigned(2368, 12), 1674 => to_unsigned(1904, 12), 1675 => to_unsigned(2271, 12), 1676 => to_unsigned(2180, 12), 1677 => to_unsigned(2270, 12), 1678 => to_unsigned(2153, 12), 1679 => to_unsigned(2066, 12), 1680 => to_unsigned(1727, 12), 1681 => to_unsigned(2278, 12), 1682 => to_unsigned(2812, 12), 1683 => to_unsigned(1736, 12), 1684 => to_unsigned(1980, 12), 1685 => to_unsigned(1628, 12), 1686 => to_unsigned(1932, 12), 1687 => to_unsigned(1963, 12), 1688 => to_unsigned(1159, 12), 1689 => to_unsigned(1709, 12), 1690 => to_unsigned(2218, 12), 1691 => to_unsigned(2496, 12), 1692 => to_unsigned(1937, 12), 1693 => to_unsigned(2656, 12), 1694 => to_unsigned(1526, 12), 1695 => to_unsigned(1946, 12), 1696 => to_unsigned(1766, 12), 1697 => to_unsigned(2367, 12), 1698 => to_unsigned(2902, 12), 1699 => to_unsigned(2174, 12), 1700 => to_unsigned(2383, 12), 1701 => to_unsigned(2053, 12), 1702 => to_unsigned(2183, 12), 1703 => to_unsigned(2417, 12), 1704 => to_unsigned(2844, 12), 1705 => to_unsigned(2045, 12), 1706 => to_unsigned(1726, 12), 1707 => to_unsigned(2384, 12), 1708 => to_unsigned(2566, 12), 1709 => to_unsigned(1992, 12), 1710 => to_unsigned(2247, 12), 1711 => to_unsigned(1851, 12), 1712 => to_unsigned(1509, 12), 1713 => to_unsigned(2172, 12), 1714 => to_unsigned(2301, 12), 1715 => to_unsigned(2219, 12), 1716 => to_unsigned(2046, 12), 1717 => to_unsigned(2205, 12), 1718 => to_unsigned(1610, 12), 1719 => to_unsigned(2031, 12), 1720 => to_unsigned(2285, 12), 1721 => to_unsigned(1987, 12), 1722 => to_unsigned(2677, 12), 1723 => to_unsigned(2030, 12), 1724 => to_unsigned(2358, 12), 1725 => to_unsigned(2452, 12), 1726 => to_unsigned(2145, 12), 1727 => to_unsigned(1444, 12), 1728 => to_unsigned(2465, 12), 1729 => to_unsigned(1647, 12), 1730 => to_unsigned(973, 12), 1731 => to_unsigned(1906, 12), 1732 => to_unsigned(2641, 12), 1733 => to_unsigned(1727, 12), 1734 => to_unsigned(2471, 12), 1735 => to_unsigned(2478, 12), 1736 => to_unsigned(1674, 12), 1737 => to_unsigned(1978, 12), 1738 => to_unsigned(2016, 12), 1739 => to_unsigned(1958, 12), 1740 => to_unsigned(1847, 12), 1741 => to_unsigned(2600, 12), 1742 => to_unsigned(1487, 12), 1743 => to_unsigned(2193, 12), 1744 => to_unsigned(1394, 12), 1745 => to_unsigned(2412, 12), 1746 => to_unsigned(1701, 12), 1747 => to_unsigned(2163, 12), 1748 => to_unsigned(2227, 12), 1749 => to_unsigned(2202, 12), 1750 => to_unsigned(1959, 12), 1751 => to_unsigned(2046, 12), 1752 => to_unsigned(1998, 12), 1753 => to_unsigned(2881, 12), 1754 => to_unsigned(1893, 12), 1755 => to_unsigned(2743, 12), 1756 => to_unsigned(2096, 12), 1757 => to_unsigned(2090, 12), 1758 => to_unsigned(2685, 12), 1759 => to_unsigned(1847, 12), 1760 => to_unsigned(1451, 12), 1761 => to_unsigned(1721, 12), 1762 => to_unsigned(2282, 12), 1763 => to_unsigned(1983, 12), 1764 => to_unsigned(1593, 12), 1765 => to_unsigned(2328, 12), 1766 => to_unsigned(2235, 12), 1767 => to_unsigned(2160, 12), 1768 => to_unsigned(3126, 12), 1769 => to_unsigned(1634, 12), 1770 => to_unsigned(1536, 12), 1771 => to_unsigned(1832, 12), 1772 => to_unsigned(3135, 12), 1773 => to_unsigned(2038, 12), 1774 => to_unsigned(2702, 12), 1775 => to_unsigned(1820, 12), 1776 => to_unsigned(1738, 12), 1777 => to_unsigned(2059, 12), 1778 => to_unsigned(1989, 12), 1779 => to_unsigned(2144, 12), 1780 => to_unsigned(2122, 12), 1781 => to_unsigned(2568, 12), 1782 => to_unsigned(1972, 12), 1783 => to_unsigned(1598, 12), 1784 => to_unsigned(2169, 12), 1785 => to_unsigned(2319, 12), 1786 => to_unsigned(2036, 12), 1787 => to_unsigned(1714, 12), 1788 => to_unsigned(1852, 12), 1789 => to_unsigned(2352, 12), 1790 => to_unsigned(2509, 12), 1791 => to_unsigned(1920, 12), 1792 => to_unsigned(2237, 12), 1793 => to_unsigned(2066, 12), 1794 => to_unsigned(1659, 12), 1795 => to_unsigned(2136, 12), 1796 => to_unsigned(2008, 12), 1797 => to_unsigned(2225, 12), 1798 => to_unsigned(1832, 12), 1799 => to_unsigned(2213, 12), 1800 => to_unsigned(2747, 12), 1801 => to_unsigned(2009, 12), 1802 => to_unsigned(2209, 12), 1803 => to_unsigned(1304, 12), 1804 => to_unsigned(2744, 12), 1805 => to_unsigned(1928, 12), 1806 => to_unsigned(2138, 12), 1807 => to_unsigned(1824, 12), 1808 => to_unsigned(2136, 12), 1809 => to_unsigned(1749, 12), 1810 => to_unsigned(2620, 12), 1811 => to_unsigned(1699, 12), 1812 => to_unsigned(2096, 12), 1813 => to_unsigned(1238, 12), 1814 => to_unsigned(2130, 12), 1815 => to_unsigned(1897, 12), 1816 => to_unsigned(2642, 12), 1817 => to_unsigned(2166, 12), 1818 => to_unsigned(2735, 12), 1819 => to_unsigned(2553, 12), 1820 => to_unsigned(2252, 12), 1821 => to_unsigned(1573, 12), 1822 => to_unsigned(1649, 12), 1823 => to_unsigned(2242, 12), 1824 => to_unsigned(2276, 12), 1825 => to_unsigned(1963, 12), 1826 => to_unsigned(1797, 12), 1827 => to_unsigned(2048, 12), 1828 => to_unsigned(1959, 12), 1829 => to_unsigned(2299, 12), 1830 => to_unsigned(1874, 12), 1831 => to_unsigned(2145, 12), 1832 => to_unsigned(2194, 12), 1833 => to_unsigned(1899, 12), 1834 => to_unsigned(1801, 12), 1835 => to_unsigned(1376, 12), 1836 => to_unsigned(2567, 12), 1837 => to_unsigned(1739, 12), 1838 => to_unsigned(2327, 12), 1839 => to_unsigned(2174, 12), 1840 => to_unsigned(2169, 12), 1841 => to_unsigned(1594, 12), 1842 => to_unsigned(2044, 12), 1843 => to_unsigned(1582, 12), 1844 => to_unsigned(2261, 12), 1845 => to_unsigned(2131, 12), 1846 => to_unsigned(1965, 12), 1847 => to_unsigned(2042, 12), 1848 => to_unsigned(1286, 12), 1849 => to_unsigned(1731, 12), 1850 => to_unsigned(1108, 12), 1851 => to_unsigned(1658, 12), 1852 => to_unsigned(1993, 12), 1853 => to_unsigned(2317, 12), 1854 => to_unsigned(2000, 12), 1855 => to_unsigned(1932, 12), 1856 => to_unsigned(2668, 12), 1857 => to_unsigned(2389, 12), 1858 => to_unsigned(1983, 12), 1859 => to_unsigned(1958, 12), 1860 => to_unsigned(1900, 12), 1861 => to_unsigned(2243, 12), 1862 => to_unsigned(1516, 12), 1863 => to_unsigned(1810, 12), 1864 => to_unsigned(2175, 12), 1865 => to_unsigned(2541, 12), 1866 => to_unsigned(2020, 12), 1867 => to_unsigned(2500, 12), 1868 => to_unsigned(2022, 12), 1869 => to_unsigned(1832, 12), 1870 => to_unsigned(1574, 12), 1871 => to_unsigned(1905, 12), 1872 => to_unsigned(1839, 12), 1873 => to_unsigned(1507, 12), 1874 => to_unsigned(1588, 12), 1875 => to_unsigned(1906, 12), 1876 => to_unsigned(2327, 12), 1877 => to_unsigned(2257, 12), 1878 => to_unsigned(1699, 12), 1879 => to_unsigned(1734, 12), 1880 => to_unsigned(2080, 12), 1881 => to_unsigned(1579, 12), 1882 => to_unsigned(2189, 12), 1883 => to_unsigned(1344, 12), 1884 => to_unsigned(2057, 12), 1885 => to_unsigned(1847, 12), 1886 => to_unsigned(2492, 12), 1887 => to_unsigned(1741, 12), 1888 => to_unsigned(1627, 12), 1889 => to_unsigned(2195, 12), 1890 => to_unsigned(1766, 12), 1891 => to_unsigned(2707, 12), 1892 => to_unsigned(2492, 12), 1893 => to_unsigned(1895, 12), 1894 => to_unsigned(1803, 12), 1895 => to_unsigned(1608, 12), 1896 => to_unsigned(1839, 12), 1897 => to_unsigned(2156, 12), 1898 => to_unsigned(1995, 12), 1899 => to_unsigned(2308, 12), 1900 => to_unsigned(2218, 12), 1901 => to_unsigned(2121, 12), 1902 => to_unsigned(2011, 12), 1903 => to_unsigned(2189, 12), 1904 => to_unsigned(2246, 12), 1905 => to_unsigned(2394, 12), 1906 => to_unsigned(2117, 12), 1907 => to_unsigned(2358, 12), 1908 => to_unsigned(2364, 12), 1909 => to_unsigned(2889, 12), 1910 => to_unsigned(2194, 12), 1911 => to_unsigned(2550, 12), 1912 => to_unsigned(2049, 12), 1913 => to_unsigned(1595, 12), 1914 => to_unsigned(2381, 12), 1915 => to_unsigned(2343, 12), 1916 => to_unsigned(1714, 12), 1917 => to_unsigned(2618, 12), 1918 => to_unsigned(2163, 12), 1919 => to_unsigned(2519, 12), 1920 => to_unsigned(1604, 12), 1921 => to_unsigned(1955, 12), 1922 => to_unsigned(1819, 12), 1923 => to_unsigned(2563, 12), 1924 => to_unsigned(2261, 12), 1925 => to_unsigned(1799, 12), 1926 => to_unsigned(2352, 12), 1927 => to_unsigned(2456, 12), 1928 => to_unsigned(1655, 12), 1929 => to_unsigned(1499, 12), 1930 => to_unsigned(1770, 12), 1931 => to_unsigned(2016, 12), 1932 => to_unsigned(1735, 12), 1933 => to_unsigned(1805, 12), 1934 => to_unsigned(1970, 12), 1935 => to_unsigned(2662, 12), 1936 => to_unsigned(2095, 12), 1937 => to_unsigned(2186, 12), 1938 => to_unsigned(1626, 12), 1939 => to_unsigned(1971, 12), 1940 => to_unsigned(1578, 12), 1941 => to_unsigned(1487, 12), 1942 => to_unsigned(1980, 12), 1943 => to_unsigned(1619, 12), 1944 => to_unsigned(1900, 12), 1945 => to_unsigned(2268, 12), 1946 => to_unsigned(2219, 12), 1947 => to_unsigned(1779, 12), 1948 => to_unsigned(2518, 12), 1949 => to_unsigned(1880, 12), 1950 => to_unsigned(2008, 12), 1951 => to_unsigned(1252, 12), 1952 => to_unsigned(2599, 12), 1953 => to_unsigned(1868, 12), 1954 => to_unsigned(1901, 12), 1955 => to_unsigned(1582, 12), 1956 => to_unsigned(2085, 12), 1957 => to_unsigned(2110, 12), 1958 => to_unsigned(1956, 12), 1959 => to_unsigned(1906, 12), 1960 => to_unsigned(1599, 12), 1961 => to_unsigned(2158, 12), 1962 => to_unsigned(1834, 12), 1963 => to_unsigned(2113, 12), 1964 => to_unsigned(2107, 12), 1965 => to_unsigned(1997, 12), 1966 => to_unsigned(1621, 12), 1967 => to_unsigned(1690, 12), 1968 => to_unsigned(1635, 12), 1969 => to_unsigned(2525, 12), 1970 => to_unsigned(2332, 12), 1971 => to_unsigned(2052, 12), 1972 => to_unsigned(2087, 12), 1973 => to_unsigned(1922, 12), 1974 => to_unsigned(2205, 12), 1975 => to_unsigned(1618, 12), 1976 => to_unsigned(1536, 12), 1977 => to_unsigned(2134, 12), 1978 => to_unsigned(1822, 12), 1979 => to_unsigned(2601, 12), 1980 => to_unsigned(2163, 12), 1981 => to_unsigned(2121, 12), 1982 => to_unsigned(2261, 12), 1983 => to_unsigned(1595, 12), 1984 => to_unsigned(2153, 12), 1985 => to_unsigned(1892, 12), 1986 => to_unsigned(1635, 12), 1987 => to_unsigned(2390, 12), 1988 => to_unsigned(1691, 12), 1989 => to_unsigned(1921, 12), 1990 => to_unsigned(2171, 12), 1991 => to_unsigned(1757, 12), 1992 => to_unsigned(1681, 12), 1993 => to_unsigned(1957, 12), 1994 => to_unsigned(1427, 12), 1995 => to_unsigned(2054, 12), 1996 => to_unsigned(1530, 12), 1997 => to_unsigned(1819, 12), 1998 => to_unsigned(2071, 12), 1999 => to_unsigned(1857, 12), 2000 => to_unsigned(1474, 12), 2001 => to_unsigned(2192, 12), 2002 => to_unsigned(1445, 12), 2003 => to_unsigned(2282, 12), 2004 => to_unsigned(2001, 12), 2005 => to_unsigned(2437, 12), 2006 => to_unsigned(2272, 12), 2007 => to_unsigned(2110, 12), 2008 => to_unsigned(2134, 12), 2009 => to_unsigned(2030, 12), 2010 => to_unsigned(1207, 12), 2011 => to_unsigned(2077, 12), 2012 => to_unsigned(2197, 12), 2013 => to_unsigned(1967, 12), 2014 => to_unsigned(2049, 12), 2015 => to_unsigned(2121, 12), 2016 => to_unsigned(2153, 12), 2017 => to_unsigned(2459, 12), 2018 => to_unsigned(1977, 12), 2019 => to_unsigned(1641, 12), 2020 => to_unsigned(2075, 12), 2021 => to_unsigned(1391, 12), 2022 => to_unsigned(2086, 12), 2023 => to_unsigned(1924, 12), 2024 => to_unsigned(2460, 12), 2025 => to_unsigned(1653, 12), 2026 => to_unsigned(2319, 12), 2027 => to_unsigned(2698, 12), 2028 => to_unsigned(2581, 12), 2029 => to_unsigned(2462, 12), 2030 => to_unsigned(2690, 12), 2031 => to_unsigned(2042, 12), 2032 => to_unsigned(2223, 12), 2033 => to_unsigned(1787, 12), 2034 => to_unsigned(2097, 12), 2035 => to_unsigned(1995, 12), 2036 => to_unsigned(2136, 12), 2037 => to_unsigned(1541, 12), 2038 => to_unsigned(2041, 12), 2039 => to_unsigned(2057, 12), 2040 => to_unsigned(2072, 12), 2041 => to_unsigned(2004, 12), 2042 => to_unsigned(1920, 12), 2043 => to_unsigned(2102, 12), 2044 => to_unsigned(2012, 12), 2045 => to_unsigned(1839, 12), 2046 => to_unsigned(2472, 12), 2047 => to_unsigned(2240, 12)),
        1 => (0 => to_unsigned(1531, 12), 1 => to_unsigned(2102, 12), 2 => to_unsigned(1927, 12), 3 => to_unsigned(2651, 12), 4 => to_unsigned(2410, 12), 5 => to_unsigned(1658, 12), 6 => to_unsigned(2642, 12), 7 => to_unsigned(2424, 12), 8 => to_unsigned(2169, 12), 9 => to_unsigned(1929, 12), 10 => to_unsigned(1565, 12), 11 => to_unsigned(1874, 12), 12 => to_unsigned(1261, 12), 13 => to_unsigned(2258, 12), 14 => to_unsigned(2082, 12), 15 => to_unsigned(1983, 12), 16 => to_unsigned(2588, 12), 17 => to_unsigned(2198, 12), 18 => to_unsigned(2647, 12), 19 => to_unsigned(2525, 12), 20 => to_unsigned(1641, 12), 21 => to_unsigned(1931, 12), 22 => to_unsigned(2340, 12), 23 => to_unsigned(2434, 12), 24 => to_unsigned(2933, 12), 25 => to_unsigned(2734, 12), 26 => to_unsigned(1867, 12), 27 => to_unsigned(1483, 12), 28 => to_unsigned(2259, 12), 29 => to_unsigned(1503, 12), 30 => to_unsigned(1976, 12), 31 => to_unsigned(1435, 12), 32 => to_unsigned(2112, 12), 33 => to_unsigned(1842, 12), 34 => to_unsigned(1386, 12), 35 => to_unsigned(2154, 12), 36 => to_unsigned(3102, 12), 37 => to_unsigned(1753, 12), 38 => to_unsigned(2740, 12), 39 => to_unsigned(2237, 12), 40 => to_unsigned(1832, 12), 41 => to_unsigned(2779, 12), 42 => to_unsigned(2199, 12), 43 => to_unsigned(2189, 12), 44 => to_unsigned(2154, 12), 45 => to_unsigned(2985, 12), 46 => to_unsigned(1976, 12), 47 => to_unsigned(2725, 12), 48 => to_unsigned(1652, 12), 49 => to_unsigned(1821, 12), 50 => to_unsigned(2281, 12), 51 => to_unsigned(2593, 12), 52 => to_unsigned(1945, 12), 53 => to_unsigned(1825, 12), 54 => to_unsigned(1801, 12), 55 => to_unsigned(2856, 12), 56 => to_unsigned(2361, 12), 57 => to_unsigned(2082, 12), 58 => to_unsigned(1696, 12), 59 => to_unsigned(1592, 12), 60 => to_unsigned(1246, 12), 61 => to_unsigned(2181, 12), 62 => to_unsigned(1281, 12), 63 => to_unsigned(1530, 12), 64 => to_unsigned(2732, 12), 65 => to_unsigned(1786, 12), 66 => to_unsigned(1826, 12), 67 => to_unsigned(1584, 12), 68 => to_unsigned(2154, 12), 69 => to_unsigned(2712, 12), 70 => to_unsigned(2397, 12), 71 => to_unsigned(1832, 12), 72 => to_unsigned(2481, 12), 73 => to_unsigned(1783, 12), 74 => to_unsigned(2416, 12), 75 => to_unsigned(2473, 12), 76 => to_unsigned(2229, 12), 77 => to_unsigned(2066, 12), 78 => to_unsigned(2457, 12), 79 => to_unsigned(2034, 12), 80 => to_unsigned(2171, 12), 81 => to_unsigned(2326, 12), 82 => to_unsigned(1858, 12), 83 => to_unsigned(2593, 12), 84 => to_unsigned(2009, 12), 85 => to_unsigned(1657, 12), 86 => to_unsigned(1855, 12), 87 => to_unsigned(1320, 12), 88 => to_unsigned(2165, 12), 89 => to_unsigned(1593, 12), 90 => to_unsigned(2066, 12), 91 => to_unsigned(1702, 12), 92 => to_unsigned(2236, 12), 93 => to_unsigned(1744, 12), 94 => to_unsigned(1729, 12), 95 => to_unsigned(2658, 12), 96 => to_unsigned(2140, 12), 97 => to_unsigned(1981, 12), 98 => to_unsigned(2242, 12), 99 => to_unsigned(1205, 12), 100 => to_unsigned(2066, 12), 101 => to_unsigned(2188, 12), 102 => to_unsigned(1809, 12), 103 => to_unsigned(2424, 12), 104 => to_unsigned(2654, 12), 105 => to_unsigned(2480, 12), 106 => to_unsigned(2296, 12), 107 => to_unsigned(1689, 12), 108 => to_unsigned(2205, 12), 109 => to_unsigned(2519, 12), 110 => to_unsigned(2026, 12), 111 => to_unsigned(1774, 12), 112 => to_unsigned(1384, 12), 113 => to_unsigned(2168, 12), 114 => to_unsigned(1079, 12), 115 => to_unsigned(2167, 12), 116 => to_unsigned(2436, 12), 117 => to_unsigned(2194, 12), 118 => to_unsigned(2177, 12), 119 => to_unsigned(1591, 12), 120 => to_unsigned(2404, 12), 121 => to_unsigned(2226, 12), 122 => to_unsigned(1351, 12), 123 => to_unsigned(2045, 12), 124 => to_unsigned(1370, 12), 125 => to_unsigned(1866, 12), 126 => to_unsigned(2075, 12), 127 => to_unsigned(2340, 12), 128 => to_unsigned(2071, 12), 129 => to_unsigned(2539, 12), 130 => to_unsigned(1482, 12), 131 => to_unsigned(2385, 12), 132 => to_unsigned(1617, 12), 133 => to_unsigned(2318, 12), 134 => to_unsigned(2902, 12), 135 => to_unsigned(1577, 12), 136 => to_unsigned(2232, 12), 137 => to_unsigned(2473, 12), 138 => to_unsigned(2306, 12), 139 => to_unsigned(2177, 12), 140 => to_unsigned(1464, 12), 141 => to_unsigned(1961, 12), 142 => to_unsigned(2305, 12), 143 => to_unsigned(2228, 12), 144 => to_unsigned(2835, 12), 145 => to_unsigned(2594, 12), 146 => to_unsigned(2466, 12), 147 => to_unsigned(2341, 12), 148 => to_unsigned(2338, 12), 149 => to_unsigned(1541, 12), 150 => to_unsigned(1808, 12), 151 => to_unsigned(2570, 12), 152 => to_unsigned(2166, 12), 153 => to_unsigned(1846, 12), 154 => to_unsigned(2097, 12), 155 => to_unsigned(1789, 12), 156 => to_unsigned(1955, 12), 157 => to_unsigned(2253, 12), 158 => to_unsigned(1507, 12), 159 => to_unsigned(2090, 12), 160 => to_unsigned(1395, 12), 161 => to_unsigned(1449, 12), 162 => to_unsigned(2230, 12), 163 => to_unsigned(1599, 12), 164 => to_unsigned(2023, 12), 165 => to_unsigned(1520, 12), 166 => to_unsigned(1650, 12), 167 => to_unsigned(2149, 12), 168 => to_unsigned(2184, 12), 169 => to_unsigned(1575, 12), 170 => to_unsigned(1327, 12), 171 => to_unsigned(1693, 12), 172 => to_unsigned(1943, 12), 173 => to_unsigned(2092, 12), 174 => to_unsigned(2018, 12), 175 => to_unsigned(2077, 12), 176 => to_unsigned(2258, 12), 177 => to_unsigned(2029, 12), 178 => to_unsigned(1329, 12), 179 => to_unsigned(2370, 12), 180 => to_unsigned(2477, 12), 181 => to_unsigned(1753, 12), 182 => to_unsigned(2278, 12), 183 => to_unsigned(1854, 12), 184 => to_unsigned(1689, 12), 185 => to_unsigned(2171, 12), 186 => to_unsigned(1548, 12), 187 => to_unsigned(2115, 12), 188 => to_unsigned(2196, 12), 189 => to_unsigned(1534, 12), 190 => to_unsigned(2098, 12), 191 => to_unsigned(1975, 12), 192 => to_unsigned(2413, 12), 193 => to_unsigned(1920, 12), 194 => to_unsigned(1431, 12), 195 => to_unsigned(2752, 12), 196 => to_unsigned(1675, 12), 197 => to_unsigned(1601, 12), 198 => to_unsigned(2273, 12), 199 => to_unsigned(2429, 12), 200 => to_unsigned(2527, 12), 201 => to_unsigned(1999, 12), 202 => to_unsigned(2123, 12), 203 => to_unsigned(1884, 12), 204 => to_unsigned(1920, 12), 205 => to_unsigned(2539, 12), 206 => to_unsigned(2534, 12), 207 => to_unsigned(2390, 12), 208 => to_unsigned(2155, 12), 209 => to_unsigned(2323, 12), 210 => to_unsigned(1964, 12), 211 => to_unsigned(1480, 12), 212 => to_unsigned(2334, 12), 213 => to_unsigned(1815, 12), 214 => to_unsigned(2048, 12), 215 => to_unsigned(2013, 12), 216 => to_unsigned(1602, 12), 217 => to_unsigned(2478, 12), 218 => to_unsigned(1668, 12), 219 => to_unsigned(1834, 12), 220 => to_unsigned(1580, 12), 221 => to_unsigned(1851, 12), 222 => to_unsigned(2049, 12), 223 => to_unsigned(1771, 12), 224 => to_unsigned(2159, 12), 225 => to_unsigned(1701, 12), 226 => to_unsigned(1839, 12), 227 => to_unsigned(1801, 12), 228 => to_unsigned(2506, 12), 229 => to_unsigned(3021, 12), 230 => to_unsigned(1998, 12), 231 => to_unsigned(2035, 12), 232 => to_unsigned(2414, 12), 233 => to_unsigned(1778, 12), 234 => to_unsigned(1735, 12), 235 => to_unsigned(1907, 12), 236 => to_unsigned(1208, 12), 237 => to_unsigned(1854, 12), 238 => to_unsigned(2232, 12), 239 => to_unsigned(2243, 12), 240 => to_unsigned(1948, 12), 241 => to_unsigned(1703, 12), 242 => to_unsigned(1914, 12), 243 => to_unsigned(1498, 12), 244 => to_unsigned(2219, 12), 245 => to_unsigned(1242, 12), 246 => to_unsigned(1937, 12), 247 => to_unsigned(2564, 12), 248 => to_unsigned(2645, 12), 249 => to_unsigned(1593, 12), 250 => to_unsigned(1857, 12), 251 => to_unsigned(1753, 12), 252 => to_unsigned(2332, 12), 253 => to_unsigned(2235, 12), 254 => to_unsigned(2655, 12), 255 => to_unsigned(2238, 12), 256 => to_unsigned(2077, 12), 257 => to_unsigned(2373, 12), 258 => to_unsigned(2052, 12), 259 => to_unsigned(2348, 12), 260 => to_unsigned(2207, 12), 261 => to_unsigned(1926, 12), 262 => to_unsigned(2397, 12), 263 => to_unsigned(1876, 12), 264 => to_unsigned(2417, 12), 265 => to_unsigned(2245, 12), 266 => to_unsigned(1805, 12), 267 => to_unsigned(1580, 12), 268 => to_unsigned(2233, 12), 269 => to_unsigned(2169, 12), 270 => to_unsigned(2000, 12), 271 => to_unsigned(1652, 12), 272 => to_unsigned(1511, 12), 273 => to_unsigned(1485, 12), 274 => to_unsigned(919, 12), 275 => to_unsigned(2117, 12), 276 => to_unsigned(1999, 12), 277 => to_unsigned(1435, 12), 278 => to_unsigned(2225, 12), 279 => to_unsigned(2516, 12), 280 => to_unsigned(2696, 12), 281 => to_unsigned(1775, 12), 282 => to_unsigned(2156, 12), 283 => to_unsigned(2148, 12), 284 => to_unsigned(2469, 12), 285 => to_unsigned(2182, 12), 286 => to_unsigned(1987, 12), 287 => to_unsigned(2341, 12), 288 => to_unsigned(1658, 12), 289 => to_unsigned(2513, 12), 290 => to_unsigned(2241, 12), 291 => to_unsigned(2181, 12), 292 => to_unsigned(1936, 12), 293 => to_unsigned(2277, 12), 294 => to_unsigned(2252, 12), 295 => to_unsigned(2115, 12), 296 => to_unsigned(2092, 12), 297 => to_unsigned(2384, 12), 298 => to_unsigned(1825, 12), 299 => to_unsigned(2118, 12), 300 => to_unsigned(1486, 12), 301 => to_unsigned(1876, 12), 302 => to_unsigned(1616, 12), 303 => to_unsigned(2175, 12), 304 => to_unsigned(2379, 12), 305 => to_unsigned(1952, 12), 306 => to_unsigned(2425, 12), 307 => to_unsigned(1852, 12), 308 => to_unsigned(1675, 12), 309 => to_unsigned(1904, 12), 310 => to_unsigned(1703, 12), 311 => to_unsigned(1649, 12), 312 => to_unsigned(1356, 12), 313 => to_unsigned(2241, 12), 314 => to_unsigned(1692, 12), 315 => to_unsigned(2097, 12), 316 => to_unsigned(1942, 12), 317 => to_unsigned(2132, 12), 318 => to_unsigned(1650, 12), 319 => to_unsigned(2309, 12), 320 => to_unsigned(2298, 12), 321 => to_unsigned(2288, 12), 322 => to_unsigned(1714, 12), 323 => to_unsigned(2095, 12), 324 => to_unsigned(1954, 12), 325 => to_unsigned(2142, 12), 326 => to_unsigned(2035, 12), 327 => to_unsigned(2625, 12), 328 => to_unsigned(2458, 12), 329 => to_unsigned(2235, 12), 330 => to_unsigned(2298, 12), 331 => to_unsigned(1921, 12), 332 => to_unsigned(1668, 12), 333 => to_unsigned(2238, 12), 334 => to_unsigned(2320, 12), 335 => to_unsigned(1778, 12), 336 => to_unsigned(2419, 12), 337 => to_unsigned(1968, 12), 338 => to_unsigned(2519, 12), 339 => to_unsigned(2179, 12), 340 => to_unsigned(2695, 12), 341 => to_unsigned(1781, 12), 342 => to_unsigned(1717, 12), 343 => to_unsigned(2079, 12), 344 => to_unsigned(1808, 12), 345 => to_unsigned(1531, 12), 346 => to_unsigned(1897, 12), 347 => to_unsigned(2286, 12), 348 => to_unsigned(3084, 12), 349 => to_unsigned(1531, 12), 350 => to_unsigned(2152, 12), 351 => to_unsigned(2436, 12), 352 => to_unsigned(2376, 12), 353 => to_unsigned(2175, 12), 354 => to_unsigned(2463, 12), 355 => to_unsigned(2255, 12), 356 => to_unsigned(2017, 12), 357 => to_unsigned(2291, 12), 358 => to_unsigned(2007, 12), 359 => to_unsigned(2776, 12), 360 => to_unsigned(2121, 12), 361 => to_unsigned(1689, 12), 362 => to_unsigned(2048, 12), 363 => to_unsigned(2339, 12), 364 => to_unsigned(1398, 12), 365 => to_unsigned(1966, 12), 366 => to_unsigned(3111, 12), 367 => to_unsigned(2294, 12), 368 => to_unsigned(2228, 12), 369 => to_unsigned(2167, 12), 370 => to_unsigned(2894, 12), 371 => to_unsigned(1642, 12), 372 => to_unsigned(1534, 12), 373 => to_unsigned(1328, 12), 374 => to_unsigned(2406, 12), 375 => to_unsigned(1813, 12), 376 => to_unsigned(2344, 12), 377 => to_unsigned(2532, 12), 378 => to_unsigned(2515, 12), 379 => to_unsigned(1863, 12), 380 => to_unsigned(2739, 12), 381 => to_unsigned(1669, 12), 382 => to_unsigned(1756, 12), 383 => to_unsigned(2552, 12), 384 => to_unsigned(1140, 12), 385 => to_unsigned(1771, 12), 386 => to_unsigned(1799, 12), 387 => to_unsigned(2115, 12), 388 => to_unsigned(2000, 12), 389 => to_unsigned(2319, 12), 390 => to_unsigned(2643, 12), 391 => to_unsigned(2415, 12), 392 => to_unsigned(1651, 12), 393 => to_unsigned(1332, 12), 394 => to_unsigned(1683, 12), 395 => to_unsigned(1347, 12), 396 => to_unsigned(1909, 12), 397 => to_unsigned(1991, 12), 398 => to_unsigned(1500, 12), 399 => to_unsigned(1605, 12), 400 => to_unsigned(1891, 12), 401 => to_unsigned(2203, 12), 402 => to_unsigned(2454, 12), 403 => to_unsigned(2571, 12), 404 => to_unsigned(2153, 12), 405 => to_unsigned(2715, 12), 406 => to_unsigned(2272, 12), 407 => to_unsigned(1558, 12), 408 => to_unsigned(1974, 12), 409 => to_unsigned(1965, 12), 410 => to_unsigned(1382, 12), 411 => to_unsigned(1570, 12), 412 => to_unsigned(2136, 12), 413 => to_unsigned(1952, 12), 414 => to_unsigned(1441, 12), 415 => to_unsigned(1344, 12), 416 => to_unsigned(2099, 12), 417 => to_unsigned(1961, 12), 418 => to_unsigned(2542, 12), 419 => to_unsigned(1285, 12), 420 => to_unsigned(2434, 12), 421 => to_unsigned(2795, 12), 422 => to_unsigned(1944, 12), 423 => to_unsigned(1902, 12), 424 => to_unsigned(2275, 12), 425 => to_unsigned(2157, 12), 426 => to_unsigned(1711, 12), 427 => to_unsigned(1871, 12), 428 => to_unsigned(2434, 12), 429 => to_unsigned(2344, 12), 430 => to_unsigned(1956, 12), 431 => to_unsigned(2160, 12), 432 => to_unsigned(2196, 12), 433 => to_unsigned(2652, 12), 434 => to_unsigned(2520, 12), 435 => to_unsigned(1996, 12), 436 => to_unsigned(1565, 12), 437 => to_unsigned(2293, 12), 438 => to_unsigned(2496, 12), 439 => to_unsigned(2256, 12), 440 => to_unsigned(2057, 12), 441 => to_unsigned(1868, 12), 442 => to_unsigned(1982, 12), 443 => to_unsigned(2831, 12), 444 => to_unsigned(2165, 12), 445 => to_unsigned(1753, 12), 446 => to_unsigned(1485, 12), 447 => to_unsigned(2760, 12), 448 => to_unsigned(2337, 12), 449 => to_unsigned(1967, 12), 450 => to_unsigned(2366, 12), 451 => to_unsigned(1850, 12), 452 => to_unsigned(1994, 12), 453 => to_unsigned(2183, 12), 454 => to_unsigned(2398, 12), 455 => to_unsigned(2007, 12), 456 => to_unsigned(1361, 12), 457 => to_unsigned(2074, 12), 458 => to_unsigned(2041, 12), 459 => to_unsigned(1648, 12), 460 => to_unsigned(2369, 12), 461 => to_unsigned(2118, 12), 462 => to_unsigned(1903, 12), 463 => to_unsigned(2408, 12), 464 => to_unsigned(1827, 12), 465 => to_unsigned(2084, 12), 466 => to_unsigned(2269, 12), 467 => to_unsigned(2331, 12), 468 => to_unsigned(2032, 12), 469 => to_unsigned(2105, 12), 470 => to_unsigned(2679, 12), 471 => to_unsigned(1310, 12), 472 => to_unsigned(1924, 12), 473 => to_unsigned(2213, 12), 474 => to_unsigned(1925, 12), 475 => to_unsigned(2206, 12), 476 => to_unsigned(1959, 12), 477 => to_unsigned(1896, 12), 478 => to_unsigned(1617, 12), 479 => to_unsigned(2332, 12), 480 => to_unsigned(2115, 12), 481 => to_unsigned(2314, 12), 482 => to_unsigned(2050, 12), 483 => to_unsigned(1192, 12), 484 => to_unsigned(2312, 12), 485 => to_unsigned(2188, 12), 486 => to_unsigned(1922, 12), 487 => to_unsigned(2052, 12), 488 => to_unsigned(1883, 12), 489 => to_unsigned(1901, 12), 490 => to_unsigned(2763, 12), 491 => to_unsigned(2022, 12), 492 => to_unsigned(1288, 12), 493 => to_unsigned(1925, 12), 494 => to_unsigned(1113, 12), 495 => to_unsigned(2111, 12), 496 => to_unsigned(2117, 12), 497 => to_unsigned(2357, 12), 498 => to_unsigned(2038, 12), 499 => to_unsigned(1780, 12), 500 => to_unsigned(2269, 12), 501 => to_unsigned(1538, 12), 502 => to_unsigned(2326, 12), 503 => to_unsigned(2193, 12), 504 => to_unsigned(1953, 12), 505 => to_unsigned(1827, 12), 506 => to_unsigned(2996, 12), 507 => to_unsigned(2684, 12), 508 => to_unsigned(2212, 12), 509 => to_unsigned(2681, 12), 510 => to_unsigned(2298, 12), 511 => to_unsigned(1790, 12), 512 => to_unsigned(1835, 12), 513 => to_unsigned(1856, 12), 514 => to_unsigned(2241, 12), 515 => to_unsigned(1838, 12), 516 => to_unsigned(1444, 12), 517 => to_unsigned(2534, 12), 518 => to_unsigned(1658, 12), 519 => to_unsigned(1747, 12), 520 => to_unsigned(1908, 12), 521 => to_unsigned(1963, 12), 522 => to_unsigned(1877, 12), 523 => to_unsigned(2341, 12), 524 => to_unsigned(2175, 12), 525 => to_unsigned(2373, 12), 526 => to_unsigned(1717, 12), 527 => to_unsigned(2262, 12), 528 => to_unsigned(2418, 12), 529 => to_unsigned(2563, 12), 530 => to_unsigned(2080, 12), 531 => to_unsigned(1768, 12), 532 => to_unsigned(2103, 12), 533 => to_unsigned(1371, 12), 534 => to_unsigned(1701, 12), 535 => to_unsigned(1947, 12), 536 => to_unsigned(1399, 12), 537 => to_unsigned(2053, 12), 538 => to_unsigned(1744, 12), 539 => to_unsigned(2223, 12), 540 => to_unsigned(2320, 12), 541 => to_unsigned(1926, 12), 542 => to_unsigned(2459, 12), 543 => to_unsigned(2240, 12), 544 => to_unsigned(1959, 12), 545 => to_unsigned(2218, 12), 546 => to_unsigned(2609, 12), 547 => to_unsigned(2311, 12), 548 => to_unsigned(2203, 12), 549 => to_unsigned(2014, 12), 550 => to_unsigned(1255, 12), 551 => to_unsigned(2063, 12), 552 => to_unsigned(1856, 12), 553 => to_unsigned(2120, 12), 554 => to_unsigned(2605, 12), 555 => to_unsigned(1919, 12), 556 => to_unsigned(1140, 12), 557 => to_unsigned(1647, 12), 558 => to_unsigned(1458, 12), 559 => to_unsigned(1845, 12), 560 => to_unsigned(1918, 12), 561 => to_unsigned(2021, 12), 562 => to_unsigned(1707, 12), 563 => to_unsigned(1297, 12), 564 => to_unsigned(2518, 12), 565 => to_unsigned(2504, 12), 566 => to_unsigned(2578, 12), 567 => to_unsigned(1940, 12), 568 => to_unsigned(1439, 12), 569 => to_unsigned(2419, 12), 570 => to_unsigned(2264, 12), 571 => to_unsigned(2009, 12), 572 => to_unsigned(1394, 12), 573 => to_unsigned(1856, 12), 574 => to_unsigned(1839, 12), 575 => to_unsigned(2690, 12), 576 => to_unsigned(1380, 12), 577 => to_unsigned(2310, 12), 578 => to_unsigned(1701, 12), 579 => to_unsigned(1914, 12), 580 => to_unsigned(2390, 12), 581 => to_unsigned(2112, 12), 582 => to_unsigned(2567, 12), 583 => to_unsigned(2152, 12), 584 => to_unsigned(2105, 12), 585 => to_unsigned(2718, 12), 586 => to_unsigned(2315, 12), 587 => to_unsigned(1893, 12), 588 => to_unsigned(1980, 12), 589 => to_unsigned(2697, 12), 590 => to_unsigned(2142, 12), 591 => to_unsigned(1558, 12), 592 => to_unsigned(1803, 12), 593 => to_unsigned(2459, 12), 594 => to_unsigned(2224, 12), 595 => to_unsigned(2309, 12), 596 => to_unsigned(2106, 12), 597 => to_unsigned(1987, 12), 598 => to_unsigned(2136, 12), 599 => to_unsigned(1726, 12), 600 => to_unsigned(2691, 12), 601 => to_unsigned(2287, 12), 602 => to_unsigned(2487, 12), 603 => to_unsigned(1956, 12), 604 => to_unsigned(3012, 12), 605 => to_unsigned(2058, 12), 606 => to_unsigned(1995, 12), 607 => to_unsigned(2438, 12), 608 => to_unsigned(2799, 12), 609 => to_unsigned(1594, 12), 610 => to_unsigned(1608, 12), 611 => to_unsigned(1708, 12), 612 => to_unsigned(2330, 12), 613 => to_unsigned(1981, 12), 614 => to_unsigned(1933, 12), 615 => to_unsigned(2376, 12), 616 => to_unsigned(1824, 12), 617 => to_unsigned(2296, 12), 618 => to_unsigned(2520, 12), 619 => to_unsigned(2035, 12), 620 => to_unsigned(2172, 12), 621 => to_unsigned(1683, 12), 622 => to_unsigned(1561, 12), 623 => to_unsigned(2202, 12), 624 => to_unsigned(1826, 12), 625 => to_unsigned(2125, 12), 626 => to_unsigned(1403, 12), 627 => to_unsigned(1792, 12), 628 => to_unsigned(2293, 12), 629 => to_unsigned(2265, 12), 630 => to_unsigned(2171, 12), 631 => to_unsigned(2677, 12), 632 => to_unsigned(2381, 12), 633 => to_unsigned(2807, 12), 634 => to_unsigned(1989, 12), 635 => to_unsigned(2670, 12), 636 => to_unsigned(1706, 12), 637 => to_unsigned(1791, 12), 638 => to_unsigned(2549, 12), 639 => to_unsigned(2251, 12), 640 => to_unsigned(2083, 12), 641 => to_unsigned(2145, 12), 642 => to_unsigned(2158, 12), 643 => to_unsigned(2231, 12), 644 => to_unsigned(2130, 12), 645 => to_unsigned(1257, 12), 646 => to_unsigned(2089, 12), 647 => to_unsigned(1760, 12), 648 => to_unsigned(2512, 12), 649 => to_unsigned(2304, 12), 650 => to_unsigned(2205, 12), 651 => to_unsigned(2818, 12), 652 => to_unsigned(1718, 12), 653 => to_unsigned(1878, 12), 654 => to_unsigned(1722, 12), 655 => to_unsigned(1174, 12), 656 => to_unsigned(2188, 12), 657 => to_unsigned(1962, 12), 658 => to_unsigned(1995, 12), 659 => to_unsigned(2062, 12), 660 => to_unsigned(2507, 12), 661 => to_unsigned(1496, 12), 662 => to_unsigned(2101, 12), 663 => to_unsigned(1699, 12), 664 => to_unsigned(1850, 12), 665 => to_unsigned(1985, 12), 666 => to_unsigned(2125, 12), 667 => to_unsigned(2122, 12), 668 => to_unsigned(2545, 12), 669 => to_unsigned(1915, 12), 670 => to_unsigned(2177, 12), 671 => to_unsigned(3051, 12), 672 => to_unsigned(1489, 12), 673 => to_unsigned(2105, 12), 674 => to_unsigned(2192, 12), 675 => to_unsigned(1672, 12), 676 => to_unsigned(1848, 12), 677 => to_unsigned(2006, 12), 678 => to_unsigned(1564, 12), 679 => to_unsigned(2217, 12), 680 => to_unsigned(2149, 12), 681 => to_unsigned(1694, 12), 682 => to_unsigned(1981, 12), 683 => to_unsigned(1750, 12), 684 => to_unsigned(2326, 12), 685 => to_unsigned(2043, 12), 686 => to_unsigned(2519, 12), 687 => to_unsigned(2335, 12), 688 => to_unsigned(2128, 12), 689 => to_unsigned(2554, 12), 690 => to_unsigned(2307, 12), 691 => to_unsigned(1909, 12), 692 => to_unsigned(1874, 12), 693 => to_unsigned(1708, 12), 694 => to_unsigned(2280, 12), 695 => to_unsigned(2228, 12), 696 => to_unsigned(1664, 12), 697 => to_unsigned(1816, 12), 698 => to_unsigned(2207, 12), 699 => to_unsigned(2296, 12), 700 => to_unsigned(1942, 12), 701 => to_unsigned(2637, 12), 702 => to_unsigned(1666, 12), 703 => to_unsigned(2020, 12), 704 => to_unsigned(2292, 12), 705 => to_unsigned(2248, 12), 706 => to_unsigned(2087, 12), 707 => to_unsigned(1840, 12), 708 => to_unsigned(1578, 12), 709 => to_unsigned(1340, 12), 710 => to_unsigned(2722, 12), 711 => to_unsigned(2040, 12), 712 => to_unsigned(1666, 12), 713 => to_unsigned(1389, 12), 714 => to_unsigned(2965, 12), 715 => to_unsigned(1497, 12), 716 => to_unsigned(3098, 12), 717 => to_unsigned(1819, 12), 718 => to_unsigned(2551, 12), 719 => to_unsigned(2146, 12), 720 => to_unsigned(1786, 12), 721 => to_unsigned(1975, 12), 722 => to_unsigned(2252, 12), 723 => to_unsigned(1847, 12), 724 => to_unsigned(2638, 12), 725 => to_unsigned(2212, 12), 726 => to_unsigned(2376, 12), 727 => to_unsigned(2353, 12), 728 => to_unsigned(2123, 12), 729 => to_unsigned(1525, 12), 730 => to_unsigned(1360, 12), 731 => to_unsigned(2160, 12), 732 => to_unsigned(2696, 12), 733 => to_unsigned(1489, 12), 734 => to_unsigned(2228, 12), 735 => to_unsigned(2269, 12), 736 => to_unsigned(1842, 12), 737 => to_unsigned(1053, 12), 738 => to_unsigned(1890, 12), 739 => to_unsigned(1878, 12), 740 => to_unsigned(2450, 12), 741 => to_unsigned(1566, 12), 742 => to_unsigned(1911, 12), 743 => to_unsigned(1975, 12), 744 => to_unsigned(1799, 12), 745 => to_unsigned(2430, 12), 746 => to_unsigned(2490, 12), 747 => to_unsigned(2578, 12), 748 => to_unsigned(2491, 12), 749 => to_unsigned(1756, 12), 750 => to_unsigned(2284, 12), 751 => to_unsigned(1724, 12), 752 => to_unsigned(2598, 12), 753 => to_unsigned(2231, 12), 754 => to_unsigned(2493, 12), 755 => to_unsigned(1817, 12), 756 => to_unsigned(1554, 12), 757 => to_unsigned(2260, 12), 758 => to_unsigned(2391, 12), 759 => to_unsigned(2192, 12), 760 => to_unsigned(1753, 12), 761 => to_unsigned(2460, 12), 762 => to_unsigned(2139, 12), 763 => to_unsigned(2154, 12), 764 => to_unsigned(1698, 12), 765 => to_unsigned(2443, 12), 766 => to_unsigned(1552, 12), 767 => to_unsigned(2135, 12), 768 => to_unsigned(1265, 12), 769 => to_unsigned(1764, 12), 770 => to_unsigned(1865, 12), 771 => to_unsigned(2364, 12), 772 => to_unsigned(3079, 12), 773 => to_unsigned(2224, 12), 774 => to_unsigned(2669, 12), 775 => to_unsigned(2101, 12), 776 => to_unsigned(1946, 12), 777 => to_unsigned(2122, 12), 778 => to_unsigned(1724, 12), 779 => to_unsigned(2081, 12), 780 => to_unsigned(2218, 12), 781 => to_unsigned(1907, 12), 782 => to_unsigned(2841, 12), 783 => to_unsigned(2198, 12), 784 => to_unsigned(2217, 12), 785 => to_unsigned(1923, 12), 786 => to_unsigned(2100, 12), 787 => to_unsigned(2384, 12), 788 => to_unsigned(1971, 12), 789 => to_unsigned(1777, 12), 790 => to_unsigned(2355, 12), 791 => to_unsigned(2186, 12), 792 => to_unsigned(1964, 12), 793 => to_unsigned(2271, 12), 794 => to_unsigned(1483, 12), 795 => to_unsigned(2315, 12), 796 => to_unsigned(1407, 12), 797 => to_unsigned(1672, 12), 798 => to_unsigned(2351, 12), 799 => to_unsigned(2494, 12), 800 => to_unsigned(2161, 12), 801 => to_unsigned(1310, 12), 802 => to_unsigned(2306, 12), 803 => to_unsigned(2013, 12), 804 => to_unsigned(2400, 12), 805 => to_unsigned(2432, 12), 806 => to_unsigned(1116, 12), 807 => to_unsigned(2228, 12), 808 => to_unsigned(1999, 12), 809 => to_unsigned(2373, 12), 810 => to_unsigned(1926, 12), 811 => to_unsigned(1993, 12), 812 => to_unsigned(1799, 12), 813 => to_unsigned(1679, 12), 814 => to_unsigned(2508, 12), 815 => to_unsigned(1649, 12), 816 => to_unsigned(2030, 12), 817 => to_unsigned(1922, 12), 818 => to_unsigned(1628, 12), 819 => to_unsigned(2457, 12), 820 => to_unsigned(2441, 12), 821 => to_unsigned(1746, 12), 822 => to_unsigned(1296, 12), 823 => to_unsigned(1825, 12), 824 => to_unsigned(1478, 12), 825 => to_unsigned(1444, 12), 826 => to_unsigned(2232, 12), 827 => to_unsigned(1663, 12), 828 => to_unsigned(1818, 12), 829 => to_unsigned(2674, 12), 830 => to_unsigned(2306, 12), 831 => to_unsigned(2614, 12), 832 => to_unsigned(2683, 12), 833 => to_unsigned(1684, 12), 834 => to_unsigned(2148, 12), 835 => to_unsigned(2124, 12), 836 => to_unsigned(1965, 12), 837 => to_unsigned(2316, 12), 838 => to_unsigned(1410, 12), 839 => to_unsigned(2104, 12), 840 => to_unsigned(2325, 12), 841 => to_unsigned(1909, 12), 842 => to_unsigned(1775, 12), 843 => to_unsigned(2022, 12), 844 => to_unsigned(2339, 12), 845 => to_unsigned(2137, 12), 846 => to_unsigned(1870, 12), 847 => to_unsigned(1902, 12), 848 => to_unsigned(2122, 12), 849 => to_unsigned(2197, 12), 850 => to_unsigned(2537, 12), 851 => to_unsigned(2196, 12), 852 => to_unsigned(1823, 12), 853 => to_unsigned(2197, 12), 854 => to_unsigned(1735, 12), 855 => to_unsigned(1967, 12), 856 => to_unsigned(1850, 12), 857 => to_unsigned(1968, 12), 858 => to_unsigned(2000, 12), 859 => to_unsigned(1551, 12), 860 => to_unsigned(1424, 12), 861 => to_unsigned(1855, 12), 862 => to_unsigned(1957, 12), 863 => to_unsigned(1126, 12), 864 => to_unsigned(1980, 12), 865 => to_unsigned(2056, 12), 866 => to_unsigned(2216, 12), 867 => to_unsigned(2534, 12), 868 => to_unsigned(1589, 12), 869 => to_unsigned(2423, 12), 870 => to_unsigned(1686, 12), 871 => to_unsigned(1775, 12), 872 => to_unsigned(1945, 12), 873 => to_unsigned(1973, 12), 874 => to_unsigned(1463, 12), 875 => to_unsigned(1888, 12), 876 => to_unsigned(1385, 12), 877 => to_unsigned(2069, 12), 878 => to_unsigned(1938, 12), 879 => to_unsigned(1985, 12), 880 => to_unsigned(2405, 12), 881 => to_unsigned(2098, 12), 882 => to_unsigned(1985, 12), 883 => to_unsigned(2441, 12), 884 => to_unsigned(1640, 12), 885 => to_unsigned(2406, 12), 886 => to_unsigned(2249, 12), 887 => to_unsigned(1759, 12), 888 => to_unsigned(2510, 12), 889 => to_unsigned(2549, 12), 890 => to_unsigned(2382, 12), 891 => to_unsigned(2619, 12), 892 => to_unsigned(2325, 12), 893 => to_unsigned(2964, 12), 894 => to_unsigned(1625, 12), 895 => to_unsigned(2280, 12), 896 => to_unsigned(2122, 12), 897 => to_unsigned(1855, 12), 898 => to_unsigned(1938, 12), 899 => to_unsigned(2565, 12), 900 => to_unsigned(2105, 12), 901 => to_unsigned(2293, 12), 902 => to_unsigned(1617, 12), 903 => to_unsigned(1689, 12), 904 => to_unsigned(2476, 12), 905 => to_unsigned(2013, 12), 906 => to_unsigned(1387, 12), 907 => to_unsigned(1809, 12), 908 => to_unsigned(1938, 12), 909 => to_unsigned(1948, 12), 910 => to_unsigned(1818, 12), 911 => to_unsigned(2411, 12), 912 => to_unsigned(2128, 12), 913 => to_unsigned(2114, 12), 914 => to_unsigned(3009, 12), 915 => to_unsigned(1912, 12), 916 => to_unsigned(2209, 12), 917 => to_unsigned(1551, 12), 918 => to_unsigned(1910, 12), 919 => to_unsigned(1583, 12), 920 => to_unsigned(1950, 12), 921 => to_unsigned(2148, 12), 922 => to_unsigned(2080, 12), 923 => to_unsigned(2198, 12), 924 => to_unsigned(1430, 12), 925 => to_unsigned(1929, 12), 926 => to_unsigned(2814, 12), 927 => to_unsigned(1976, 12), 928 => to_unsigned(2126, 12), 929 => to_unsigned(1721, 12), 930 => to_unsigned(2561, 12), 931 => to_unsigned(2161, 12), 932 => to_unsigned(1960, 12), 933 => to_unsigned(2580, 12), 934 => to_unsigned(1941, 12), 935 => to_unsigned(2231, 12), 936 => to_unsigned(1988, 12), 937 => to_unsigned(1799, 12), 938 => to_unsigned(2377, 12), 939 => to_unsigned(2363, 12), 940 => to_unsigned(2369, 12), 941 => to_unsigned(1904, 12), 942 => to_unsigned(2062, 12), 943 => to_unsigned(2153, 12), 944 => to_unsigned(2356, 12), 945 => to_unsigned(2557, 12), 946 => to_unsigned(2437, 12), 947 => to_unsigned(2055, 12), 948 => to_unsigned(2095, 12), 949 => to_unsigned(1599, 12), 950 => to_unsigned(968, 12), 951 => to_unsigned(2318, 12), 952 => to_unsigned(1580, 12), 953 => to_unsigned(2184, 12), 954 => to_unsigned(2172, 12), 955 => to_unsigned(1769, 12), 956 => to_unsigned(1705, 12), 957 => to_unsigned(1969, 12), 958 => to_unsigned(2916, 12), 959 => to_unsigned(1604, 12), 960 => to_unsigned(2532, 12), 961 => to_unsigned(2477, 12), 962 => to_unsigned(3107, 12), 963 => to_unsigned(2133, 12), 964 => to_unsigned(1660, 12), 965 => to_unsigned(1499, 12), 966 => to_unsigned(1508, 12), 967 => to_unsigned(2386, 12), 968 => to_unsigned(1961, 12), 969 => to_unsigned(1712, 12), 970 => to_unsigned(2810, 12), 971 => to_unsigned(2314, 12), 972 => to_unsigned(1927, 12), 973 => to_unsigned(1592, 12), 974 => to_unsigned(2256, 12), 975 => to_unsigned(1743, 12), 976 => to_unsigned(2373, 12), 977 => to_unsigned(1878, 12), 978 => to_unsigned(1641, 12), 979 => to_unsigned(2133, 12), 980 => to_unsigned(2301, 12), 981 => to_unsigned(1975, 12), 982 => to_unsigned(2330, 12), 983 => to_unsigned(1992, 12), 984 => to_unsigned(2029, 12), 985 => to_unsigned(2114, 12), 986 => to_unsigned(1643, 12), 987 => to_unsigned(1923, 12), 988 => to_unsigned(1537, 12), 989 => to_unsigned(2282, 12), 990 => to_unsigned(2170, 12), 991 => to_unsigned(1498, 12), 992 => to_unsigned(1786, 12), 993 => to_unsigned(1756, 12), 994 => to_unsigned(1905, 12), 995 => to_unsigned(1479, 12), 996 => to_unsigned(2214, 12), 997 => to_unsigned(2278, 12), 998 => to_unsigned(2510, 12), 999 => to_unsigned(2038, 12), 1000 => to_unsigned(2873, 12), 1001 => to_unsigned(1655, 12), 1002 => to_unsigned(1872, 12), 1003 => to_unsigned(1814, 12), 1004 => to_unsigned(2256, 12), 1005 => to_unsigned(2272, 12), 1006 => to_unsigned(1720, 12), 1007 => to_unsigned(2188, 12), 1008 => to_unsigned(2499, 12), 1009 => to_unsigned(1597, 12), 1010 => to_unsigned(2856, 12), 1011 => to_unsigned(2481, 12), 1012 => to_unsigned(2449, 12), 1013 => to_unsigned(1745, 12), 1014 => to_unsigned(1800, 12), 1015 => to_unsigned(1790, 12), 1016 => to_unsigned(2412, 12), 1017 => to_unsigned(2118, 12), 1018 => to_unsigned(1350, 12), 1019 => to_unsigned(1748, 12), 1020 => to_unsigned(1870, 12), 1021 => to_unsigned(1919, 12), 1022 => to_unsigned(1489, 12), 1023 => to_unsigned(1364, 12), 1024 => to_unsigned(1645, 12), 1025 => to_unsigned(1737, 12), 1026 => to_unsigned(1878, 12), 1027 => to_unsigned(1462, 12), 1028 => to_unsigned(2074, 12), 1029 => to_unsigned(1664, 12), 1030 => to_unsigned(2448, 12), 1031 => to_unsigned(2018, 12), 1032 => to_unsigned(1696, 12), 1033 => to_unsigned(2093, 12), 1034 => to_unsigned(1767, 12), 1035 => to_unsigned(1340, 12), 1036 => to_unsigned(2149, 12), 1037 => to_unsigned(1287, 12), 1038 => to_unsigned(2111, 12), 1039 => to_unsigned(1878, 12), 1040 => to_unsigned(2579, 12), 1041 => to_unsigned(2284, 12), 1042 => to_unsigned(1988, 12), 1043 => to_unsigned(1872, 12), 1044 => to_unsigned(2170, 12), 1045 => to_unsigned(1772, 12), 1046 => to_unsigned(2640, 12), 1047 => to_unsigned(1924, 12), 1048 => to_unsigned(1753, 12), 1049 => to_unsigned(2087, 12), 1050 => to_unsigned(1939, 12), 1051 => to_unsigned(2018, 12), 1052 => to_unsigned(1302, 12), 1053 => to_unsigned(1642, 12), 1054 => to_unsigned(1945, 12), 1055 => to_unsigned(1576, 12), 1056 => to_unsigned(2270, 12), 1057 => to_unsigned(1589, 12), 1058 => to_unsigned(1845, 12), 1059 => to_unsigned(2342, 12), 1060 => to_unsigned(2462, 12), 1061 => to_unsigned(1534, 12), 1062 => to_unsigned(2221, 12), 1063 => to_unsigned(2157, 12), 1064 => to_unsigned(1895, 12), 1065 => to_unsigned(2229, 12), 1066 => to_unsigned(1849, 12), 1067 => to_unsigned(2655, 12), 1068 => to_unsigned(2326, 12), 1069 => to_unsigned(2035, 12), 1070 => to_unsigned(2299, 12), 1071 => to_unsigned(1727, 12), 1072 => to_unsigned(1836, 12), 1073 => to_unsigned(1999, 12), 1074 => to_unsigned(1791, 12), 1075 => to_unsigned(2527, 12), 1076 => to_unsigned(1954, 12), 1077 => to_unsigned(1942, 12), 1078 => to_unsigned(2365, 12), 1079 => to_unsigned(1794, 12), 1080 => to_unsigned(2110, 12), 1081 => to_unsigned(2393, 12), 1082 => to_unsigned(2139, 12), 1083 => to_unsigned(2542, 12), 1084 => to_unsigned(1514, 12), 1085 => to_unsigned(2161, 12), 1086 => to_unsigned(2430, 12), 1087 => to_unsigned(2479, 12), 1088 => to_unsigned(2597, 12), 1089 => to_unsigned(2594, 12), 1090 => to_unsigned(2627, 12), 1091 => to_unsigned(1822, 12), 1092 => to_unsigned(2417, 12), 1093 => to_unsigned(1715, 12), 1094 => to_unsigned(1472, 12), 1095 => to_unsigned(1899, 12), 1096 => to_unsigned(1952, 12), 1097 => to_unsigned(2196, 12), 1098 => to_unsigned(2680, 12), 1099 => to_unsigned(1765, 12), 1100 => to_unsigned(1573, 12), 1101 => to_unsigned(2323, 12), 1102 => to_unsigned(2037, 12), 1103 => to_unsigned(2422, 12), 1104 => to_unsigned(1526, 12), 1105 => to_unsigned(1537, 12), 1106 => to_unsigned(1889, 12), 1107 => to_unsigned(2030, 12), 1108 => to_unsigned(1699, 12), 1109 => to_unsigned(1952, 12), 1110 => to_unsigned(2001, 12), 1111 => to_unsigned(2583, 12), 1112 => to_unsigned(2777, 12), 1113 => to_unsigned(1893, 12), 1114 => to_unsigned(1432, 12), 1115 => to_unsigned(2447, 12), 1116 => to_unsigned(2185, 12), 1117 => to_unsigned(2240, 12), 1118 => to_unsigned(2236, 12), 1119 => to_unsigned(2082, 12), 1120 => to_unsigned(2265, 12), 1121 => to_unsigned(2407, 12), 1122 => to_unsigned(1912, 12), 1123 => to_unsigned(1835, 12), 1124 => to_unsigned(2557, 12), 1125 => to_unsigned(2071, 12), 1126 => to_unsigned(2085, 12), 1127 => to_unsigned(2559, 12), 1128 => to_unsigned(2572, 12), 1129 => to_unsigned(2505, 12), 1130 => to_unsigned(2224, 12), 1131 => to_unsigned(2259, 12), 1132 => to_unsigned(1819, 12), 1133 => to_unsigned(2517, 12), 1134 => to_unsigned(2651, 12), 1135 => to_unsigned(2276, 12), 1136 => to_unsigned(2107, 12), 1137 => to_unsigned(2473, 12), 1138 => to_unsigned(2254, 12), 1139 => to_unsigned(1746, 12), 1140 => to_unsigned(2142, 12), 1141 => to_unsigned(2242, 12), 1142 => to_unsigned(2127, 12), 1143 => to_unsigned(2531, 12), 1144 => to_unsigned(1633, 12), 1145 => to_unsigned(1997, 12), 1146 => to_unsigned(2245, 12), 1147 => to_unsigned(2112, 12), 1148 => to_unsigned(1913, 12), 1149 => to_unsigned(2695, 12), 1150 => to_unsigned(1639, 12), 1151 => to_unsigned(2027, 12), 1152 => to_unsigned(1850, 12), 1153 => to_unsigned(2673, 12), 1154 => to_unsigned(2287, 12), 1155 => to_unsigned(2402, 12), 1156 => to_unsigned(2153, 12), 1157 => to_unsigned(2483, 12), 1158 => to_unsigned(2024, 12), 1159 => to_unsigned(2175, 12), 1160 => to_unsigned(1664, 12), 1161 => to_unsigned(1496, 12), 1162 => to_unsigned(1622, 12), 1163 => to_unsigned(1896, 12), 1164 => to_unsigned(2125, 12), 1165 => to_unsigned(2420, 12), 1166 => to_unsigned(2588, 12), 1167 => to_unsigned(1685, 12), 1168 => to_unsigned(2020, 12), 1169 => to_unsigned(2007, 12), 1170 => to_unsigned(1811, 12), 1171 => to_unsigned(1595, 12), 1172 => to_unsigned(2688, 12), 1173 => to_unsigned(2798, 12), 1174 => to_unsigned(1940, 12), 1175 => to_unsigned(1783, 12), 1176 => to_unsigned(2114, 12), 1177 => to_unsigned(2473, 12), 1178 => to_unsigned(2829, 12), 1179 => to_unsigned(1626, 12), 1180 => to_unsigned(2001, 12), 1181 => to_unsigned(1515, 12), 1182 => to_unsigned(1919, 12), 1183 => to_unsigned(1627, 12), 1184 => to_unsigned(1946, 12), 1185 => to_unsigned(1903, 12), 1186 => to_unsigned(2146, 12), 1187 => to_unsigned(1905, 12), 1188 => to_unsigned(1740, 12), 1189 => to_unsigned(2071, 12), 1190 => to_unsigned(2236, 12), 1191 => to_unsigned(2173, 12), 1192 => to_unsigned(2474, 12), 1193 => to_unsigned(1774, 12), 1194 => to_unsigned(1789, 12), 1195 => to_unsigned(2507, 12), 1196 => to_unsigned(2030, 12), 1197 => to_unsigned(2553, 12), 1198 => to_unsigned(2504, 12), 1199 => to_unsigned(2394, 12), 1200 => to_unsigned(1690, 12), 1201 => to_unsigned(2171, 12), 1202 => to_unsigned(2739, 12), 1203 => to_unsigned(1715, 12), 1204 => to_unsigned(1728, 12), 1205 => to_unsigned(2349, 12), 1206 => to_unsigned(2163, 12), 1207 => to_unsigned(2184, 12), 1208 => to_unsigned(1903, 12), 1209 => to_unsigned(1514, 12), 1210 => to_unsigned(2205, 12), 1211 => to_unsigned(1933, 12), 1212 => to_unsigned(2675, 12), 1213 => to_unsigned(2510, 12), 1214 => to_unsigned(1989, 12), 1215 => to_unsigned(1975, 12), 1216 => to_unsigned(1653, 12), 1217 => to_unsigned(2411, 12), 1218 => to_unsigned(2357, 12), 1219 => to_unsigned(1495, 12), 1220 => to_unsigned(2086, 12), 1221 => to_unsigned(2286, 12), 1222 => to_unsigned(1767, 12), 1223 => to_unsigned(1720, 12), 1224 => to_unsigned(1898, 12), 1225 => to_unsigned(1492, 12), 1226 => to_unsigned(2371, 12), 1227 => to_unsigned(2205, 12), 1228 => to_unsigned(2022, 12), 1229 => to_unsigned(1785, 12), 1230 => to_unsigned(2858, 12), 1231 => to_unsigned(2525, 12), 1232 => to_unsigned(1850, 12), 1233 => to_unsigned(2355, 12), 1234 => to_unsigned(2075, 12), 1235 => to_unsigned(1689, 12), 1236 => to_unsigned(1782, 12), 1237 => to_unsigned(2074, 12), 1238 => to_unsigned(2436, 12), 1239 => to_unsigned(2638, 12), 1240 => to_unsigned(2390, 12), 1241 => to_unsigned(2126, 12), 1242 => to_unsigned(1884, 12), 1243 => to_unsigned(1706, 12), 1244 => to_unsigned(1431, 12), 1245 => to_unsigned(2437, 12), 1246 => to_unsigned(2036, 12), 1247 => to_unsigned(2256, 12), 1248 => to_unsigned(1709, 12), 1249 => to_unsigned(2070, 12), 1250 => to_unsigned(2150, 12), 1251 => to_unsigned(1134, 12), 1252 => to_unsigned(859, 12), 1253 => to_unsigned(1611, 12), 1254 => to_unsigned(2215, 12), 1255 => to_unsigned(2230, 12), 1256 => to_unsigned(1578, 12), 1257 => to_unsigned(1800, 12), 1258 => to_unsigned(1930, 12), 1259 => to_unsigned(1854, 12), 1260 => to_unsigned(1758, 12), 1261 => to_unsigned(1804, 12), 1262 => to_unsigned(2482, 12), 1263 => to_unsigned(1612, 12), 1264 => to_unsigned(1880, 12), 1265 => to_unsigned(2507, 12), 1266 => to_unsigned(1572, 12), 1267 => to_unsigned(1747, 12), 1268 => to_unsigned(1270, 12), 1269 => to_unsigned(2264, 12), 1270 => to_unsigned(2388, 12), 1271 => to_unsigned(2443, 12), 1272 => to_unsigned(2705, 12), 1273 => to_unsigned(1805, 12), 1274 => to_unsigned(1556, 12), 1275 => to_unsigned(2139, 12), 1276 => to_unsigned(2606, 12), 1277 => to_unsigned(2511, 12), 1278 => to_unsigned(2351, 12), 1279 => to_unsigned(1514, 12), 1280 => to_unsigned(2088, 12), 1281 => to_unsigned(2686, 12), 1282 => to_unsigned(2200, 12), 1283 => to_unsigned(2262, 12), 1284 => to_unsigned(2474, 12), 1285 => to_unsigned(2052, 12), 1286 => to_unsigned(2318, 12), 1287 => to_unsigned(2244, 12), 1288 => to_unsigned(1775, 12), 1289 => to_unsigned(2442, 12), 1290 => to_unsigned(1915, 12), 1291 => to_unsigned(1999, 12), 1292 => to_unsigned(1473, 12), 1293 => to_unsigned(1244, 12), 1294 => to_unsigned(1892, 12), 1295 => to_unsigned(1577, 12), 1296 => to_unsigned(1795, 12), 1297 => to_unsigned(2794, 12), 1298 => to_unsigned(2100, 12), 1299 => to_unsigned(1501, 12), 1300 => to_unsigned(1731, 12), 1301 => to_unsigned(1691, 12), 1302 => to_unsigned(1777, 12), 1303 => to_unsigned(2488, 12), 1304 => to_unsigned(2123, 12), 1305 => to_unsigned(1332, 12), 1306 => to_unsigned(2118, 12), 1307 => to_unsigned(2418, 12), 1308 => to_unsigned(2385, 12), 1309 => to_unsigned(2113, 12), 1310 => to_unsigned(1962, 12), 1311 => to_unsigned(2217, 12), 1312 => to_unsigned(1841, 12), 1313 => to_unsigned(2147, 12), 1314 => to_unsigned(2249, 12), 1315 => to_unsigned(1892, 12), 1316 => to_unsigned(2420, 12), 1317 => to_unsigned(1406, 12), 1318 => to_unsigned(1759, 12), 1319 => to_unsigned(2260, 12), 1320 => to_unsigned(2299, 12), 1321 => to_unsigned(2531, 12), 1322 => to_unsigned(1669, 12), 1323 => to_unsigned(1495, 12), 1324 => to_unsigned(2560, 12), 1325 => to_unsigned(2435, 12), 1326 => to_unsigned(2374, 12), 1327 => to_unsigned(2611, 12), 1328 => to_unsigned(2317, 12), 1329 => to_unsigned(1785, 12), 1330 => to_unsigned(2509, 12), 1331 => to_unsigned(2017, 12), 1332 => to_unsigned(2420, 12), 1333 => to_unsigned(1717, 12), 1334 => to_unsigned(2361, 12), 1335 => to_unsigned(2118, 12), 1336 => to_unsigned(2164, 12), 1337 => to_unsigned(1697, 12), 1338 => to_unsigned(1932, 12), 1339 => to_unsigned(2038, 12), 1340 => to_unsigned(1829, 12), 1341 => to_unsigned(1370, 12), 1342 => to_unsigned(1729, 12), 1343 => to_unsigned(1624, 12), 1344 => to_unsigned(1344, 12), 1345 => to_unsigned(2040, 12), 1346 => to_unsigned(1835, 12), 1347 => to_unsigned(2376, 12), 1348 => to_unsigned(1576, 12), 1349 => to_unsigned(2245, 12), 1350 => to_unsigned(1822, 12), 1351 => to_unsigned(1705, 12), 1352 => to_unsigned(2065, 12), 1353 => to_unsigned(1938, 12), 1354 => to_unsigned(1777, 12), 1355 => to_unsigned(1889, 12), 1356 => to_unsigned(2362, 12), 1357 => to_unsigned(2154, 12), 1358 => to_unsigned(1427, 12), 1359 => to_unsigned(2081, 12), 1360 => to_unsigned(2593, 12), 1361 => to_unsigned(1646, 12), 1362 => to_unsigned(1911, 12), 1363 => to_unsigned(2330, 12), 1364 => to_unsigned(2455, 12), 1365 => to_unsigned(1257, 12), 1366 => to_unsigned(1530, 12), 1367 => to_unsigned(1915, 12), 1368 => to_unsigned(1853, 12), 1369 => to_unsigned(2438, 12), 1370 => to_unsigned(1786, 12), 1371 => to_unsigned(2594, 12), 1372 => to_unsigned(2128, 12), 1373 => to_unsigned(1996, 12), 1374 => to_unsigned(1820, 12), 1375 => to_unsigned(2469, 12), 1376 => to_unsigned(1647, 12), 1377 => to_unsigned(2379, 12), 1378 => to_unsigned(1975, 12), 1379 => to_unsigned(2372, 12), 1380 => to_unsigned(2218, 12), 1381 => to_unsigned(2246, 12), 1382 => to_unsigned(2510, 12), 1383 => to_unsigned(2617, 12), 1384 => to_unsigned(2405, 12), 1385 => to_unsigned(1824, 12), 1386 => to_unsigned(1905, 12), 1387 => to_unsigned(1673, 12), 1388 => to_unsigned(2069, 12), 1389 => to_unsigned(1896, 12), 1390 => to_unsigned(2151, 12), 1391 => to_unsigned(2609, 12), 1392 => to_unsigned(2158, 12), 1393 => to_unsigned(1946, 12), 1394 => to_unsigned(2151, 12), 1395 => to_unsigned(1905, 12), 1396 => to_unsigned(2042, 12), 1397 => to_unsigned(2135, 12), 1398 => to_unsigned(2351, 12), 1399 => to_unsigned(1959, 12), 1400 => to_unsigned(1826, 12), 1401 => to_unsigned(2161, 12), 1402 => to_unsigned(1517, 12), 1403 => to_unsigned(2368, 12), 1404 => to_unsigned(1884, 12), 1405 => to_unsigned(1763, 12), 1406 => to_unsigned(1995, 12), 1407 => to_unsigned(2636, 12), 1408 => to_unsigned(1661, 12), 1409 => to_unsigned(2784, 12), 1410 => to_unsigned(2028, 12), 1411 => to_unsigned(2061, 12), 1412 => to_unsigned(2047, 12), 1413 => to_unsigned(1860, 12), 1414 => to_unsigned(1603, 12), 1415 => to_unsigned(1216, 12), 1416 => to_unsigned(2385, 12), 1417 => to_unsigned(1285, 12), 1418 => to_unsigned(2262, 12), 1419 => to_unsigned(1186, 12), 1420 => to_unsigned(2958, 12), 1421 => to_unsigned(2185, 12), 1422 => to_unsigned(2460, 12), 1423 => to_unsigned(2232, 12), 1424 => to_unsigned(2131, 12), 1425 => to_unsigned(1793, 12), 1426 => to_unsigned(2283, 12), 1427 => to_unsigned(1839, 12), 1428 => to_unsigned(1408, 12), 1429 => to_unsigned(2100, 12), 1430 => to_unsigned(1958, 12), 1431 => to_unsigned(1972, 12), 1432 => to_unsigned(2042, 12), 1433 => to_unsigned(2431, 12), 1434 => to_unsigned(2278, 12), 1435 => to_unsigned(2489, 12), 1436 => to_unsigned(2322, 12), 1437 => to_unsigned(2091, 12), 1438 => to_unsigned(2043, 12), 1439 => to_unsigned(1874, 12), 1440 => to_unsigned(2886, 12), 1441 => to_unsigned(1675, 12), 1442 => to_unsigned(2162, 12), 1443 => to_unsigned(1919, 12), 1444 => to_unsigned(2569, 12), 1445 => to_unsigned(2166, 12), 1446 => to_unsigned(1623, 12), 1447 => to_unsigned(2064, 12), 1448 => to_unsigned(1495, 12), 1449 => to_unsigned(1920, 12), 1450 => to_unsigned(1765, 12), 1451 => to_unsigned(1817, 12), 1452 => to_unsigned(2083, 12), 1453 => to_unsigned(1529, 12), 1454 => to_unsigned(1818, 12), 1455 => to_unsigned(2300, 12), 1456 => to_unsigned(1192, 12), 1457 => to_unsigned(2406, 12), 1458 => to_unsigned(2203, 12), 1459 => to_unsigned(1796, 12), 1460 => to_unsigned(2221, 12), 1461 => to_unsigned(1539, 12), 1462 => to_unsigned(2337, 12), 1463 => to_unsigned(2108, 12), 1464 => to_unsigned(1752, 12), 1465 => to_unsigned(2220, 12), 1466 => to_unsigned(2202, 12), 1467 => to_unsigned(1679, 12), 1468 => to_unsigned(1755, 12), 1469 => to_unsigned(1489, 12), 1470 => to_unsigned(1927, 12), 1471 => to_unsigned(1924, 12), 1472 => to_unsigned(2225, 12), 1473 => to_unsigned(2155, 12), 1474 => to_unsigned(1655, 12), 1475 => to_unsigned(2848, 12), 1476 => to_unsigned(2318, 12), 1477 => to_unsigned(1466, 12), 1478 => to_unsigned(2296, 12), 1479 => to_unsigned(2124, 12), 1480 => to_unsigned(2126, 12), 1481 => to_unsigned(1862, 12), 1482 => to_unsigned(1406, 12), 1483 => to_unsigned(1582, 12), 1484 => to_unsigned(2368, 12), 1485 => to_unsigned(2197, 12), 1486 => to_unsigned(1662, 12), 1487 => to_unsigned(2939, 12), 1488 => to_unsigned(2117, 12), 1489 => to_unsigned(2270, 12), 1490 => to_unsigned(1905, 12), 1491 => to_unsigned(2034, 12), 1492 => to_unsigned(1990, 12), 1493 => to_unsigned(1019, 12), 1494 => to_unsigned(2225, 12), 1495 => to_unsigned(1734, 12), 1496 => to_unsigned(1824, 12), 1497 => to_unsigned(2412, 12), 1498 => to_unsigned(1882, 12), 1499 => to_unsigned(2236, 12), 1500 => to_unsigned(1995, 12), 1501 => to_unsigned(2522, 12), 1502 => to_unsigned(2819, 12), 1503 => to_unsigned(2683, 12), 1504 => to_unsigned(2155, 12), 1505 => to_unsigned(2175, 12), 1506 => to_unsigned(2204, 12), 1507 => to_unsigned(2417, 12), 1508 => to_unsigned(2338, 12), 1509 => to_unsigned(2251, 12), 1510 => to_unsigned(2021, 12), 1511 => to_unsigned(1604, 12), 1512 => to_unsigned(2138, 12), 1513 => to_unsigned(1636, 12), 1514 => to_unsigned(2460, 12), 1515 => to_unsigned(1972, 12), 1516 => to_unsigned(2021, 12), 1517 => to_unsigned(2575, 12), 1518 => to_unsigned(2219, 12), 1519 => to_unsigned(2375, 12), 1520 => to_unsigned(1783, 12), 1521 => to_unsigned(1941, 12), 1522 => to_unsigned(2006, 12), 1523 => to_unsigned(1723, 12), 1524 => to_unsigned(1939, 12), 1525 => to_unsigned(2095, 12), 1526 => to_unsigned(1572, 12), 1527 => to_unsigned(1896, 12), 1528 => to_unsigned(2254, 12), 1529 => to_unsigned(2208, 12), 1530 => to_unsigned(2628, 12), 1531 => to_unsigned(2192, 12), 1532 => to_unsigned(1501, 12), 1533 => to_unsigned(2150, 12), 1534 => to_unsigned(1810, 12), 1535 => to_unsigned(2506, 12), 1536 => to_unsigned(2567, 12), 1537 => to_unsigned(2068, 12), 1538 => to_unsigned(1482, 12), 1539 => to_unsigned(2363, 12), 1540 => to_unsigned(2549, 12), 1541 => to_unsigned(1266, 12), 1542 => to_unsigned(3027, 12), 1543 => to_unsigned(2659, 12), 1544 => to_unsigned(1845, 12), 1545 => to_unsigned(1787, 12), 1546 => to_unsigned(2007, 12), 1547 => to_unsigned(2063, 12), 1548 => to_unsigned(2312, 12), 1549 => to_unsigned(1600, 12), 1550 => to_unsigned(1843, 12), 1551 => to_unsigned(1352, 12), 1552 => to_unsigned(2661, 12), 1553 => to_unsigned(2001, 12), 1554 => to_unsigned(2072, 12), 1555 => to_unsigned(2068, 12), 1556 => to_unsigned(2067, 12), 1557 => to_unsigned(2369, 12), 1558 => to_unsigned(2396, 12), 1559 => to_unsigned(1933, 12), 1560 => to_unsigned(1729, 12), 1561 => to_unsigned(2147, 12), 1562 => to_unsigned(1853, 12), 1563 => to_unsigned(2193, 12), 1564 => to_unsigned(1202, 12), 1565 => to_unsigned(2283, 12), 1566 => to_unsigned(2010, 12), 1567 => to_unsigned(1783, 12), 1568 => to_unsigned(1993, 12), 1569 => to_unsigned(2292, 12), 1570 => to_unsigned(1308, 12), 1571 => to_unsigned(2414, 12), 1572 => to_unsigned(2383, 12), 1573 => to_unsigned(1333, 12), 1574 => to_unsigned(1905, 12), 1575 => to_unsigned(2307, 12), 1576 => to_unsigned(2406, 12), 1577 => to_unsigned(2058, 12), 1578 => to_unsigned(2233, 12), 1579 => to_unsigned(2069, 12), 1580 => to_unsigned(1716, 12), 1581 => to_unsigned(2313, 12), 1582 => to_unsigned(2266, 12), 1583 => to_unsigned(2376, 12), 1584 => to_unsigned(2593, 12), 1585 => to_unsigned(1402, 12), 1586 => to_unsigned(1460, 12), 1587 => to_unsigned(1793, 12), 1588 => to_unsigned(1523, 12), 1589 => to_unsigned(2042, 12), 1590 => to_unsigned(1844, 12), 1591 => to_unsigned(2520, 12), 1592 => to_unsigned(1626, 12), 1593 => to_unsigned(2102, 12), 1594 => to_unsigned(2301, 12), 1595 => to_unsigned(2241, 12), 1596 => to_unsigned(1390, 12), 1597 => to_unsigned(1868, 12), 1598 => to_unsigned(1601, 12), 1599 => to_unsigned(1552, 12), 1600 => to_unsigned(1908, 12), 1601 => to_unsigned(1747, 12), 1602 => to_unsigned(2394, 12), 1603 => to_unsigned(2445, 12), 1604 => to_unsigned(1499, 12), 1605 => to_unsigned(2366, 12), 1606 => to_unsigned(2047, 12), 1607 => to_unsigned(2258, 12), 1608 => to_unsigned(1921, 12), 1609 => to_unsigned(1869, 12), 1610 => to_unsigned(2012, 12), 1611 => to_unsigned(1883, 12), 1612 => to_unsigned(2009, 12), 1613 => to_unsigned(2338, 12), 1614 => to_unsigned(1835, 12), 1615 => to_unsigned(1967, 12), 1616 => to_unsigned(2106, 12), 1617 => to_unsigned(1841, 12), 1618 => to_unsigned(1911, 12), 1619 => to_unsigned(1706, 12), 1620 => to_unsigned(1757, 12), 1621 => to_unsigned(2102, 12), 1622 => to_unsigned(1513, 12), 1623 => to_unsigned(1923, 12), 1624 => to_unsigned(1354, 12), 1625 => to_unsigned(2507, 12), 1626 => to_unsigned(2379, 12), 1627 => to_unsigned(2245, 12), 1628 => to_unsigned(2235, 12), 1629 => to_unsigned(2195, 12), 1630 => to_unsigned(2244, 12), 1631 => to_unsigned(2008, 12), 1632 => to_unsigned(2065, 12), 1633 => to_unsigned(1517, 12), 1634 => to_unsigned(2304, 12), 1635 => to_unsigned(1515, 12), 1636 => to_unsigned(1583, 12), 1637 => to_unsigned(1939, 12), 1638 => to_unsigned(1900, 12), 1639 => to_unsigned(2720, 12), 1640 => to_unsigned(1960, 12), 1641 => to_unsigned(2735, 12), 1642 => to_unsigned(1748, 12), 1643 => to_unsigned(1667, 12), 1644 => to_unsigned(2090, 12), 1645 => to_unsigned(1908, 12), 1646 => to_unsigned(2359, 12), 1647 => to_unsigned(1945, 12), 1648 => to_unsigned(2271, 12), 1649 => to_unsigned(2309, 12), 1650 => to_unsigned(2194, 12), 1651 => to_unsigned(2663, 12), 1652 => to_unsigned(2641, 12), 1653 => to_unsigned(2332, 12), 1654 => to_unsigned(1830, 12), 1655 => to_unsigned(2521, 12), 1656 => to_unsigned(2570, 12), 1657 => to_unsigned(2663, 12), 1658 => to_unsigned(1746, 12), 1659 => to_unsigned(1867, 12), 1660 => to_unsigned(2178, 12), 1661 => to_unsigned(2178, 12), 1662 => to_unsigned(1858, 12), 1663 => to_unsigned(2413, 12), 1664 => to_unsigned(2058, 12), 1665 => to_unsigned(1288, 12), 1666 => to_unsigned(2469, 12), 1667 => to_unsigned(2219, 12), 1668 => to_unsigned(2483, 12), 1669 => to_unsigned(1988, 12), 1670 => to_unsigned(2452, 12), 1671 => to_unsigned(2216, 12), 1672 => to_unsigned(1621, 12), 1673 => to_unsigned(1500, 12), 1674 => to_unsigned(1955, 12), 1675 => to_unsigned(2307, 12), 1676 => to_unsigned(2315, 12), 1677 => to_unsigned(1467, 12), 1678 => to_unsigned(2000, 12), 1679 => to_unsigned(1839, 12), 1680 => to_unsigned(2570, 12), 1681 => to_unsigned(1674, 12), 1682 => to_unsigned(1579, 12), 1683 => to_unsigned(2235, 12), 1684 => to_unsigned(1759, 12), 1685 => to_unsigned(2403, 12), 1686 => to_unsigned(2810, 12), 1687 => to_unsigned(2071, 12), 1688 => to_unsigned(1990, 12), 1689 => to_unsigned(1692, 12), 1690 => to_unsigned(1935, 12), 1691 => to_unsigned(2625, 12), 1692 => to_unsigned(1831, 12), 1693 => to_unsigned(2761, 12), 1694 => to_unsigned(2156, 12), 1695 => to_unsigned(2227, 12), 1696 => to_unsigned(1846, 12), 1697 => to_unsigned(1767, 12), 1698 => to_unsigned(1346, 12), 1699 => to_unsigned(2035, 12), 1700 => to_unsigned(1775, 12), 1701 => to_unsigned(2026, 12), 1702 => to_unsigned(2568, 12), 1703 => to_unsigned(2435, 12), 1704 => to_unsigned(1876, 12), 1705 => to_unsigned(2146, 12), 1706 => to_unsigned(2171, 12), 1707 => to_unsigned(2244, 12), 1708 => to_unsigned(1935, 12), 1709 => to_unsigned(2414, 12), 1710 => to_unsigned(1969, 12), 1711 => to_unsigned(2389, 12), 1712 => to_unsigned(2587, 12), 1713 => to_unsigned(2238, 12), 1714 => to_unsigned(2097, 12), 1715 => to_unsigned(1728, 12), 1716 => to_unsigned(1642, 12), 1717 => to_unsigned(2020, 12), 1718 => to_unsigned(2158, 12), 1719 => to_unsigned(1860, 12), 1720 => to_unsigned(1781, 12), 1721 => to_unsigned(2073, 12), 1722 => to_unsigned(2295, 12), 1723 => to_unsigned(1869, 12), 1724 => to_unsigned(2014, 12), 1725 => to_unsigned(1336, 12), 1726 => to_unsigned(1980, 12), 1727 => to_unsigned(2157, 12), 1728 => to_unsigned(1987, 12), 1729 => to_unsigned(1647, 12), 1730 => to_unsigned(1756, 12), 1731 => to_unsigned(2807, 12), 1732 => to_unsigned(2549, 12), 1733 => to_unsigned(2389, 12), 1734 => to_unsigned(1306, 12), 1735 => to_unsigned(1808, 12), 1736 => to_unsigned(2639, 12), 1737 => to_unsigned(1939, 12), 1738 => to_unsigned(1434, 12), 1739 => to_unsigned(2227, 12), 1740 => to_unsigned(2076, 12), 1741 => to_unsigned(2146, 12), 1742 => to_unsigned(1581, 12), 1743 => to_unsigned(2378, 12), 1744 => to_unsigned(1972, 12), 1745 => to_unsigned(1628, 12), 1746 => to_unsigned(1689, 12), 1747 => to_unsigned(1823, 12), 1748 => to_unsigned(2039, 12), 1749 => to_unsigned(1884, 12), 1750 => to_unsigned(1853, 12), 1751 => to_unsigned(2589, 12), 1752 => to_unsigned(1660, 12), 1753 => to_unsigned(1909, 12), 1754 => to_unsigned(2362, 12), 1755 => to_unsigned(2110, 12), 1756 => to_unsigned(2024, 12), 1757 => to_unsigned(2556, 12), 1758 => to_unsigned(2097, 12), 1759 => to_unsigned(2533, 12), 1760 => to_unsigned(2289, 12), 1761 => to_unsigned(1764, 12), 1762 => to_unsigned(1895, 12), 1763 => to_unsigned(1895, 12), 1764 => to_unsigned(2268, 12), 1765 => to_unsigned(2545, 12), 1766 => to_unsigned(2290, 12), 1767 => to_unsigned(2656, 12), 1768 => to_unsigned(2917, 12), 1769 => to_unsigned(1876, 12), 1770 => to_unsigned(1534, 12), 1771 => to_unsigned(1919, 12), 1772 => to_unsigned(1955, 12), 1773 => to_unsigned(1506, 12), 1774 => to_unsigned(1939, 12), 1775 => to_unsigned(2170, 12), 1776 => to_unsigned(2761, 12), 1777 => to_unsigned(2210, 12), 1778 => to_unsigned(1741, 12), 1779 => to_unsigned(2517, 12), 1780 => to_unsigned(1661, 12), 1781 => to_unsigned(1590, 12), 1782 => to_unsigned(2269, 12), 1783 => to_unsigned(1726, 12), 1784 => to_unsigned(2332, 12), 1785 => to_unsigned(1781, 12), 1786 => to_unsigned(2140, 12), 1787 => to_unsigned(2335, 12), 1788 => to_unsigned(2194, 12), 1789 => to_unsigned(1582, 12), 1790 => to_unsigned(2077, 12), 1791 => to_unsigned(1903, 12), 1792 => to_unsigned(1889, 12), 1793 => to_unsigned(2272, 12), 1794 => to_unsigned(1767, 12), 1795 => to_unsigned(2457, 12), 1796 => to_unsigned(2331, 12), 1797 => to_unsigned(1573, 12), 1798 => to_unsigned(1991, 12), 1799 => to_unsigned(1879, 12), 1800 => to_unsigned(1392, 12), 1801 => to_unsigned(2195, 12), 1802 => to_unsigned(2346, 12), 1803 => to_unsigned(2178, 12), 1804 => to_unsigned(1826, 12), 1805 => to_unsigned(2041, 12), 1806 => to_unsigned(2379, 12), 1807 => to_unsigned(2101, 12), 1808 => to_unsigned(2346, 12), 1809 => to_unsigned(1919, 12), 1810 => to_unsigned(1495, 12), 1811 => to_unsigned(2146, 12), 1812 => to_unsigned(1889, 12), 1813 => to_unsigned(2160, 12), 1814 => to_unsigned(2149, 12), 1815 => to_unsigned(1610, 12), 1816 => to_unsigned(2112, 12), 1817 => to_unsigned(2005, 12), 1818 => to_unsigned(2244, 12), 1819 => to_unsigned(2362, 12), 1820 => to_unsigned(1613, 12), 1821 => to_unsigned(1307, 12), 1822 => to_unsigned(1811, 12), 1823 => to_unsigned(2340, 12), 1824 => to_unsigned(1887, 12), 1825 => to_unsigned(1763, 12), 1826 => to_unsigned(2518, 12), 1827 => to_unsigned(1841, 12), 1828 => to_unsigned(1768, 12), 1829 => to_unsigned(1879, 12), 1830 => to_unsigned(2456, 12), 1831 => to_unsigned(2688, 12), 1832 => to_unsigned(2576, 12), 1833 => to_unsigned(2750, 12), 1834 => to_unsigned(1564, 12), 1835 => to_unsigned(2392, 12), 1836 => to_unsigned(2209, 12), 1837 => to_unsigned(1778, 12), 1838 => to_unsigned(2126, 12), 1839 => to_unsigned(1412, 12), 1840 => to_unsigned(2108, 12), 1841 => to_unsigned(2330, 12), 1842 => to_unsigned(2167, 12), 1843 => to_unsigned(1420, 12), 1844 => to_unsigned(1532, 12), 1845 => to_unsigned(2122, 12), 1846 => to_unsigned(2025, 12), 1847 => to_unsigned(1986, 12), 1848 => to_unsigned(2555, 12), 1849 => to_unsigned(2452, 12), 1850 => to_unsigned(2285, 12), 1851 => to_unsigned(2291, 12), 1852 => to_unsigned(2527, 12), 1853 => to_unsigned(2203, 12), 1854 => to_unsigned(2033, 12), 1855 => to_unsigned(1406, 12), 1856 => to_unsigned(2351, 12), 1857 => to_unsigned(2387, 12), 1858 => to_unsigned(1767, 12), 1859 => to_unsigned(1755, 12), 1860 => to_unsigned(2391, 12), 1861 => to_unsigned(1755, 12), 1862 => to_unsigned(2204, 12), 1863 => to_unsigned(1716, 12), 1864 => to_unsigned(2016, 12), 1865 => to_unsigned(1710, 12), 1866 => to_unsigned(2006, 12), 1867 => to_unsigned(2240, 12), 1868 => to_unsigned(2669, 12), 1869 => to_unsigned(2101, 12), 1870 => to_unsigned(2090, 12), 1871 => to_unsigned(1601, 12), 1872 => to_unsigned(1139, 12), 1873 => to_unsigned(2040, 12), 1874 => to_unsigned(1359, 12), 1875 => to_unsigned(1781, 12), 1876 => to_unsigned(2262, 12), 1877 => to_unsigned(2154, 12), 1878 => to_unsigned(2034, 12), 1879 => to_unsigned(2253, 12), 1880 => to_unsigned(2341, 12), 1881 => to_unsigned(1503, 12), 1882 => to_unsigned(1830, 12), 1883 => to_unsigned(1597, 12), 1884 => to_unsigned(1441, 12), 1885 => to_unsigned(1689, 12), 1886 => to_unsigned(1711, 12), 1887 => to_unsigned(1559, 12), 1888 => to_unsigned(2224, 12), 1889 => to_unsigned(2222, 12), 1890 => to_unsigned(2185, 12), 1891 => to_unsigned(2157, 12), 1892 => to_unsigned(1683, 12), 1893 => to_unsigned(1141, 12), 1894 => to_unsigned(2514, 12), 1895 => to_unsigned(1853, 12), 1896 => to_unsigned(1991, 12), 1897 => to_unsigned(1950, 12), 1898 => to_unsigned(1781, 12), 1899 => to_unsigned(1649, 12), 1900 => to_unsigned(2117, 12), 1901 => to_unsigned(2078, 12), 1902 => to_unsigned(1819, 12), 1903 => to_unsigned(3055, 12), 1904 => to_unsigned(2348, 12), 1905 => to_unsigned(2055, 12), 1906 => to_unsigned(2351, 12), 1907 => to_unsigned(1968, 12), 1908 => to_unsigned(2174, 12), 1909 => to_unsigned(2288, 12), 1910 => to_unsigned(2009, 12), 1911 => to_unsigned(2230, 12), 1912 => to_unsigned(1580, 12), 1913 => to_unsigned(1772, 12), 1914 => to_unsigned(1810, 12), 1915 => to_unsigned(2110, 12), 1916 => to_unsigned(1683, 12), 1917 => to_unsigned(2311, 12), 1918 => to_unsigned(1868, 12), 1919 => to_unsigned(2132, 12), 1920 => to_unsigned(2221, 12), 1921 => to_unsigned(1576, 12), 1922 => to_unsigned(1902, 12), 1923 => to_unsigned(2109, 12), 1924 => to_unsigned(2391, 12), 1925 => to_unsigned(1576, 12), 1926 => to_unsigned(1796, 12), 1927 => to_unsigned(1860, 12), 1928 => to_unsigned(2198, 12), 1929 => to_unsigned(2124, 12), 1930 => to_unsigned(2125, 12), 1931 => to_unsigned(2064, 12), 1932 => to_unsigned(1957, 12), 1933 => to_unsigned(1846, 12), 1934 => to_unsigned(1803, 12), 1935 => to_unsigned(1555, 12), 1936 => to_unsigned(2270, 12), 1937 => to_unsigned(1985, 12), 1938 => to_unsigned(1696, 12), 1939 => to_unsigned(1726, 12), 1940 => to_unsigned(2287, 12), 1941 => to_unsigned(2815, 12), 1942 => to_unsigned(2432, 12), 1943 => to_unsigned(1748, 12), 1944 => to_unsigned(1878, 12), 1945 => to_unsigned(1266, 12), 1946 => to_unsigned(2061, 12), 1947 => to_unsigned(1758, 12), 1948 => to_unsigned(2323, 12), 1949 => to_unsigned(2467, 12), 1950 => to_unsigned(2017, 12), 1951 => to_unsigned(2878, 12), 1952 => to_unsigned(1780, 12), 1953 => to_unsigned(1979, 12), 1954 => to_unsigned(1981, 12), 1955 => to_unsigned(1712, 12), 1956 => to_unsigned(1540, 12), 1957 => to_unsigned(2144, 12), 1958 => to_unsigned(1706, 12), 1959 => to_unsigned(1913, 12), 1960 => to_unsigned(1501, 12), 1961 => to_unsigned(2357, 12), 1962 => to_unsigned(1725, 12), 1963 => to_unsigned(1865, 12), 1964 => to_unsigned(2441, 12), 1965 => to_unsigned(2297, 12), 1966 => to_unsigned(2509, 12), 1967 => to_unsigned(2384, 12), 1968 => to_unsigned(1806, 12), 1969 => to_unsigned(2490, 12), 1970 => to_unsigned(1842, 12), 1971 => to_unsigned(1364, 12), 1972 => to_unsigned(1976, 12), 1973 => to_unsigned(1730, 12), 1974 => to_unsigned(2027, 12), 1975 => to_unsigned(2747, 12), 1976 => to_unsigned(1882, 12), 1977 => to_unsigned(1536, 12), 1978 => to_unsigned(1488, 12), 1979 => to_unsigned(1557, 12), 1980 => to_unsigned(1800, 12), 1981 => to_unsigned(1568, 12), 1982 => to_unsigned(1564, 12), 1983 => to_unsigned(2042, 12), 1984 => to_unsigned(2164, 12), 1985 => to_unsigned(2250, 12), 1986 => to_unsigned(2224, 12), 1987 => to_unsigned(1943, 12), 1988 => to_unsigned(1704, 12), 1989 => to_unsigned(2501, 12), 1990 => to_unsigned(2381, 12), 1991 => to_unsigned(2185, 12), 1992 => to_unsigned(2362, 12), 1993 => to_unsigned(2015, 12), 1994 => to_unsigned(1845, 12), 1995 => to_unsigned(2180, 12), 1996 => to_unsigned(2186, 12), 1997 => to_unsigned(2496, 12), 1998 => to_unsigned(2475, 12), 1999 => to_unsigned(2093, 12), 2000 => to_unsigned(2096, 12), 2001 => to_unsigned(2006, 12), 2002 => to_unsigned(2168, 12), 2003 => to_unsigned(2238, 12), 2004 => to_unsigned(2235, 12), 2005 => to_unsigned(1874, 12), 2006 => to_unsigned(1927, 12), 2007 => to_unsigned(1410, 12), 2008 => to_unsigned(1990, 12), 2009 => to_unsigned(2352, 12), 2010 => to_unsigned(1942, 12), 2011 => to_unsigned(1388, 12), 2012 => to_unsigned(2485, 12), 2013 => to_unsigned(2091, 12), 2014 => to_unsigned(2294, 12), 2015 => to_unsigned(1623, 12), 2016 => to_unsigned(1960, 12), 2017 => to_unsigned(1720, 12), 2018 => to_unsigned(2001, 12), 2019 => to_unsigned(2468, 12), 2020 => to_unsigned(2012, 12), 2021 => to_unsigned(1671, 12), 2022 => to_unsigned(1590, 12), 2023 => to_unsigned(1765, 12), 2024 => to_unsigned(2517, 12), 2025 => to_unsigned(1777, 12), 2026 => to_unsigned(2661, 12), 2027 => to_unsigned(2102, 12), 2028 => to_unsigned(2293, 12), 2029 => to_unsigned(2459, 12), 2030 => to_unsigned(2506, 12), 2031 => to_unsigned(2143, 12), 2032 => to_unsigned(2379, 12), 2033 => to_unsigned(2592, 12), 2034 => to_unsigned(1379, 12), 2035 => to_unsigned(1884, 12), 2036 => to_unsigned(1745, 12), 2037 => to_unsigned(1957, 12), 2038 => to_unsigned(1820, 12), 2039 => to_unsigned(1980, 12), 2040 => to_unsigned(2355, 12), 2041 => to_unsigned(2190, 12), 2042 => to_unsigned(2337, 12), 2043 => to_unsigned(1802, 12), 2044 => to_unsigned(2177, 12), 2045 => to_unsigned(1967, 12), 2046 => to_unsigned(2458, 12), 2047 => to_unsigned(1485, 12)),
        2 => (0 => to_unsigned(2541, 12), 1 => to_unsigned(2211, 12), 2 => to_unsigned(2253, 12), 3 => to_unsigned(1983, 12), 4 => to_unsigned(1895, 12), 5 => to_unsigned(1797, 12), 6 => to_unsigned(2129, 12), 7 => to_unsigned(1925, 12), 8 => to_unsigned(2652, 12), 9 => to_unsigned(2042, 12), 10 => to_unsigned(1654, 12), 11 => to_unsigned(2230, 12), 12 => to_unsigned(2059, 12), 13 => to_unsigned(1965, 12), 14 => to_unsigned(2329, 12), 15 => to_unsigned(2093, 12), 16 => to_unsigned(2220, 12), 17 => to_unsigned(2161, 12), 18 => to_unsigned(1740, 12), 19 => to_unsigned(2612, 12), 20 => to_unsigned(1977, 12), 21 => to_unsigned(1747, 12), 22 => to_unsigned(1895, 12), 23 => to_unsigned(1899, 12), 24 => to_unsigned(1871, 12), 25 => to_unsigned(1562, 12), 26 => to_unsigned(2575, 12), 27 => to_unsigned(2628, 12), 28 => to_unsigned(2347, 12), 29 => to_unsigned(1926, 12), 30 => to_unsigned(1373, 12), 31 => to_unsigned(1914, 12), 32 => to_unsigned(2064, 12), 33 => to_unsigned(2009, 12), 34 => to_unsigned(2290, 12), 35 => to_unsigned(1591, 12), 36 => to_unsigned(2080, 12), 37 => to_unsigned(1783, 12), 38 => to_unsigned(1361, 12), 39 => to_unsigned(1579, 12), 40 => to_unsigned(1789, 12), 41 => to_unsigned(1695, 12), 42 => to_unsigned(1451, 12), 43 => to_unsigned(1844, 12), 44 => to_unsigned(2217, 12), 45 => to_unsigned(2256, 12), 46 => to_unsigned(2722, 12), 47 => to_unsigned(2147, 12), 48 => to_unsigned(2371, 12), 49 => to_unsigned(2464, 12), 50 => to_unsigned(2648, 12), 51 => to_unsigned(1802, 12), 52 => to_unsigned(1713, 12), 53 => to_unsigned(1441, 12), 54 => to_unsigned(2194, 12), 55 => to_unsigned(2070, 12), 56 => to_unsigned(1611, 12), 57 => to_unsigned(1473, 12), 58 => to_unsigned(2463, 12), 59 => to_unsigned(2281, 12), 60 => to_unsigned(2346, 12), 61 => to_unsigned(2344, 12), 62 => to_unsigned(1516, 12), 63 => to_unsigned(1787, 12), 64 => to_unsigned(2120, 12), 65 => to_unsigned(1983, 12), 66 => to_unsigned(1155, 12), 67 => to_unsigned(1980, 12), 68 => to_unsigned(2327, 12), 69 => to_unsigned(2429, 12), 70 => to_unsigned(2242, 12), 71 => to_unsigned(2412, 12), 72 => to_unsigned(1913, 12), 73 => to_unsigned(2268, 12), 74 => to_unsigned(2010, 12), 75 => to_unsigned(2077, 12), 76 => to_unsigned(2096, 12), 77 => to_unsigned(2200, 12), 78 => to_unsigned(1914, 12), 79 => to_unsigned(2178, 12), 80 => to_unsigned(1545, 12), 81 => to_unsigned(2101, 12), 82 => to_unsigned(2112, 12), 83 => to_unsigned(2431, 12), 84 => to_unsigned(1599, 12), 85 => to_unsigned(1928, 12), 86 => to_unsigned(2337, 12), 87 => to_unsigned(1855, 12), 88 => to_unsigned(2286, 12), 89 => to_unsigned(1385, 12), 90 => to_unsigned(2047, 12), 91 => to_unsigned(2285, 12), 92 => to_unsigned(2583, 12), 93 => to_unsigned(2080, 12), 94 => to_unsigned(1977, 12), 95 => to_unsigned(1503, 12), 96 => to_unsigned(1765, 12), 97 => to_unsigned(2608, 12), 98 => to_unsigned(2923, 12), 99 => to_unsigned(2136, 12), 100 => to_unsigned(2089, 12), 101 => to_unsigned(2657, 12), 102 => to_unsigned(1344, 12), 103 => to_unsigned(2434, 12), 104 => to_unsigned(3241, 12), 105 => to_unsigned(2160, 12), 106 => to_unsigned(1684, 12), 107 => to_unsigned(2447, 12), 108 => to_unsigned(1191, 12), 109 => to_unsigned(2335, 12), 110 => to_unsigned(2383, 12), 111 => to_unsigned(1826, 12), 112 => to_unsigned(2596, 12), 113 => to_unsigned(1896, 12), 114 => to_unsigned(1667, 12), 115 => to_unsigned(1646, 12), 116 => to_unsigned(1767, 12), 117 => to_unsigned(2277, 12), 118 => to_unsigned(2020, 12), 119 => to_unsigned(2147, 12), 120 => to_unsigned(2146, 12), 121 => to_unsigned(2859, 12), 122 => to_unsigned(1999, 12), 123 => to_unsigned(1870, 12), 124 => to_unsigned(1864, 12), 125 => to_unsigned(2876, 12), 126 => to_unsigned(2245, 12), 127 => to_unsigned(2045, 12), 128 => to_unsigned(2279, 12), 129 => to_unsigned(2545, 12), 130 => to_unsigned(1605, 12), 131 => to_unsigned(2358, 12), 132 => to_unsigned(2748, 12), 133 => to_unsigned(1794, 12), 134 => to_unsigned(1477, 12), 135 => to_unsigned(1863, 12), 136 => to_unsigned(2186, 12), 137 => to_unsigned(1859, 12), 138 => to_unsigned(1470, 12), 139 => to_unsigned(1666, 12), 140 => to_unsigned(2914, 12), 141 => to_unsigned(2270, 12), 142 => to_unsigned(2121, 12), 143 => to_unsigned(2326, 12), 144 => to_unsigned(1429, 12), 145 => to_unsigned(1502, 12), 146 => to_unsigned(1772, 12), 147 => to_unsigned(1976, 12), 148 => to_unsigned(2172, 12), 149 => to_unsigned(2103, 12), 150 => to_unsigned(1973, 12), 151 => to_unsigned(1790, 12), 152 => to_unsigned(2691, 12), 153 => to_unsigned(1660, 12), 154 => to_unsigned(2169, 12), 155 => to_unsigned(1198, 12), 156 => to_unsigned(2494, 12), 157 => to_unsigned(2571, 12), 158 => to_unsigned(2241, 12), 159 => to_unsigned(1785, 12), 160 => to_unsigned(2686, 12), 161 => to_unsigned(2042, 12), 162 => to_unsigned(1659, 12), 163 => to_unsigned(1891, 12), 164 => to_unsigned(1695, 12), 165 => to_unsigned(1904, 12), 166 => to_unsigned(2197, 12), 167 => to_unsigned(2414, 12), 168 => to_unsigned(2582, 12), 169 => to_unsigned(2383, 12), 170 => to_unsigned(1679, 12), 171 => to_unsigned(1499, 12), 172 => to_unsigned(1874, 12), 173 => to_unsigned(1682, 12), 174 => to_unsigned(1851, 12), 175 => to_unsigned(1685, 12), 176 => to_unsigned(1906, 12), 177 => to_unsigned(1636, 12), 178 => to_unsigned(1540, 12), 179 => to_unsigned(2376, 12), 180 => to_unsigned(1838, 12), 181 => to_unsigned(1967, 12), 182 => to_unsigned(2073, 12), 183 => to_unsigned(2120, 12), 184 => to_unsigned(2205, 12), 185 => to_unsigned(2241, 12), 186 => to_unsigned(1677, 12), 187 => to_unsigned(2803, 12), 188 => to_unsigned(792, 12), 189 => to_unsigned(2221, 12), 190 => to_unsigned(1665, 12), 191 => to_unsigned(2540, 12), 192 => to_unsigned(2001, 12), 193 => to_unsigned(2358, 12), 194 => to_unsigned(2531, 12), 195 => to_unsigned(1757, 12), 196 => to_unsigned(2150, 12), 197 => to_unsigned(2152, 12), 198 => to_unsigned(2043, 12), 199 => to_unsigned(1936, 12), 200 => to_unsigned(1396, 12), 201 => to_unsigned(1130, 12), 202 => to_unsigned(2968, 12), 203 => to_unsigned(2219, 12), 204 => to_unsigned(2445, 12), 205 => to_unsigned(1742, 12), 206 => to_unsigned(2183, 12), 207 => to_unsigned(1689, 12), 208 => to_unsigned(2305, 12), 209 => to_unsigned(2412, 12), 210 => to_unsigned(1559, 12), 211 => to_unsigned(1998, 12), 212 => to_unsigned(2111, 12), 213 => to_unsigned(827, 12), 214 => to_unsigned(2294, 12), 215 => to_unsigned(2193, 12), 216 => to_unsigned(1726, 12), 217 => to_unsigned(2104, 12), 218 => to_unsigned(1861, 12), 219 => to_unsigned(2145, 12), 220 => to_unsigned(2258, 12), 221 => to_unsigned(1031, 12), 222 => to_unsigned(2084, 12), 223 => to_unsigned(2811, 12), 224 => to_unsigned(2111, 12), 225 => to_unsigned(2000, 12), 226 => to_unsigned(2004, 12), 227 => to_unsigned(1585, 12), 228 => to_unsigned(2383, 12), 229 => to_unsigned(2669, 12), 230 => to_unsigned(2069, 12), 231 => to_unsigned(2240, 12), 232 => to_unsigned(1747, 12), 233 => to_unsigned(2629, 12), 234 => to_unsigned(1802, 12), 235 => to_unsigned(2717, 12), 236 => to_unsigned(1454, 12), 237 => to_unsigned(1934, 12), 238 => to_unsigned(2049, 12), 239 => to_unsigned(2011, 12), 240 => to_unsigned(2005, 12), 241 => to_unsigned(2005, 12), 242 => to_unsigned(1899, 12), 243 => to_unsigned(1163, 12), 244 => to_unsigned(2293, 12), 245 => to_unsigned(1546, 12), 246 => to_unsigned(2357, 12), 247 => to_unsigned(2441, 12), 248 => to_unsigned(2198, 12), 249 => to_unsigned(2161, 12), 250 => to_unsigned(1926, 12), 251 => to_unsigned(1738, 12), 252 => to_unsigned(2541, 12), 253 => to_unsigned(1759, 12), 254 => to_unsigned(2055, 12), 255 => to_unsigned(1832, 12), 256 => to_unsigned(2865, 12), 257 => to_unsigned(2748, 12), 258 => to_unsigned(2462, 12), 259 => to_unsigned(2402, 12), 260 => to_unsigned(2080, 12), 261 => to_unsigned(2659, 12), 262 => to_unsigned(3042, 12), 263 => to_unsigned(1578, 12), 264 => to_unsigned(1749, 12), 265 => to_unsigned(2102, 12), 266 => to_unsigned(1840, 12), 267 => to_unsigned(2870, 12), 268 => to_unsigned(2353, 12), 269 => to_unsigned(2471, 12), 270 => to_unsigned(1924, 12), 271 => to_unsigned(1570, 12), 272 => to_unsigned(2176, 12), 273 => to_unsigned(2696, 12), 274 => to_unsigned(2264, 12), 275 => to_unsigned(2744, 12), 276 => to_unsigned(1924, 12), 277 => to_unsigned(1747, 12), 278 => to_unsigned(2848, 12), 279 => to_unsigned(1723, 12), 280 => to_unsigned(2509, 12), 281 => to_unsigned(2207, 12), 282 => to_unsigned(1842, 12), 283 => to_unsigned(2457, 12), 284 => to_unsigned(2343, 12), 285 => to_unsigned(1747, 12), 286 => to_unsigned(1165, 12), 287 => to_unsigned(1955, 12), 288 => to_unsigned(1861, 12), 289 => to_unsigned(1899, 12), 290 => to_unsigned(1365, 12), 291 => to_unsigned(3295, 12), 292 => to_unsigned(1848, 12), 293 => to_unsigned(1356, 12), 294 => to_unsigned(2191, 12), 295 => to_unsigned(2053, 12), 296 => to_unsigned(1969, 12), 297 => to_unsigned(1681, 12), 298 => to_unsigned(2393, 12), 299 => to_unsigned(2264, 12), 300 => to_unsigned(1725, 12), 301 => to_unsigned(2128, 12), 302 => to_unsigned(2195, 12), 303 => to_unsigned(2816, 12), 304 => to_unsigned(1400, 12), 305 => to_unsigned(2309, 12), 306 => to_unsigned(2354, 12), 307 => to_unsigned(1621, 12), 308 => to_unsigned(1821, 12), 309 => to_unsigned(1451, 12), 310 => to_unsigned(1463, 12), 311 => to_unsigned(2629, 12), 312 => to_unsigned(2606, 12), 313 => to_unsigned(1681, 12), 314 => to_unsigned(1978, 12), 315 => to_unsigned(2069, 12), 316 => to_unsigned(2565, 12), 317 => to_unsigned(2482, 12), 318 => to_unsigned(2180, 12), 319 => to_unsigned(2174, 12), 320 => to_unsigned(1840, 12), 321 => to_unsigned(2008, 12), 322 => to_unsigned(1405, 12), 323 => to_unsigned(2797, 12), 324 => to_unsigned(1161, 12), 325 => to_unsigned(2692, 12), 326 => to_unsigned(2637, 12), 327 => to_unsigned(2149, 12), 328 => to_unsigned(1806, 12), 329 => to_unsigned(2028, 12), 330 => to_unsigned(2042, 12), 331 => to_unsigned(1707, 12), 332 => to_unsigned(1644, 12), 333 => to_unsigned(1801, 12), 334 => to_unsigned(1803, 12), 335 => to_unsigned(1930, 12), 336 => to_unsigned(1721, 12), 337 => to_unsigned(2437, 12), 338 => to_unsigned(2162, 12), 339 => to_unsigned(2204, 12), 340 => to_unsigned(2346, 12), 341 => to_unsigned(1894, 12), 342 => to_unsigned(2446, 12), 343 => to_unsigned(2430, 12), 344 => to_unsigned(2356, 12), 345 => to_unsigned(2049, 12), 346 => to_unsigned(1914, 12), 347 => to_unsigned(2657, 12), 348 => to_unsigned(1382, 12), 349 => to_unsigned(1935, 12), 350 => to_unsigned(1844, 12), 351 => to_unsigned(1694, 12), 352 => to_unsigned(2288, 12), 353 => to_unsigned(1738, 12), 354 => to_unsigned(2556, 12), 355 => to_unsigned(2059, 12), 356 => to_unsigned(1644, 12), 357 => to_unsigned(1914, 12), 358 => to_unsigned(2085, 12), 359 => to_unsigned(2215, 12), 360 => to_unsigned(1561, 12), 361 => to_unsigned(1746, 12), 362 => to_unsigned(2190, 12), 363 => to_unsigned(2157, 12), 364 => to_unsigned(2207, 12), 365 => to_unsigned(2707, 12), 366 => to_unsigned(1980, 12), 367 => to_unsigned(1539, 12), 368 => to_unsigned(1651, 12), 369 => to_unsigned(1929, 12), 370 => to_unsigned(2324, 12), 371 => to_unsigned(1847, 12), 372 => to_unsigned(2467, 12), 373 => to_unsigned(2496, 12), 374 => to_unsigned(1555, 12), 375 => to_unsigned(1611, 12), 376 => to_unsigned(1959, 12), 377 => to_unsigned(1977, 12), 378 => to_unsigned(1642, 12), 379 => to_unsigned(2443, 12), 380 => to_unsigned(2264, 12), 381 => to_unsigned(1688, 12), 382 => to_unsigned(2008, 12), 383 => to_unsigned(1892, 12), 384 => to_unsigned(2147, 12), 385 => to_unsigned(1230, 12), 386 => to_unsigned(1939, 12), 387 => to_unsigned(2519, 12), 388 => to_unsigned(2686, 12), 389 => to_unsigned(1335, 12), 390 => to_unsigned(2373, 12), 391 => to_unsigned(2290, 12), 392 => to_unsigned(1950, 12), 393 => to_unsigned(1912, 12), 394 => to_unsigned(1495, 12), 395 => to_unsigned(2055, 12), 396 => to_unsigned(1751, 12), 397 => to_unsigned(2362, 12), 398 => to_unsigned(2224, 12), 399 => to_unsigned(1875, 12), 400 => to_unsigned(2257, 12), 401 => to_unsigned(2996, 12), 402 => to_unsigned(2298, 12), 403 => to_unsigned(1792, 12), 404 => to_unsigned(2383, 12), 405 => to_unsigned(2136, 12), 406 => to_unsigned(1720, 12), 407 => to_unsigned(2043, 12), 408 => to_unsigned(1707, 12), 409 => to_unsigned(2012, 12), 410 => to_unsigned(2150, 12), 411 => to_unsigned(1558, 12), 412 => to_unsigned(2169, 12), 413 => to_unsigned(2132, 12), 414 => to_unsigned(2194, 12), 415 => to_unsigned(2344, 12), 416 => to_unsigned(2374, 12), 417 => to_unsigned(2603, 12), 418 => to_unsigned(2473, 12), 419 => to_unsigned(1332, 12), 420 => to_unsigned(2694, 12), 421 => to_unsigned(1968, 12), 422 => to_unsigned(1815, 12), 423 => to_unsigned(1800, 12), 424 => to_unsigned(2075, 12), 425 => to_unsigned(2259, 12), 426 => to_unsigned(2472, 12), 427 => to_unsigned(1815, 12), 428 => to_unsigned(2455, 12), 429 => to_unsigned(1665, 12), 430 => to_unsigned(1844, 12), 431 => to_unsigned(1494, 12), 432 => to_unsigned(2045, 12), 433 => to_unsigned(2635, 12), 434 => to_unsigned(2247, 12), 435 => to_unsigned(2455, 12), 436 => to_unsigned(1883, 12), 437 => to_unsigned(2005, 12), 438 => to_unsigned(1564, 12), 439 => to_unsigned(1692, 12), 440 => to_unsigned(2048, 12), 441 => to_unsigned(1939, 12), 442 => to_unsigned(2430, 12), 443 => to_unsigned(1914, 12), 444 => to_unsigned(2519, 12), 445 => to_unsigned(2033, 12), 446 => to_unsigned(1997, 12), 447 => to_unsigned(2277, 12), 448 => to_unsigned(1716, 12), 449 => to_unsigned(2410, 12), 450 => to_unsigned(1990, 12), 451 => to_unsigned(1926, 12), 452 => to_unsigned(1906, 12), 453 => to_unsigned(2418, 12), 454 => to_unsigned(2067, 12), 455 => to_unsigned(1800, 12), 456 => to_unsigned(1068, 12), 457 => to_unsigned(1946, 12), 458 => to_unsigned(2149, 12), 459 => to_unsigned(2386, 12), 460 => to_unsigned(1593, 12), 461 => to_unsigned(2189, 12), 462 => to_unsigned(2042, 12), 463 => to_unsigned(1841, 12), 464 => to_unsigned(1647, 12), 465 => to_unsigned(1557, 12), 466 => to_unsigned(1553, 12), 467 => to_unsigned(2464, 12), 468 => to_unsigned(2294, 12), 469 => to_unsigned(1550, 12), 470 => to_unsigned(2329, 12), 471 => to_unsigned(2317, 12), 472 => to_unsigned(2543, 12), 473 => to_unsigned(3199, 12), 474 => to_unsigned(1823, 12), 475 => to_unsigned(2491, 12), 476 => to_unsigned(1804, 12), 477 => to_unsigned(2416, 12), 478 => to_unsigned(1545, 12), 479 => to_unsigned(1988, 12), 480 => to_unsigned(2392, 12), 481 => to_unsigned(3006, 12), 482 => to_unsigned(1560, 12), 483 => to_unsigned(2255, 12), 484 => to_unsigned(2392, 12), 485 => to_unsigned(1816, 12), 486 => to_unsigned(1855, 12), 487 => to_unsigned(2186, 12), 488 => to_unsigned(2011, 12), 489 => to_unsigned(2706, 12), 490 => to_unsigned(1795, 12), 491 => to_unsigned(1860, 12), 492 => to_unsigned(2530, 12), 493 => to_unsigned(2063, 12), 494 => to_unsigned(2144, 12), 495 => to_unsigned(1777, 12), 496 => to_unsigned(2640, 12), 497 => to_unsigned(2493, 12), 498 => to_unsigned(2385, 12), 499 => to_unsigned(1735, 12), 500 => to_unsigned(1706, 12), 501 => to_unsigned(2182, 12), 502 => to_unsigned(1773, 12), 503 => to_unsigned(1748, 12), 504 => to_unsigned(1704, 12), 505 => to_unsigned(2561, 12), 506 => to_unsigned(2135, 12), 507 => to_unsigned(2724, 12), 508 => to_unsigned(2384, 12), 509 => to_unsigned(2057, 12), 510 => to_unsigned(2029, 12), 511 => to_unsigned(2230, 12), 512 => to_unsigned(1649, 12), 513 => to_unsigned(1729, 12), 514 => to_unsigned(2407, 12), 515 => to_unsigned(1498, 12), 516 => to_unsigned(1063, 12), 517 => to_unsigned(2344, 12), 518 => to_unsigned(2018, 12), 519 => to_unsigned(1553, 12), 520 => to_unsigned(2285, 12), 521 => to_unsigned(1984, 12), 522 => to_unsigned(1556, 12), 523 => to_unsigned(1414, 12), 524 => to_unsigned(1886, 12), 525 => to_unsigned(1656, 12), 526 => to_unsigned(1527, 12), 527 => to_unsigned(1643, 12), 528 => to_unsigned(1887, 12), 529 => to_unsigned(1929, 12), 530 => to_unsigned(1996, 12), 531 => to_unsigned(2460, 12), 532 => to_unsigned(2593, 12), 533 => to_unsigned(1917, 12), 534 => to_unsigned(1932, 12), 535 => to_unsigned(1314, 12), 536 => to_unsigned(2652, 12), 537 => to_unsigned(2494, 12), 538 => to_unsigned(2482, 12), 539 => to_unsigned(1913, 12), 540 => to_unsigned(1696, 12), 541 => to_unsigned(2430, 12), 542 => to_unsigned(1807, 12), 543 => to_unsigned(1952, 12), 544 => to_unsigned(1692, 12), 545 => to_unsigned(2086, 12), 546 => to_unsigned(1662, 12), 547 => to_unsigned(1991, 12), 548 => to_unsigned(2182, 12), 549 => to_unsigned(2243, 12), 550 => to_unsigned(2433, 12), 551 => to_unsigned(2279, 12), 552 => to_unsigned(2238, 12), 553 => to_unsigned(1542, 12), 554 => to_unsigned(1718, 12), 555 => to_unsigned(2345, 12), 556 => to_unsigned(2246, 12), 557 => to_unsigned(2490, 12), 558 => to_unsigned(2568, 12), 559 => to_unsigned(2322, 12), 560 => to_unsigned(1588, 12), 561 => to_unsigned(2681, 12), 562 => to_unsigned(2579, 12), 563 => to_unsigned(2070, 12), 564 => to_unsigned(1502, 12), 565 => to_unsigned(1475, 12), 566 => to_unsigned(2337, 12), 567 => to_unsigned(2218, 12), 568 => to_unsigned(2043, 12), 569 => to_unsigned(1685, 12), 570 => to_unsigned(1550, 12), 571 => to_unsigned(1787, 12), 572 => to_unsigned(1389, 12), 573 => to_unsigned(2016, 12), 574 => to_unsigned(1957, 12), 575 => to_unsigned(1767, 12), 576 => to_unsigned(2369, 12), 577 => to_unsigned(1544, 12), 578 => to_unsigned(2668, 12), 579 => to_unsigned(2310, 12), 580 => to_unsigned(2249, 12), 581 => to_unsigned(1726, 12), 582 => to_unsigned(1997, 12), 583 => to_unsigned(2480, 12), 584 => to_unsigned(1465, 12), 585 => to_unsigned(1876, 12), 586 => to_unsigned(1799, 12), 587 => to_unsigned(1848, 12), 588 => to_unsigned(1634, 12), 589 => to_unsigned(1715, 12), 590 => to_unsigned(2001, 12), 591 => to_unsigned(2253, 12), 592 => to_unsigned(1902, 12), 593 => to_unsigned(1878, 12), 594 => to_unsigned(1842, 12), 595 => to_unsigned(1402, 12), 596 => to_unsigned(1395, 12), 597 => to_unsigned(1731, 12), 598 => to_unsigned(2248, 12), 599 => to_unsigned(2337, 12), 600 => to_unsigned(1687, 12), 601 => to_unsigned(1803, 12), 602 => to_unsigned(1671, 12), 603 => to_unsigned(1643, 12), 604 => to_unsigned(1902, 12), 605 => to_unsigned(1627, 12), 606 => to_unsigned(2395, 12), 607 => to_unsigned(2080, 12), 608 => to_unsigned(2058, 12), 609 => to_unsigned(2464, 12), 610 => to_unsigned(2137, 12), 611 => to_unsigned(1956, 12), 612 => to_unsigned(2080, 12), 613 => to_unsigned(2602, 12), 614 => to_unsigned(1465, 12), 615 => to_unsigned(2418, 12), 616 => to_unsigned(1749, 12), 617 => to_unsigned(1806, 12), 618 => to_unsigned(2672, 12), 619 => to_unsigned(1982, 12), 620 => to_unsigned(2116, 12), 621 => to_unsigned(1981, 12), 622 => to_unsigned(2147, 12), 623 => to_unsigned(2146, 12), 624 => to_unsigned(1459, 12), 625 => to_unsigned(1446, 12), 626 => to_unsigned(2182, 12), 627 => to_unsigned(1708, 12), 628 => to_unsigned(2302, 12), 629 => to_unsigned(2246, 12), 630 => to_unsigned(1934, 12), 631 => to_unsigned(1999, 12), 632 => to_unsigned(2356, 12), 633 => to_unsigned(1870, 12), 634 => to_unsigned(2535, 12), 635 => to_unsigned(2410, 12), 636 => to_unsigned(1544, 12), 637 => to_unsigned(1972, 12), 638 => to_unsigned(2317, 12), 639 => to_unsigned(2066, 12), 640 => to_unsigned(2109, 12), 641 => to_unsigned(1768, 12), 642 => to_unsigned(1996, 12), 643 => to_unsigned(2227, 12), 644 => to_unsigned(1816, 12), 645 => to_unsigned(1370, 12), 646 => to_unsigned(1369, 12), 647 => to_unsigned(2325, 12), 648 => to_unsigned(1777, 12), 649 => to_unsigned(2128, 12), 650 => to_unsigned(2231, 12), 651 => to_unsigned(2697, 12), 652 => to_unsigned(2101, 12), 653 => to_unsigned(1905, 12), 654 => to_unsigned(2414, 12), 655 => to_unsigned(1947, 12), 656 => to_unsigned(2364, 12), 657 => to_unsigned(1612, 12), 658 => to_unsigned(2056, 12), 659 => to_unsigned(1928, 12), 660 => to_unsigned(1517, 12), 661 => to_unsigned(2443, 12), 662 => to_unsigned(1970, 12), 663 => to_unsigned(2340, 12), 664 => to_unsigned(2457, 12), 665 => to_unsigned(2208, 12), 666 => to_unsigned(2167, 12), 667 => to_unsigned(2221, 12), 668 => to_unsigned(1687, 12), 669 => to_unsigned(1606, 12), 670 => to_unsigned(2095, 12), 671 => to_unsigned(1721, 12), 672 => to_unsigned(2692, 12), 673 => to_unsigned(1636, 12), 674 => to_unsigned(2263, 12), 675 => to_unsigned(2071, 12), 676 => to_unsigned(1438, 12), 677 => to_unsigned(2871, 12), 678 => to_unsigned(2118, 12), 679 => to_unsigned(2046, 12), 680 => to_unsigned(2195, 12), 681 => to_unsigned(2653, 12), 682 => to_unsigned(2010, 12), 683 => to_unsigned(2743, 12), 684 => to_unsigned(1478, 12), 685 => to_unsigned(2664, 12), 686 => to_unsigned(2573, 12), 687 => to_unsigned(2064, 12), 688 => to_unsigned(2311, 12), 689 => to_unsigned(1768, 12), 690 => to_unsigned(1519, 12), 691 => to_unsigned(1144, 12), 692 => to_unsigned(1703, 12), 693 => to_unsigned(1989, 12), 694 => to_unsigned(1884, 12), 695 => to_unsigned(1776, 12), 696 => to_unsigned(2149, 12), 697 => to_unsigned(1628, 12), 698 => to_unsigned(2673, 12), 699 => to_unsigned(2398, 12), 700 => to_unsigned(1728, 12), 701 => to_unsigned(2121, 12), 702 => to_unsigned(1901, 12), 703 => to_unsigned(1786, 12), 704 => to_unsigned(1345, 12), 705 => to_unsigned(2751, 12), 706 => to_unsigned(1605, 12), 707 => to_unsigned(1523, 12), 708 => to_unsigned(2637, 12), 709 => to_unsigned(2658, 12), 710 => to_unsigned(1745, 12), 711 => to_unsigned(2371, 12), 712 => to_unsigned(1736, 12), 713 => to_unsigned(2429, 12), 714 => to_unsigned(2082, 12), 715 => to_unsigned(1377, 12), 716 => to_unsigned(2041, 12), 717 => to_unsigned(1996, 12), 718 => to_unsigned(2324, 12), 719 => to_unsigned(2498, 12), 720 => to_unsigned(2081, 12), 721 => to_unsigned(2951, 12), 722 => to_unsigned(2011, 12), 723 => to_unsigned(2546, 12), 724 => to_unsigned(2029, 12), 725 => to_unsigned(1069, 12), 726 => to_unsigned(1530, 12), 727 => to_unsigned(1728, 12), 728 => to_unsigned(1661, 12), 729 => to_unsigned(2044, 12), 730 => to_unsigned(1369, 12), 731 => to_unsigned(2884, 12), 732 => to_unsigned(1913, 12), 733 => to_unsigned(2701, 12), 734 => to_unsigned(2461, 12), 735 => to_unsigned(1989, 12), 736 => to_unsigned(1579, 12), 737 => to_unsigned(1841, 12), 738 => to_unsigned(1557, 12), 739 => to_unsigned(2547, 12), 740 => to_unsigned(1620, 12), 741 => to_unsigned(2032, 12), 742 => to_unsigned(1588, 12), 743 => to_unsigned(2195, 12), 744 => to_unsigned(2548, 12), 745 => to_unsigned(1731, 12), 746 => to_unsigned(2488, 12), 747 => to_unsigned(1876, 12), 748 => to_unsigned(2290, 12), 749 => to_unsigned(2260, 12), 750 => to_unsigned(1902, 12), 751 => to_unsigned(1939, 12), 752 => to_unsigned(2033, 12), 753 => to_unsigned(1463, 12), 754 => to_unsigned(2696, 12), 755 => to_unsigned(1978, 12), 756 => to_unsigned(1596, 12), 757 => to_unsigned(2099, 12), 758 => to_unsigned(2560, 12), 759 => to_unsigned(1999, 12), 760 => to_unsigned(2181, 12), 761 => to_unsigned(1785, 12), 762 => to_unsigned(2381, 12), 763 => to_unsigned(1106, 12), 764 => to_unsigned(1283, 12), 765 => to_unsigned(2649, 12), 766 => to_unsigned(2466, 12), 767 => to_unsigned(1482, 12), 768 => to_unsigned(1763, 12), 769 => to_unsigned(2237, 12), 770 => to_unsigned(1749, 12), 771 => to_unsigned(1505, 12), 772 => to_unsigned(1711, 12), 773 => to_unsigned(1835, 12), 774 => to_unsigned(2243, 12), 775 => to_unsigned(2094, 12), 776 => to_unsigned(2001, 12), 777 => to_unsigned(1902, 12), 778 => to_unsigned(1097, 12), 779 => to_unsigned(2164, 12), 780 => to_unsigned(2480, 12), 781 => to_unsigned(2306, 12), 782 => to_unsigned(2295, 12), 783 => to_unsigned(1760, 12), 784 => to_unsigned(2434, 12), 785 => to_unsigned(1921, 12), 786 => to_unsigned(2518, 12), 787 => to_unsigned(1910, 12), 788 => to_unsigned(1672, 12), 789 => to_unsigned(1346, 12), 790 => to_unsigned(2053, 12), 791 => to_unsigned(1894, 12), 792 => to_unsigned(2567, 12), 793 => to_unsigned(1866, 12), 794 => to_unsigned(2605, 12), 795 => to_unsigned(1451, 12), 796 => to_unsigned(2210, 12), 797 => to_unsigned(2142, 12), 798 => to_unsigned(2695, 12), 799 => to_unsigned(1364, 12), 800 => to_unsigned(1510, 12), 801 => to_unsigned(2049, 12), 802 => to_unsigned(1684, 12), 803 => to_unsigned(1671, 12), 804 => to_unsigned(1577, 12), 805 => to_unsigned(1503, 12), 806 => to_unsigned(1993, 12), 807 => to_unsigned(1656, 12), 808 => to_unsigned(2628, 12), 809 => to_unsigned(1841, 12), 810 => to_unsigned(1878, 12), 811 => to_unsigned(1793, 12), 812 => to_unsigned(2245, 12), 813 => to_unsigned(2037, 12), 814 => to_unsigned(1755, 12), 815 => to_unsigned(1864, 12), 816 => to_unsigned(1959, 12), 817 => to_unsigned(1977, 12), 818 => to_unsigned(2122, 12), 819 => to_unsigned(1637, 12), 820 => to_unsigned(2565, 12), 821 => to_unsigned(1897, 12), 822 => to_unsigned(1886, 12), 823 => to_unsigned(2009, 12), 824 => to_unsigned(2100, 12), 825 => to_unsigned(1922, 12), 826 => to_unsigned(2032, 12), 827 => to_unsigned(1635, 12), 828 => to_unsigned(2525, 12), 829 => to_unsigned(2083, 12), 830 => to_unsigned(1533, 12), 831 => to_unsigned(1506, 12), 832 => to_unsigned(2496, 12), 833 => to_unsigned(2040, 12), 834 => to_unsigned(2101, 12), 835 => to_unsigned(1247, 12), 836 => to_unsigned(1634, 12), 837 => to_unsigned(2052, 12), 838 => to_unsigned(2530, 12), 839 => to_unsigned(2133, 12), 840 => to_unsigned(2357, 12), 841 => to_unsigned(1713, 12), 842 => to_unsigned(2620, 12), 843 => to_unsigned(1809, 12), 844 => to_unsigned(2589, 12), 845 => to_unsigned(1938, 12), 846 => to_unsigned(1707, 12), 847 => to_unsigned(2061, 12), 848 => to_unsigned(1598, 12), 849 => to_unsigned(1952, 12), 850 => to_unsigned(2258, 12), 851 => to_unsigned(2365, 12), 852 => to_unsigned(2241, 12), 853 => to_unsigned(1849, 12), 854 => to_unsigned(2295, 12), 855 => to_unsigned(2186, 12), 856 => to_unsigned(2242, 12), 857 => to_unsigned(1810, 12), 858 => to_unsigned(2420, 12), 859 => to_unsigned(1690, 12), 860 => to_unsigned(2651, 12), 861 => to_unsigned(1569, 12), 862 => to_unsigned(1861, 12), 863 => to_unsigned(2339, 12), 864 => to_unsigned(1877, 12), 865 => to_unsigned(2247, 12), 866 => to_unsigned(2335, 12), 867 => to_unsigned(2180, 12), 868 => to_unsigned(1605, 12), 869 => to_unsigned(2391, 12), 870 => to_unsigned(1503, 12), 871 => to_unsigned(1574, 12), 872 => to_unsigned(1944, 12), 873 => to_unsigned(2398, 12), 874 => to_unsigned(1138, 12), 875 => to_unsigned(1697, 12), 876 => to_unsigned(1688, 12), 877 => to_unsigned(1713, 12), 878 => to_unsigned(2171, 12), 879 => to_unsigned(2039, 12), 880 => to_unsigned(1955, 12), 881 => to_unsigned(1859, 12), 882 => to_unsigned(2086, 12), 883 => to_unsigned(1358, 12), 884 => to_unsigned(1713, 12), 885 => to_unsigned(2287, 12), 886 => to_unsigned(1151, 12), 887 => to_unsigned(2434, 12), 888 => to_unsigned(1955, 12), 889 => to_unsigned(1976, 12), 890 => to_unsigned(2194, 12), 891 => to_unsigned(2429, 12), 892 => to_unsigned(2535, 12), 893 => to_unsigned(1826, 12), 894 => to_unsigned(1590, 12), 895 => to_unsigned(1962, 12), 896 => to_unsigned(2868, 12), 897 => to_unsigned(2060, 12), 898 => to_unsigned(1501, 12), 899 => to_unsigned(2480, 12), 900 => to_unsigned(1382, 12), 901 => to_unsigned(1698, 12), 902 => to_unsigned(1886, 12), 903 => to_unsigned(1804, 12), 904 => to_unsigned(1971, 12), 905 => to_unsigned(2511, 12), 906 => to_unsigned(1782, 12), 907 => to_unsigned(2050, 12), 908 => to_unsigned(2219, 12), 909 => to_unsigned(1935, 12), 910 => to_unsigned(2633, 12), 911 => to_unsigned(2064, 12), 912 => to_unsigned(1695, 12), 913 => to_unsigned(2928, 12), 914 => to_unsigned(2068, 12), 915 => to_unsigned(2369, 12), 916 => to_unsigned(1532, 12), 917 => to_unsigned(1475, 12), 918 => to_unsigned(2091, 12), 919 => to_unsigned(1485, 12), 920 => to_unsigned(2189, 12), 921 => to_unsigned(1651, 12), 922 => to_unsigned(2658, 12), 923 => to_unsigned(2168, 12), 924 => to_unsigned(1703, 12), 925 => to_unsigned(1543, 12), 926 => to_unsigned(2410, 12), 927 => to_unsigned(2429, 12), 928 => to_unsigned(1869, 12), 929 => to_unsigned(1959, 12), 930 => to_unsigned(1911, 12), 931 => to_unsigned(1841, 12), 932 => to_unsigned(2261, 12), 933 => to_unsigned(1807, 12), 934 => to_unsigned(2059, 12), 935 => to_unsigned(2007, 12), 936 => to_unsigned(2452, 12), 937 => to_unsigned(1752, 12), 938 => to_unsigned(1729, 12), 939 => to_unsigned(1931, 12), 940 => to_unsigned(2130, 12), 941 => to_unsigned(1577, 12), 942 => to_unsigned(1237, 12), 943 => to_unsigned(2894, 12), 944 => to_unsigned(1765, 12), 945 => to_unsigned(2588, 12), 946 => to_unsigned(1874, 12), 947 => to_unsigned(1517, 12), 948 => to_unsigned(1362, 12), 949 => to_unsigned(2046, 12), 950 => to_unsigned(1980, 12), 951 => to_unsigned(1630, 12), 952 => to_unsigned(2328, 12), 953 => to_unsigned(1931, 12), 954 => to_unsigned(2276, 12), 955 => to_unsigned(2493, 12), 956 => to_unsigned(2225, 12), 957 => to_unsigned(2047, 12), 958 => to_unsigned(2538, 12), 959 => to_unsigned(1785, 12), 960 => to_unsigned(2203, 12), 961 => to_unsigned(2047, 12), 962 => to_unsigned(2656, 12), 963 => to_unsigned(2440, 12), 964 => to_unsigned(2198, 12), 965 => to_unsigned(2295, 12), 966 => to_unsigned(1551, 12), 967 => to_unsigned(2469, 12), 968 => to_unsigned(2158, 12), 969 => to_unsigned(1367, 12), 970 => to_unsigned(2092, 12), 971 => to_unsigned(2157, 12), 972 => to_unsigned(2177, 12), 973 => to_unsigned(1375, 12), 974 => to_unsigned(1996, 12), 975 => to_unsigned(1763, 12), 976 => to_unsigned(2291, 12), 977 => to_unsigned(2181, 12), 978 => to_unsigned(2471, 12), 979 => to_unsigned(2415, 12), 980 => to_unsigned(1944, 12), 981 => to_unsigned(2100, 12), 982 => to_unsigned(1443, 12), 983 => to_unsigned(1822, 12), 984 => to_unsigned(1985, 12), 985 => to_unsigned(2395, 12), 986 => to_unsigned(2287, 12), 987 => to_unsigned(2132, 12), 988 => to_unsigned(1595, 12), 989 => to_unsigned(2265, 12), 990 => to_unsigned(2380, 12), 991 => to_unsigned(1850, 12), 992 => to_unsigned(1222, 12), 993 => to_unsigned(1641, 12), 994 => to_unsigned(2482, 12), 995 => to_unsigned(1892, 12), 996 => to_unsigned(2015, 12), 997 => to_unsigned(1885, 12), 998 => to_unsigned(1566, 12), 999 => to_unsigned(2760, 12), 1000 => to_unsigned(2777, 12), 1001 => to_unsigned(2540, 12), 1002 => to_unsigned(1994, 12), 1003 => to_unsigned(2076, 12), 1004 => to_unsigned(1537, 12), 1005 => to_unsigned(2185, 12), 1006 => to_unsigned(2087, 12), 1007 => to_unsigned(1761, 12), 1008 => to_unsigned(2203, 12), 1009 => to_unsigned(1723, 12), 1010 => to_unsigned(1936, 12), 1011 => to_unsigned(2103, 12), 1012 => to_unsigned(1520, 12), 1013 => to_unsigned(2240, 12), 1014 => to_unsigned(1812, 12), 1015 => to_unsigned(1998, 12), 1016 => to_unsigned(1582, 12), 1017 => to_unsigned(1171, 12), 1018 => to_unsigned(2144, 12), 1019 => to_unsigned(2264, 12), 1020 => to_unsigned(1221, 12), 1021 => to_unsigned(2277, 12), 1022 => to_unsigned(1775, 12), 1023 => to_unsigned(1703, 12), 1024 => to_unsigned(2080, 12), 1025 => to_unsigned(2001, 12), 1026 => to_unsigned(1869, 12), 1027 => to_unsigned(2297, 12), 1028 => to_unsigned(2181, 12), 1029 => to_unsigned(2473, 12), 1030 => to_unsigned(1828, 12), 1031 => to_unsigned(2401, 12), 1032 => to_unsigned(2140, 12), 1033 => to_unsigned(2534, 12), 1034 => to_unsigned(1755, 12), 1035 => to_unsigned(2172, 12), 1036 => to_unsigned(1134, 12), 1037 => to_unsigned(1899, 12), 1038 => to_unsigned(1946, 12), 1039 => to_unsigned(2761, 12), 1040 => to_unsigned(2348, 12), 1041 => to_unsigned(1343, 12), 1042 => to_unsigned(1534, 12), 1043 => to_unsigned(1849, 12), 1044 => to_unsigned(1323, 12), 1045 => to_unsigned(1632, 12), 1046 => to_unsigned(1487, 12), 1047 => to_unsigned(2293, 12), 1048 => to_unsigned(2119, 12), 1049 => to_unsigned(1726, 12), 1050 => to_unsigned(2034, 12), 1051 => to_unsigned(1939, 12), 1052 => to_unsigned(1486, 12), 1053 => to_unsigned(1632, 12), 1054 => to_unsigned(1970, 12), 1055 => to_unsigned(1836, 12), 1056 => to_unsigned(2422, 12), 1057 => to_unsigned(1923, 12), 1058 => to_unsigned(2081, 12), 1059 => to_unsigned(2721, 12), 1060 => to_unsigned(1979, 12), 1061 => to_unsigned(2051, 12), 1062 => to_unsigned(1938, 12), 1063 => to_unsigned(2399, 12), 1064 => to_unsigned(2220, 12), 1065 => to_unsigned(2449, 12), 1066 => to_unsigned(2126, 12), 1067 => to_unsigned(2460, 12), 1068 => to_unsigned(2062, 12), 1069 => to_unsigned(2465, 12), 1070 => to_unsigned(2464, 12), 1071 => to_unsigned(2360, 12), 1072 => to_unsigned(1877, 12), 1073 => to_unsigned(2271, 12), 1074 => to_unsigned(1625, 12), 1075 => to_unsigned(1728, 12), 1076 => to_unsigned(2016, 12), 1077 => to_unsigned(2507, 12), 1078 => to_unsigned(2335, 12), 1079 => to_unsigned(1815, 12), 1080 => to_unsigned(1798, 12), 1081 => to_unsigned(1993, 12), 1082 => to_unsigned(1790, 12), 1083 => to_unsigned(1392, 12), 1084 => to_unsigned(1633, 12), 1085 => to_unsigned(1920, 12), 1086 => to_unsigned(2381, 12), 1087 => to_unsigned(2168, 12), 1088 => to_unsigned(2323, 12), 1089 => to_unsigned(1855, 12), 1090 => to_unsigned(1627, 12), 1091 => to_unsigned(2003, 12), 1092 => to_unsigned(1961, 12), 1093 => to_unsigned(2567, 12), 1094 => to_unsigned(1513, 12), 1095 => to_unsigned(2167, 12), 1096 => to_unsigned(2316, 12), 1097 => to_unsigned(2414, 12), 1098 => to_unsigned(1937, 12), 1099 => to_unsigned(2092, 12), 1100 => to_unsigned(2000, 12), 1101 => to_unsigned(1990, 12), 1102 => to_unsigned(1873, 12), 1103 => to_unsigned(1862, 12), 1104 => to_unsigned(1999, 12), 1105 => to_unsigned(1862, 12), 1106 => to_unsigned(2023, 12), 1107 => to_unsigned(1627, 12), 1108 => to_unsigned(1750, 12), 1109 => to_unsigned(2802, 12), 1110 => to_unsigned(2279, 12), 1111 => to_unsigned(2967, 12), 1112 => to_unsigned(1817, 12), 1113 => to_unsigned(1408, 12), 1114 => to_unsigned(2125, 12), 1115 => to_unsigned(2135, 12), 1116 => to_unsigned(1699, 12), 1117 => to_unsigned(1954, 12), 1118 => to_unsigned(2383, 12), 1119 => to_unsigned(2442, 12), 1120 => to_unsigned(2167, 12), 1121 => to_unsigned(2341, 12), 1122 => to_unsigned(1834, 12), 1123 => to_unsigned(2072, 12), 1124 => to_unsigned(2125, 12), 1125 => to_unsigned(1807, 12), 1126 => to_unsigned(2311, 12), 1127 => to_unsigned(2252, 12), 1128 => to_unsigned(2246, 12), 1129 => to_unsigned(2094, 12), 1130 => to_unsigned(2140, 12), 1131 => to_unsigned(2202, 12), 1132 => to_unsigned(1311, 12), 1133 => to_unsigned(2400, 12), 1134 => to_unsigned(2071, 12), 1135 => to_unsigned(2272, 12), 1136 => to_unsigned(2472, 12), 1137 => to_unsigned(2091, 12), 1138 => to_unsigned(2366, 12), 1139 => to_unsigned(1807, 12), 1140 => to_unsigned(2855, 12), 1141 => to_unsigned(2361, 12), 1142 => to_unsigned(3158, 12), 1143 => to_unsigned(2697, 12), 1144 => to_unsigned(1942, 12), 1145 => to_unsigned(2158, 12), 1146 => to_unsigned(2145, 12), 1147 => to_unsigned(1623, 12), 1148 => to_unsigned(1838, 12), 1149 => to_unsigned(1922, 12), 1150 => to_unsigned(2740, 12), 1151 => to_unsigned(1774, 12), 1152 => to_unsigned(1871, 12), 1153 => to_unsigned(1837, 12), 1154 => to_unsigned(1891, 12), 1155 => to_unsigned(2139, 12), 1156 => to_unsigned(2654, 12), 1157 => to_unsigned(2175, 12), 1158 => to_unsigned(1738, 12), 1159 => to_unsigned(1685, 12), 1160 => to_unsigned(2469, 12), 1161 => to_unsigned(2323, 12), 1162 => to_unsigned(3126, 12), 1163 => to_unsigned(1767, 12), 1164 => to_unsigned(1437, 12), 1165 => to_unsigned(2034, 12), 1166 => to_unsigned(1766, 12), 1167 => to_unsigned(1762, 12), 1168 => to_unsigned(2136, 12), 1169 => to_unsigned(2078, 12), 1170 => to_unsigned(1930, 12), 1171 => to_unsigned(2426, 12), 1172 => to_unsigned(1984, 12), 1173 => to_unsigned(2838, 12), 1174 => to_unsigned(1658, 12), 1175 => to_unsigned(2116, 12), 1176 => to_unsigned(1502, 12), 1177 => to_unsigned(2335, 12), 1178 => to_unsigned(2344, 12), 1179 => to_unsigned(2585, 12), 1180 => to_unsigned(1742, 12), 1181 => to_unsigned(1866, 12), 1182 => to_unsigned(1846, 12), 1183 => to_unsigned(2232, 12), 1184 => to_unsigned(2539, 12), 1185 => to_unsigned(1908, 12), 1186 => to_unsigned(2708, 12), 1187 => to_unsigned(1178, 12), 1188 => to_unsigned(1930, 12), 1189 => to_unsigned(2362, 12), 1190 => to_unsigned(1994, 12), 1191 => to_unsigned(1776, 12), 1192 => to_unsigned(2269, 12), 1193 => to_unsigned(930, 12), 1194 => to_unsigned(2145, 12), 1195 => to_unsigned(2351, 12), 1196 => to_unsigned(1446, 12), 1197 => to_unsigned(2085, 12), 1198 => to_unsigned(3049, 12), 1199 => to_unsigned(1563, 12), 1200 => to_unsigned(1771, 12), 1201 => to_unsigned(2097, 12), 1202 => to_unsigned(2476, 12), 1203 => to_unsigned(2673, 12), 1204 => to_unsigned(2708, 12), 1205 => to_unsigned(2137, 12), 1206 => to_unsigned(1724, 12), 1207 => to_unsigned(1910, 12), 1208 => to_unsigned(1721, 12), 1209 => to_unsigned(2497, 12), 1210 => to_unsigned(2334, 12), 1211 => to_unsigned(1807, 12), 1212 => to_unsigned(1855, 12), 1213 => to_unsigned(1696, 12), 1214 => to_unsigned(2373, 12), 1215 => to_unsigned(2039, 12), 1216 => to_unsigned(1991, 12), 1217 => to_unsigned(2375, 12), 1218 => to_unsigned(2545, 12), 1219 => to_unsigned(2299, 12), 1220 => to_unsigned(1367, 12), 1221 => to_unsigned(1974, 12), 1222 => to_unsigned(1900, 12), 1223 => to_unsigned(2320, 12), 1224 => to_unsigned(1841, 12), 1225 => to_unsigned(1882, 12), 1226 => to_unsigned(1730, 12), 1227 => to_unsigned(1720, 12), 1228 => to_unsigned(2365, 12), 1229 => to_unsigned(2372, 12), 1230 => to_unsigned(1680, 12), 1231 => to_unsigned(1459, 12), 1232 => to_unsigned(2144, 12), 1233 => to_unsigned(1375, 12), 1234 => to_unsigned(1853, 12), 1235 => to_unsigned(1801, 12), 1236 => to_unsigned(2467, 12), 1237 => to_unsigned(2445, 12), 1238 => to_unsigned(1994, 12), 1239 => to_unsigned(2037, 12), 1240 => to_unsigned(2203, 12), 1241 => to_unsigned(1835, 12), 1242 => to_unsigned(1627, 12), 1243 => to_unsigned(2555, 12), 1244 => to_unsigned(2305, 12), 1245 => to_unsigned(2129, 12), 1246 => to_unsigned(2161, 12), 1247 => to_unsigned(1977, 12), 1248 => to_unsigned(1785, 12), 1249 => to_unsigned(2152, 12), 1250 => to_unsigned(2066, 12), 1251 => to_unsigned(1480, 12), 1252 => to_unsigned(1986, 12), 1253 => to_unsigned(2393, 12), 1254 => to_unsigned(1864, 12), 1255 => to_unsigned(1740, 12), 1256 => to_unsigned(2276, 12), 1257 => to_unsigned(2469, 12), 1258 => to_unsigned(1361, 12), 1259 => to_unsigned(1395, 12), 1260 => to_unsigned(1594, 12), 1261 => to_unsigned(1518, 12), 1262 => to_unsigned(2282, 12), 1263 => to_unsigned(2407, 12), 1264 => to_unsigned(1435, 12), 1265 => to_unsigned(2552, 12), 1266 => to_unsigned(2508, 12), 1267 => to_unsigned(2644, 12), 1268 => to_unsigned(1649, 12), 1269 => to_unsigned(1511, 12), 1270 => to_unsigned(1995, 12), 1271 => to_unsigned(1551, 12), 1272 => to_unsigned(1872, 12), 1273 => to_unsigned(2039, 12), 1274 => to_unsigned(1645, 12), 1275 => to_unsigned(2017, 12), 1276 => to_unsigned(1852, 12), 1277 => to_unsigned(2279, 12), 1278 => to_unsigned(2044, 12), 1279 => to_unsigned(2298, 12), 1280 => to_unsigned(2481, 12), 1281 => to_unsigned(2627, 12), 1282 => to_unsigned(1619, 12), 1283 => to_unsigned(2196, 12), 1284 => to_unsigned(1367, 12), 1285 => to_unsigned(1566, 12), 1286 => to_unsigned(2109, 12), 1287 => to_unsigned(2914, 12), 1288 => to_unsigned(2004, 12), 1289 => to_unsigned(2342, 12), 1290 => to_unsigned(1920, 12), 1291 => to_unsigned(1889, 12), 1292 => to_unsigned(2477, 12), 1293 => to_unsigned(1749, 12), 1294 => to_unsigned(1370, 12), 1295 => to_unsigned(2267, 12), 1296 => to_unsigned(2106, 12), 1297 => to_unsigned(1727, 12), 1298 => to_unsigned(2007, 12), 1299 => to_unsigned(2234, 12), 1300 => to_unsigned(1551, 12), 1301 => to_unsigned(1796, 12), 1302 => to_unsigned(1807, 12), 1303 => to_unsigned(2125, 12), 1304 => to_unsigned(2749, 12), 1305 => to_unsigned(1738, 12), 1306 => to_unsigned(2132, 12), 1307 => to_unsigned(2501, 12), 1308 => to_unsigned(2254, 12), 1309 => to_unsigned(1967, 12), 1310 => to_unsigned(1695, 12), 1311 => to_unsigned(2182, 12), 1312 => to_unsigned(2374, 12), 1313 => to_unsigned(2490, 12), 1314 => to_unsigned(1897, 12), 1315 => to_unsigned(1976, 12), 1316 => to_unsigned(2153, 12), 1317 => to_unsigned(1735, 12), 1318 => to_unsigned(2148, 12), 1319 => to_unsigned(1655, 12), 1320 => to_unsigned(1943, 12), 1321 => to_unsigned(1540, 12), 1322 => to_unsigned(1668, 12), 1323 => to_unsigned(1896, 12), 1324 => to_unsigned(2683, 12), 1325 => to_unsigned(2191, 12), 1326 => to_unsigned(2475, 12), 1327 => to_unsigned(2390, 12), 1328 => to_unsigned(1815, 12), 1329 => to_unsigned(2496, 12), 1330 => to_unsigned(2107, 12), 1331 => to_unsigned(1578, 12), 1332 => to_unsigned(2264, 12), 1333 => to_unsigned(2184, 12), 1334 => to_unsigned(2359, 12), 1335 => to_unsigned(2381, 12), 1336 => to_unsigned(2621, 12), 1337 => to_unsigned(1464, 12), 1338 => to_unsigned(1961, 12), 1339 => to_unsigned(2648, 12), 1340 => to_unsigned(1756, 12), 1341 => to_unsigned(2382, 12), 1342 => to_unsigned(2097, 12), 1343 => to_unsigned(2897, 12), 1344 => to_unsigned(2273, 12), 1345 => to_unsigned(2062, 12), 1346 => to_unsigned(2519, 12), 1347 => to_unsigned(2473, 12), 1348 => to_unsigned(2413, 12), 1349 => to_unsigned(1977, 12), 1350 => to_unsigned(2023, 12), 1351 => to_unsigned(1934, 12), 1352 => to_unsigned(1323, 12), 1353 => to_unsigned(1975, 12), 1354 => to_unsigned(2521, 12), 1355 => to_unsigned(2247, 12), 1356 => to_unsigned(2345, 12), 1357 => to_unsigned(2314, 12), 1358 => to_unsigned(2117, 12), 1359 => to_unsigned(2386, 12), 1360 => to_unsigned(2081, 12), 1361 => to_unsigned(1618, 12), 1362 => to_unsigned(2077, 12), 1363 => to_unsigned(2683, 12), 1364 => to_unsigned(2375, 12), 1365 => to_unsigned(1588, 12), 1366 => to_unsigned(2226, 12), 1367 => to_unsigned(2164, 12), 1368 => to_unsigned(1855, 12), 1369 => to_unsigned(2202, 12), 1370 => to_unsigned(1289, 12), 1371 => to_unsigned(2003, 12), 1372 => to_unsigned(1852, 12), 1373 => to_unsigned(2224, 12), 1374 => to_unsigned(1393, 12), 1375 => to_unsigned(2525, 12), 1376 => to_unsigned(2094, 12), 1377 => to_unsigned(2005, 12), 1378 => to_unsigned(2373, 12), 1379 => to_unsigned(2112, 12), 1380 => to_unsigned(1879, 12), 1381 => to_unsigned(1862, 12), 1382 => to_unsigned(1723, 12), 1383 => to_unsigned(2115, 12), 1384 => to_unsigned(1651, 12), 1385 => to_unsigned(1970, 12), 1386 => to_unsigned(2150, 12), 1387 => to_unsigned(1712, 12), 1388 => to_unsigned(2022, 12), 1389 => to_unsigned(2233, 12), 1390 => to_unsigned(1825, 12), 1391 => to_unsigned(2083, 12), 1392 => to_unsigned(2416, 12), 1393 => to_unsigned(1434, 12), 1394 => to_unsigned(2126, 12), 1395 => to_unsigned(1772, 12), 1396 => to_unsigned(2169, 12), 1397 => to_unsigned(2170, 12), 1398 => to_unsigned(1874, 12), 1399 => to_unsigned(1947, 12), 1400 => to_unsigned(1682, 12), 1401 => to_unsigned(2335, 12), 1402 => to_unsigned(1810, 12), 1403 => to_unsigned(2168, 12), 1404 => to_unsigned(2542, 12), 1405 => to_unsigned(2127, 12), 1406 => to_unsigned(2548, 12), 1407 => to_unsigned(2177, 12), 1408 => to_unsigned(2336, 12), 1409 => to_unsigned(1881, 12), 1410 => to_unsigned(1705, 12), 1411 => to_unsigned(1698, 12), 1412 => to_unsigned(2406, 12), 1413 => to_unsigned(2089, 12), 1414 => to_unsigned(1801, 12), 1415 => to_unsigned(2065, 12), 1416 => to_unsigned(1441, 12), 1417 => to_unsigned(2296, 12), 1418 => to_unsigned(2223, 12), 1419 => to_unsigned(2469, 12), 1420 => to_unsigned(2506, 12), 1421 => to_unsigned(2021, 12), 1422 => to_unsigned(1986, 12), 1423 => to_unsigned(2211, 12), 1424 => to_unsigned(1451, 12), 1425 => to_unsigned(2144, 12), 1426 => to_unsigned(1038, 12), 1427 => to_unsigned(1274, 12), 1428 => to_unsigned(2125, 12), 1429 => to_unsigned(2187, 12), 1430 => to_unsigned(1778, 12), 1431 => to_unsigned(1685, 12), 1432 => to_unsigned(1849, 12), 1433 => to_unsigned(2010, 12), 1434 => to_unsigned(2701, 12), 1435 => to_unsigned(1647, 12), 1436 => to_unsigned(2673, 12), 1437 => to_unsigned(1961, 12), 1438 => to_unsigned(1909, 12), 1439 => to_unsigned(1782, 12), 1440 => to_unsigned(1683, 12), 1441 => to_unsigned(1438, 12), 1442 => to_unsigned(1736, 12), 1443 => to_unsigned(1968, 12), 1444 => to_unsigned(2206, 12), 1445 => to_unsigned(2169, 12), 1446 => to_unsigned(2172, 12), 1447 => to_unsigned(1380, 12), 1448 => to_unsigned(1472, 12), 1449 => to_unsigned(2135, 12), 1450 => to_unsigned(2125, 12), 1451 => to_unsigned(2428, 12), 1452 => to_unsigned(2330, 12), 1453 => to_unsigned(2676, 12), 1454 => to_unsigned(1731, 12), 1455 => to_unsigned(1815, 12), 1456 => to_unsigned(2257, 12), 1457 => to_unsigned(1999, 12), 1458 => to_unsigned(1822, 12), 1459 => to_unsigned(2127, 12), 1460 => to_unsigned(2018, 12), 1461 => to_unsigned(2421, 12), 1462 => to_unsigned(2016, 12), 1463 => to_unsigned(1509, 12), 1464 => to_unsigned(2335, 12), 1465 => to_unsigned(2775, 12), 1466 => to_unsigned(2121, 12), 1467 => to_unsigned(2545, 12), 1468 => to_unsigned(1991, 12), 1469 => to_unsigned(1526, 12), 1470 => to_unsigned(1311, 12), 1471 => to_unsigned(1922, 12), 1472 => to_unsigned(1416, 12), 1473 => to_unsigned(2523, 12), 1474 => to_unsigned(2401, 12), 1475 => to_unsigned(2374, 12), 1476 => to_unsigned(2015, 12), 1477 => to_unsigned(1955, 12), 1478 => to_unsigned(2025, 12), 1479 => to_unsigned(2084, 12), 1480 => to_unsigned(1867, 12), 1481 => to_unsigned(2091, 12), 1482 => to_unsigned(1812, 12), 1483 => to_unsigned(2147, 12), 1484 => to_unsigned(2750, 12), 1485 => to_unsigned(2704, 12), 1486 => to_unsigned(1920, 12), 1487 => to_unsigned(1617, 12), 1488 => to_unsigned(2165, 12), 1489 => to_unsigned(2545, 12), 1490 => to_unsigned(1808, 12), 1491 => to_unsigned(2365, 12), 1492 => to_unsigned(2454, 12), 1493 => to_unsigned(1985, 12), 1494 => to_unsigned(1381, 12), 1495 => to_unsigned(1755, 12), 1496 => to_unsigned(2062, 12), 1497 => to_unsigned(2155, 12), 1498 => to_unsigned(1434, 12), 1499 => to_unsigned(2328, 12), 1500 => to_unsigned(1943, 12), 1501 => to_unsigned(2447, 12), 1502 => to_unsigned(1474, 12), 1503 => to_unsigned(1780, 12), 1504 => to_unsigned(1919, 12), 1505 => to_unsigned(2041, 12), 1506 => to_unsigned(2854, 12), 1507 => to_unsigned(1807, 12), 1508 => to_unsigned(2136, 12), 1509 => to_unsigned(2151, 12), 1510 => to_unsigned(2204, 12), 1511 => to_unsigned(2565, 12), 1512 => to_unsigned(1841, 12), 1513 => to_unsigned(1491, 12), 1514 => to_unsigned(1339, 12), 1515 => to_unsigned(2123, 12), 1516 => to_unsigned(1956, 12), 1517 => to_unsigned(2381, 12), 1518 => to_unsigned(2436, 12), 1519 => to_unsigned(1877, 12), 1520 => to_unsigned(1925, 12), 1521 => to_unsigned(1898, 12), 1522 => to_unsigned(2095, 12), 1523 => to_unsigned(2286, 12), 1524 => to_unsigned(1847, 12), 1525 => to_unsigned(2318, 12), 1526 => to_unsigned(2180, 12), 1527 => to_unsigned(1962, 12), 1528 => to_unsigned(2304, 12), 1529 => to_unsigned(1807, 12), 1530 => to_unsigned(2243, 12), 1531 => to_unsigned(2180, 12), 1532 => to_unsigned(2499, 12), 1533 => to_unsigned(2099, 12), 1534 => to_unsigned(2376, 12), 1535 => to_unsigned(1998, 12), 1536 => to_unsigned(1737, 12), 1537 => to_unsigned(2753, 12), 1538 => to_unsigned(1734, 12), 1539 => to_unsigned(1577, 12), 1540 => to_unsigned(1590, 12), 1541 => to_unsigned(2238, 12), 1542 => to_unsigned(2015, 12), 1543 => to_unsigned(2800, 12), 1544 => to_unsigned(2194, 12), 1545 => to_unsigned(2159, 12), 1546 => to_unsigned(2333, 12), 1547 => to_unsigned(2178, 12), 1548 => to_unsigned(1766, 12), 1549 => to_unsigned(1647, 12), 1550 => to_unsigned(2496, 12), 1551 => to_unsigned(2411, 12), 1552 => to_unsigned(2182, 12), 1553 => to_unsigned(2155, 12), 1554 => to_unsigned(1586, 12), 1555 => to_unsigned(1557, 12), 1556 => to_unsigned(2215, 12), 1557 => to_unsigned(2607, 12), 1558 => to_unsigned(1567, 12), 1559 => to_unsigned(1856, 12), 1560 => to_unsigned(2734, 12), 1561 => to_unsigned(2182, 12), 1562 => to_unsigned(1941, 12), 1563 => to_unsigned(2299, 12), 1564 => to_unsigned(1997, 12), 1565 => to_unsigned(1915, 12), 1566 => to_unsigned(3264, 12), 1567 => to_unsigned(1870, 12), 1568 => to_unsigned(1648, 12), 1569 => to_unsigned(2814, 12), 1570 => to_unsigned(1436, 12), 1571 => to_unsigned(2157, 12), 1572 => to_unsigned(1175, 12), 1573 => to_unsigned(2087, 12), 1574 => to_unsigned(2396, 12), 1575 => to_unsigned(1775, 12), 1576 => to_unsigned(2542, 12), 1577 => to_unsigned(2984, 12), 1578 => to_unsigned(2079, 12), 1579 => to_unsigned(2150, 12), 1580 => to_unsigned(1416, 12), 1581 => to_unsigned(1305, 12), 1582 => to_unsigned(973, 12), 1583 => to_unsigned(1817, 12), 1584 => to_unsigned(2149, 12), 1585 => to_unsigned(2507, 12), 1586 => to_unsigned(2157, 12), 1587 => to_unsigned(2131, 12), 1588 => to_unsigned(2130, 12), 1589 => to_unsigned(1803, 12), 1590 => to_unsigned(2592, 12), 1591 => to_unsigned(1754, 12), 1592 => to_unsigned(1832, 12), 1593 => to_unsigned(2614, 12), 1594 => to_unsigned(1858, 12), 1595 => to_unsigned(2610, 12), 1596 => to_unsigned(2002, 12), 1597 => to_unsigned(1921, 12), 1598 => to_unsigned(1913, 12), 1599 => to_unsigned(1936, 12), 1600 => to_unsigned(1838, 12), 1601 => to_unsigned(2242, 12), 1602 => to_unsigned(2295, 12), 1603 => to_unsigned(3180, 12), 1604 => to_unsigned(1842, 12), 1605 => to_unsigned(1608, 12), 1606 => to_unsigned(2358, 12), 1607 => to_unsigned(2213, 12), 1608 => to_unsigned(2415, 12), 1609 => to_unsigned(1412, 12), 1610 => to_unsigned(2359, 12), 1611 => to_unsigned(1917, 12), 1612 => to_unsigned(1904, 12), 1613 => to_unsigned(2507, 12), 1614 => to_unsigned(2219, 12), 1615 => to_unsigned(2126, 12), 1616 => to_unsigned(2103, 12), 1617 => to_unsigned(1519, 12), 1618 => to_unsigned(2404, 12), 1619 => to_unsigned(2042, 12), 1620 => to_unsigned(1505, 12), 1621 => to_unsigned(1835, 12), 1622 => to_unsigned(1855, 12), 1623 => to_unsigned(1316, 12), 1624 => to_unsigned(2339, 12), 1625 => to_unsigned(2239, 12), 1626 => to_unsigned(2154, 12), 1627 => to_unsigned(2007, 12), 1628 => to_unsigned(1440, 12), 1629 => to_unsigned(2153, 12), 1630 => to_unsigned(1436, 12), 1631 => to_unsigned(2025, 12), 1632 => to_unsigned(1879, 12), 1633 => to_unsigned(2236, 12), 1634 => to_unsigned(2390, 12), 1635 => to_unsigned(2051, 12), 1636 => to_unsigned(1613, 12), 1637 => to_unsigned(2105, 12), 1638 => to_unsigned(2442, 12), 1639 => to_unsigned(1810, 12), 1640 => to_unsigned(1829, 12), 1641 => to_unsigned(2057, 12), 1642 => to_unsigned(1876, 12), 1643 => to_unsigned(2398, 12), 1644 => to_unsigned(1820, 12), 1645 => to_unsigned(1760, 12), 1646 => to_unsigned(2271, 12), 1647 => to_unsigned(2148, 12), 1648 => to_unsigned(2409, 12), 1649 => to_unsigned(1707, 12), 1650 => to_unsigned(1500, 12), 1651 => to_unsigned(1826, 12), 1652 => to_unsigned(1958, 12), 1653 => to_unsigned(2581, 12), 1654 => to_unsigned(2142, 12), 1655 => to_unsigned(2370, 12), 1656 => to_unsigned(1906, 12), 1657 => to_unsigned(1175, 12), 1658 => to_unsigned(1963, 12), 1659 => to_unsigned(2546, 12), 1660 => to_unsigned(1772, 12), 1661 => to_unsigned(1598, 12), 1662 => to_unsigned(2230, 12), 1663 => to_unsigned(1820, 12), 1664 => to_unsigned(1751, 12), 1665 => to_unsigned(1825, 12), 1666 => to_unsigned(1657, 12), 1667 => to_unsigned(2197, 12), 1668 => to_unsigned(2001, 12), 1669 => to_unsigned(2045, 12), 1670 => to_unsigned(2060, 12), 1671 => to_unsigned(2840, 12), 1672 => to_unsigned(2109, 12), 1673 => to_unsigned(1879, 12), 1674 => to_unsigned(1958, 12), 1675 => to_unsigned(1916, 12), 1676 => to_unsigned(1244, 12), 1677 => to_unsigned(2429, 12), 1678 => to_unsigned(2045, 12), 1679 => to_unsigned(2393, 12), 1680 => to_unsigned(1725, 12), 1681 => to_unsigned(2222, 12), 1682 => to_unsigned(1895, 12), 1683 => to_unsigned(2084, 12), 1684 => to_unsigned(1791, 12), 1685 => to_unsigned(1475, 12), 1686 => to_unsigned(2166, 12), 1687 => to_unsigned(2209, 12), 1688 => to_unsigned(2132, 12), 1689 => to_unsigned(1442, 12), 1690 => to_unsigned(2498, 12), 1691 => to_unsigned(1364, 12), 1692 => to_unsigned(2121, 12), 1693 => to_unsigned(1840, 12), 1694 => to_unsigned(2360, 12), 1695 => to_unsigned(1743, 12), 1696 => to_unsigned(1847, 12), 1697 => to_unsigned(1921, 12), 1698 => to_unsigned(1740, 12), 1699 => to_unsigned(2644, 12), 1700 => to_unsigned(1577, 12), 1701 => to_unsigned(2026, 12), 1702 => to_unsigned(2377, 12), 1703 => to_unsigned(1963, 12), 1704 => to_unsigned(2165, 12), 1705 => to_unsigned(2825, 12), 1706 => to_unsigned(2869, 12), 1707 => to_unsigned(1951, 12), 1708 => to_unsigned(1141, 12), 1709 => to_unsigned(1657, 12), 1710 => to_unsigned(2286, 12), 1711 => to_unsigned(1452, 12), 1712 => to_unsigned(2111, 12), 1713 => to_unsigned(2086, 12), 1714 => to_unsigned(2401, 12), 1715 => to_unsigned(2149, 12), 1716 => to_unsigned(2181, 12), 1717 => to_unsigned(1905, 12), 1718 => to_unsigned(1418, 12), 1719 => to_unsigned(1745, 12), 1720 => to_unsigned(2024, 12), 1721 => to_unsigned(2408, 12), 1722 => to_unsigned(2159, 12), 1723 => to_unsigned(2325, 12), 1724 => to_unsigned(2417, 12), 1725 => to_unsigned(2099, 12), 1726 => to_unsigned(2089, 12), 1727 => to_unsigned(2119, 12), 1728 => to_unsigned(2083, 12), 1729 => to_unsigned(2296, 12), 1730 => to_unsigned(1734, 12), 1731 => to_unsigned(1089, 12), 1732 => to_unsigned(1509, 12), 1733 => to_unsigned(1800, 12), 1734 => to_unsigned(1488, 12), 1735 => to_unsigned(1425, 12), 1736 => to_unsigned(2296, 12), 1737 => to_unsigned(1368, 12), 1738 => to_unsigned(1554, 12), 1739 => to_unsigned(2044, 12), 1740 => to_unsigned(2127, 12), 1741 => to_unsigned(2314, 12), 1742 => to_unsigned(2207, 12), 1743 => to_unsigned(2577, 12), 1744 => to_unsigned(1517, 12), 1745 => to_unsigned(2210, 12), 1746 => to_unsigned(1770, 12), 1747 => to_unsigned(1763, 12), 1748 => to_unsigned(2265, 12), 1749 => to_unsigned(2026, 12), 1750 => to_unsigned(2232, 12), 1751 => to_unsigned(2537, 12), 1752 => to_unsigned(1915, 12), 1753 => to_unsigned(1906, 12), 1754 => to_unsigned(1921, 12), 1755 => to_unsigned(2294, 12), 1756 => to_unsigned(2186, 12), 1757 => to_unsigned(1973, 12), 1758 => to_unsigned(2049, 12), 1759 => to_unsigned(2851, 12), 1760 => to_unsigned(2089, 12), 1761 => to_unsigned(2598, 12), 1762 => to_unsigned(2073, 12), 1763 => to_unsigned(1479, 12), 1764 => to_unsigned(2240, 12), 1765 => to_unsigned(1925, 12), 1766 => to_unsigned(1562, 12), 1767 => to_unsigned(1845, 12), 1768 => to_unsigned(1919, 12), 1769 => to_unsigned(1800, 12), 1770 => to_unsigned(2215, 12), 1771 => to_unsigned(2310, 12), 1772 => to_unsigned(2096, 12), 1773 => to_unsigned(2274, 12), 1774 => to_unsigned(2327, 12), 1775 => to_unsigned(2150, 12), 1776 => to_unsigned(1820, 12), 1777 => to_unsigned(2417, 12), 1778 => to_unsigned(2329, 12), 1779 => to_unsigned(2009, 12), 1780 => to_unsigned(2559, 12), 1781 => to_unsigned(2349, 12), 1782 => to_unsigned(1935, 12), 1783 => to_unsigned(3115, 12), 1784 => to_unsigned(2310, 12), 1785 => to_unsigned(2255, 12), 1786 => to_unsigned(2140, 12), 1787 => to_unsigned(2266, 12), 1788 => to_unsigned(2198, 12), 1789 => to_unsigned(1683, 12), 1790 => to_unsigned(2185, 12), 1791 => to_unsigned(2048, 12), 1792 => to_unsigned(1856, 12), 1793 => to_unsigned(2068, 12), 1794 => to_unsigned(2501, 12), 1795 => to_unsigned(1487, 12), 1796 => to_unsigned(1847, 12), 1797 => to_unsigned(2572, 12), 1798 => to_unsigned(2337, 12), 1799 => to_unsigned(1864, 12), 1800 => to_unsigned(2476, 12), 1801 => to_unsigned(2099, 12), 1802 => to_unsigned(2360, 12), 1803 => to_unsigned(1870, 12), 1804 => to_unsigned(1519, 12), 1805 => to_unsigned(1988, 12), 1806 => to_unsigned(2135, 12), 1807 => to_unsigned(1420, 12), 1808 => to_unsigned(1724, 12), 1809 => to_unsigned(2184, 12), 1810 => to_unsigned(1919, 12), 1811 => to_unsigned(1851, 12), 1812 => to_unsigned(2264, 12), 1813 => to_unsigned(1367, 12), 1814 => to_unsigned(1793, 12), 1815 => to_unsigned(1732, 12), 1816 => to_unsigned(2152, 12), 1817 => to_unsigned(2128, 12), 1818 => to_unsigned(1628, 12), 1819 => to_unsigned(2467, 12), 1820 => to_unsigned(3105, 12), 1821 => to_unsigned(1755, 12), 1822 => to_unsigned(1425, 12), 1823 => to_unsigned(2119, 12), 1824 => to_unsigned(2598, 12), 1825 => to_unsigned(1565, 12), 1826 => to_unsigned(1511, 12), 1827 => to_unsigned(2361, 12), 1828 => to_unsigned(2203, 12), 1829 => to_unsigned(1883, 12), 1830 => to_unsigned(1892, 12), 1831 => to_unsigned(2446, 12), 1832 => to_unsigned(2288, 12), 1833 => to_unsigned(1751, 12), 1834 => to_unsigned(2066, 12), 1835 => to_unsigned(1913, 12), 1836 => to_unsigned(1730, 12), 1837 => to_unsigned(1863, 12), 1838 => to_unsigned(1787, 12), 1839 => to_unsigned(2337, 12), 1840 => to_unsigned(2558, 12), 1841 => to_unsigned(1800, 12), 1842 => to_unsigned(1838, 12), 1843 => to_unsigned(2147, 12), 1844 => to_unsigned(2003, 12), 1845 => to_unsigned(1688, 12), 1846 => to_unsigned(2245, 12), 1847 => to_unsigned(2113, 12), 1848 => to_unsigned(2141, 12), 1849 => to_unsigned(2427, 12), 1850 => to_unsigned(2569, 12), 1851 => to_unsigned(2520, 12), 1852 => to_unsigned(2308, 12), 1853 => to_unsigned(1575, 12), 1854 => to_unsigned(1931, 12), 1855 => to_unsigned(1968, 12), 1856 => to_unsigned(1959, 12), 1857 => to_unsigned(1980, 12), 1858 => to_unsigned(1532, 12), 1859 => to_unsigned(2071, 12), 1860 => to_unsigned(2304, 12), 1861 => to_unsigned(2127, 12), 1862 => to_unsigned(1909, 12), 1863 => to_unsigned(2084, 12), 1864 => to_unsigned(2915, 12), 1865 => to_unsigned(2036, 12), 1866 => to_unsigned(2391, 12), 1867 => to_unsigned(2534, 12), 1868 => to_unsigned(1643, 12), 1869 => to_unsigned(1514, 12), 1870 => to_unsigned(1720, 12), 1871 => to_unsigned(2064, 12), 1872 => to_unsigned(2479, 12), 1873 => to_unsigned(2063, 12), 1874 => to_unsigned(2277, 12), 1875 => to_unsigned(2070, 12), 1876 => to_unsigned(2281, 12), 1877 => to_unsigned(1935, 12), 1878 => to_unsigned(1747, 12), 1879 => to_unsigned(1881, 12), 1880 => to_unsigned(1921, 12), 1881 => to_unsigned(2299, 12), 1882 => to_unsigned(1700, 12), 1883 => to_unsigned(2089, 12), 1884 => to_unsigned(1881, 12), 1885 => to_unsigned(2068, 12), 1886 => to_unsigned(1963, 12), 1887 => to_unsigned(1769, 12), 1888 => to_unsigned(1987, 12), 1889 => to_unsigned(1666, 12), 1890 => to_unsigned(2615, 12), 1891 => to_unsigned(2010, 12), 1892 => to_unsigned(2588, 12), 1893 => to_unsigned(2095, 12), 1894 => to_unsigned(1341, 12), 1895 => to_unsigned(1810, 12), 1896 => to_unsigned(2007, 12), 1897 => to_unsigned(2148, 12), 1898 => to_unsigned(2126, 12), 1899 => to_unsigned(1680, 12), 1900 => to_unsigned(1485, 12), 1901 => to_unsigned(2012, 12), 1902 => to_unsigned(1769, 12), 1903 => to_unsigned(1941, 12), 1904 => to_unsigned(1717, 12), 1905 => to_unsigned(2137, 12), 1906 => to_unsigned(2414, 12), 1907 => to_unsigned(1528, 12), 1908 => to_unsigned(1606, 12), 1909 => to_unsigned(1990, 12), 1910 => to_unsigned(2048, 12), 1911 => to_unsigned(1848, 12), 1912 => to_unsigned(1735, 12), 1913 => to_unsigned(2283, 12), 1914 => to_unsigned(1986, 12), 1915 => to_unsigned(2066, 12), 1916 => to_unsigned(1827, 12), 1917 => to_unsigned(2533, 12), 1918 => to_unsigned(1309, 12), 1919 => to_unsigned(3415, 12), 1920 => to_unsigned(1954, 12), 1921 => to_unsigned(1723, 12), 1922 => to_unsigned(1663, 12), 1923 => to_unsigned(1860, 12), 1924 => to_unsigned(2056, 12), 1925 => to_unsigned(1634, 12), 1926 => to_unsigned(2083, 12), 1927 => to_unsigned(2094, 12), 1928 => to_unsigned(2216, 12), 1929 => to_unsigned(2289, 12), 1930 => to_unsigned(1748, 12), 1931 => to_unsigned(2313, 12), 1932 => to_unsigned(1836, 12), 1933 => to_unsigned(2145, 12), 1934 => to_unsigned(2306, 12), 1935 => to_unsigned(2290, 12), 1936 => to_unsigned(2191, 12), 1937 => to_unsigned(2101, 12), 1938 => to_unsigned(2104, 12), 1939 => to_unsigned(2196, 12), 1940 => to_unsigned(2060, 12), 1941 => to_unsigned(1918, 12), 1942 => to_unsigned(1750, 12), 1943 => to_unsigned(2256, 12), 1944 => to_unsigned(2208, 12), 1945 => to_unsigned(1780, 12), 1946 => to_unsigned(2107, 12), 1947 => to_unsigned(2126, 12), 1948 => to_unsigned(2269, 12), 1949 => to_unsigned(1652, 12), 1950 => to_unsigned(2182, 12), 1951 => to_unsigned(1741, 12), 1952 => to_unsigned(2031, 12), 1953 => to_unsigned(1560, 12), 1954 => to_unsigned(2336, 12), 1955 => to_unsigned(1591, 12), 1956 => to_unsigned(2031, 12), 1957 => to_unsigned(2488, 12), 1958 => to_unsigned(1360, 12), 1959 => to_unsigned(2332, 12), 1960 => to_unsigned(1920, 12), 1961 => to_unsigned(1737, 12), 1962 => to_unsigned(2360, 12), 1963 => to_unsigned(1868, 12), 1964 => to_unsigned(1666, 12), 1965 => to_unsigned(2122, 12), 1966 => to_unsigned(2105, 12), 1967 => to_unsigned(1391, 12), 1968 => to_unsigned(2069, 12), 1969 => to_unsigned(2211, 12), 1970 => to_unsigned(1804, 12), 1971 => to_unsigned(2699, 12), 1972 => to_unsigned(1637, 12), 1973 => to_unsigned(2377, 12), 1974 => to_unsigned(2269, 12), 1975 => to_unsigned(1928, 12), 1976 => to_unsigned(1779, 12), 1977 => to_unsigned(1997, 12), 1978 => to_unsigned(2564, 12), 1979 => to_unsigned(1615, 12), 1980 => to_unsigned(2122, 12), 1981 => to_unsigned(1764, 12), 1982 => to_unsigned(1993, 12), 1983 => to_unsigned(2008, 12), 1984 => to_unsigned(2624, 12), 1985 => to_unsigned(2298, 12), 1986 => to_unsigned(1886, 12), 1987 => to_unsigned(1873, 12), 1988 => to_unsigned(2191, 12), 1989 => to_unsigned(1878, 12), 1990 => to_unsigned(1972, 12), 1991 => to_unsigned(2748, 12), 1992 => to_unsigned(2164, 12), 1993 => to_unsigned(3053, 12), 1994 => to_unsigned(2171, 12), 1995 => to_unsigned(2196, 12), 1996 => to_unsigned(2204, 12), 1997 => to_unsigned(1806, 12), 1998 => to_unsigned(2007, 12), 1999 => to_unsigned(2209, 12), 2000 => to_unsigned(2251, 12), 2001 => to_unsigned(2168, 12), 2002 => to_unsigned(1326, 12), 2003 => to_unsigned(1226, 12), 2004 => to_unsigned(2044, 12), 2005 => to_unsigned(1756, 12), 2006 => to_unsigned(2265, 12), 2007 => to_unsigned(2249, 12), 2008 => to_unsigned(2115, 12), 2009 => to_unsigned(2218, 12), 2010 => to_unsigned(1822, 12), 2011 => to_unsigned(1890, 12), 2012 => to_unsigned(2175, 12), 2013 => to_unsigned(1199, 12), 2014 => to_unsigned(1630, 12), 2015 => to_unsigned(1903, 12), 2016 => to_unsigned(2876, 12), 2017 => to_unsigned(2398, 12), 2018 => to_unsigned(1991, 12), 2019 => to_unsigned(1831, 12), 2020 => to_unsigned(2055, 12), 2021 => to_unsigned(2242, 12), 2022 => to_unsigned(1664, 12), 2023 => to_unsigned(1772, 12), 2024 => to_unsigned(1298, 12), 2025 => to_unsigned(1920, 12), 2026 => to_unsigned(2227, 12), 2027 => to_unsigned(1601, 12), 2028 => to_unsigned(1907, 12), 2029 => to_unsigned(2543, 12), 2030 => to_unsigned(1820, 12), 2031 => to_unsigned(2127, 12), 2032 => to_unsigned(2668, 12), 2033 => to_unsigned(1659, 12), 2034 => to_unsigned(2177, 12), 2035 => to_unsigned(2498, 12), 2036 => to_unsigned(1649, 12), 2037 => to_unsigned(2537, 12), 2038 => to_unsigned(1872, 12), 2039 => to_unsigned(2151, 12), 2040 => to_unsigned(2057, 12), 2041 => to_unsigned(1950, 12), 2042 => to_unsigned(2523, 12), 2043 => to_unsigned(1651, 12), 2044 => to_unsigned(1298, 12), 2045 => to_unsigned(2691, 12), 2046 => to_unsigned(2041, 12), 2047 => to_unsigned(1864, 12))
    );

    pure function slice_data(data : data_t; color : integer; row : integer; pixel : integer) return vnir_pixel_t is
        variable data_color : vnir_row_window_t;
        variable data_color_row : vnir_row_t;
    begin
        data_color := data(color);
        data_color_row := data_color(row);
        return data_color_row(pixel);
    end;

begin

	-- Generate main clock signal
	clock_gen : process
	begin
		wait for clock_period / 2;
		clock <= not clock;
	end process clock_gen;
    

    test : process
        constant window_size : integer := 10;
        constant fragment_size : integer := 512;
	begin

        report "Uploading started";
        for color in 0 to 2 loop
            for row in 0 to window_size-1 loop
                for fragment in 0 to fragment_size-1 loop
                    pixels_available <= '1';
                    pixels(0) <= slice_data(data, color, row, fragment);
                    pixels(1) <= slice_data(data, color, row, fragment + fragment_size);
                    pixels(2) <= slice_data(data, color, row, fragment + fragment_size * 2);
                    pixels(3) <= slice_data(data, color, row, fragment + fragment_size * 3);
                    wait until rising_edge(clock);
                end loop;
            end loop;
        end loop;
        report "Uploading finished";

        pixels_available <= '0';
        wait until rising_edge(clock);
        assert rows_available = '1' report "********************* Rows not available";
        assert row_red = averages(0) report "********************* Red row incorrect";
        assert row_blue = averages(1) report "********************* Blue row incorrect";
        assert row_nir = averages(2) report "********************* NIR row incorrect";

        report "Finished running tests.";

        wait;
    end process test;

    collate_rows_component : collate_rows port map (
        clock => clock,
        reset_n => reset_n,
        pixels => pixels,
        pixels_available => pixels_available,
        row_red => row_red,
        row_blue => row_blue,
        row_nir => row_nir,
        rows_available => rows_available
    );

end tests;
