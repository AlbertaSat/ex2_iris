----------------------------------------------------------------
-- Copyright 2020 University of Alberta

-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at

--     http://www.apache.org/licenses/LICENSE-2.0

-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
----------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.spi_types.all;
use work.vnir_types.all;
use work.test_util.all;

entity row_collator_tb is
end entity row_collator_tb;

architecture tests of row_collator_tb is
	signal clock            : std_logic := '0';
	signal reset_n          : std_logic := '1';
    signal config           : vnir_config_t;
    signal read_config      : std_logic := '0';
    signal pixels           : vnir_pixel_vector_t(vnir_lvds_data_width-1 downto 0);
	signal pixels_available	: std_logic := '0';
	signal rows             : vnir_rows_t;
	signal rows_available   : std_logic := '0';

    component row_collator is
    port (
        clock            : in std_logic;
        reset_n          : in std_logic;
        config           : in vnir_config_t;
        read_config      : in std_logic;
        pixels           : in vnir_pixel_vector_t(vnir_lvds_data_width-1 downto 0);
        pixels_available : in std_logic;
        rows             : out vnir_rows_t;
        rows_available   : out std_logic
    );
    end component row_collator;

    constant n_colours : integer := 3;
    constant window_size : integer := 10;  -- Matches row_collator_tb_datagen.py
    type vnir_row_window_t is array(window_size-1 downto 0) of vnir_row_t;
    type data_t is array(n_colours-1 downto 0) of vnir_row_window_t;
    type averages_t is array(n_colours-1 downto 0) of vnir_row_t;
    
    constant data : data_t := (
        0 => (
            0 => (0 => to_unsigned(684, 10), 1 => to_unsigned(559, 10), 2 => to_unsigned(629, 10), 3 => to_unsigned(192, 10), 4 => to_unsigned(835, 10), 5 => to_unsigned(763, 10), 6 => to_unsigned(707, 10), 7 => to_unsigned(359, 10), 8 => to_unsigned(9, 10), 9 => to_unsigned(723, 10), 10 => to_unsigned(277, 10), 11 => to_unsigned(754, 10), 12 => to_unsigned(804, 10), 13 => to_unsigned(599, 10), 14 => to_unsigned(70, 10), 15 => to_unsigned(472, 10), 16 => to_unsigned(600, 10), 17 => to_unsigned(396, 10), 18 => to_unsigned(314, 10), 19 => to_unsigned(705, 10), 20 => to_unsigned(486, 10), 21 => to_unsigned(551, 10), 22 => to_unsigned(87, 10), 23 => to_unsigned(174, 10), 24 => to_unsigned(600, 10), 25 => to_unsigned(849, 10), 26 => to_unsigned(677, 10), 27 => to_unsigned(537, 10), 28 => to_unsigned(845, 10), 29 => to_unsigned(72, 10), 30 => to_unsigned(777, 10), 31 => to_unsigned(916, 10), 32 => to_unsigned(115, 10), 33 => to_unsigned(976, 10), 34 => to_unsigned(755, 10), 35 => to_unsigned(709, 10), 36 => to_unsigned(1022, 10), 37 => to_unsigned(847, 10), 38 => to_unsigned(431, 10), 39 => to_unsigned(448, 10), 40 => to_unsigned(850, 10), 41 => to_unsigned(99, 10), 42 => to_unsigned(984, 10), 43 => to_unsigned(177, 10), 44 => to_unsigned(755, 10), 45 => to_unsigned(797, 10), 46 => to_unsigned(659, 10), 47 => to_unsigned(147, 10), 48 => to_unsigned(910, 10), 49 => to_unsigned(423, 10), 50 => to_unsigned(288, 10), 51 => to_unsigned(961, 10), 52 => to_unsigned(265, 10), 53 => to_unsigned(697, 10), 54 => to_unsigned(639, 10), 55 => to_unsigned(544, 10), 56 => to_unsigned(543, 10), 57 => to_unsigned(714, 10), 58 => to_unsigned(244, 10), 59 => to_unsigned(151, 10), 60 => to_unsigned(675, 10), 61 => to_unsigned(510, 10), 62 => to_unsigned(459, 10), 63 => to_unsigned(882, 10), 64 => to_unsigned(183, 10), 65 => to_unsigned(28, 10), 66 => to_unsigned(802, 10), 67 => to_unsigned(128, 10), 68 => to_unsigned(128, 10), 69 => to_unsigned(932, 10), 70 => to_unsigned(53, 10), 71 => to_unsigned(901, 10), 72 => to_unsigned(550, 10), 73 => to_unsigned(488, 10), 74 => to_unsigned(756, 10), 75 => to_unsigned(273, 10), 76 => to_unsigned(335, 10), 77 => to_unsigned(388, 10), 78 => to_unsigned(617, 10), 79 => to_unsigned(42, 10), 80 => to_unsigned(442, 10), 81 => to_unsigned(543, 10), 82 => to_unsigned(888, 10), 83 => to_unsigned(257, 10), 84 => to_unsigned(321, 10), 85 => to_unsigned(999, 10), 86 => to_unsigned(937, 10), 87 => to_unsigned(57, 10), 88 => to_unsigned(291, 10), 89 => to_unsigned(870, 10), 90 => to_unsigned(119, 10), 91 => to_unsigned(779, 10), 92 => to_unsigned(430, 10), 93 => to_unsigned(82, 10), 94 => to_unsigned(91, 10), 95 => to_unsigned(896, 10), 96 => to_unsigned(398, 10), 97 => to_unsigned(611, 10), 98 => to_unsigned(565, 10), 99 => to_unsigned(908, 10), 100 => to_unsigned(633, 10), 101 => to_unsigned(938, 10), 102 => to_unsigned(84, 10), 103 => to_unsigned(203, 10), 104 => to_unsigned(324, 10), 105 => to_unsigned(774, 10), 106 => to_unsigned(964, 10), 107 => to_unsigned(47, 10), 108 => to_unsigned(639, 10), 109 => to_unsigned(1012, 10), 110 => to_unsigned(131, 10), 111 => to_unsigned(972, 10), 112 => to_unsigned(868, 10), 113 => to_unsigned(180, 10), 114 => to_unsigned(1000, 10), 115 => to_unsigned(846, 10), 116 => to_unsigned(143, 10), 117 => to_unsigned(660, 10), 118 => to_unsigned(227, 10), 119 => to_unsigned(954, 10), 120 => to_unsigned(791, 10), 121 => to_unsigned(719, 10), 122 => to_unsigned(909, 10), 123 => to_unsigned(373, 10), 124 => to_unsigned(853, 10), 125 => to_unsigned(560, 10), 126 => to_unsigned(305, 10), 127 => to_unsigned(581, 10), 128 => to_unsigned(169, 10), 129 => to_unsigned(675, 10), 130 => to_unsigned(448, 10), 131 => to_unsigned(95, 10), 132 => to_unsigned(197, 10), 133 => to_unsigned(606, 10), 134 => to_unsigned(256, 10), 135 => to_unsigned(881, 10), 136 => to_unsigned(690, 10), 137 => to_unsigned(292, 10), 138 => to_unsigned(930, 10), 139 => to_unsigned(816, 10), 140 => to_unsigned(861, 10), 141 => to_unsigned(387, 10), 142 => to_unsigned(610, 10), 143 => to_unsigned(554, 10), 144 => to_unsigned(973, 10), 145 => to_unsigned(368, 10), 146 => to_unsigned(999, 10), 147 => to_unsigned(917, 10), 148 => to_unsigned(201, 10), 149 => to_unsigned(383, 10), 150 => to_unsigned(512, 10), 151 => to_unsigned(906, 10), 152 => to_unsigned(370, 10), 153 => to_unsigned(555, 10), 154 => to_unsigned(954, 10), 155 => to_unsigned(383, 10), 156 => to_unsigned(23, 10), 157 => to_unsigned(699, 10), 158 => to_unsigned(130, 10), 159 => to_unsigned(377, 10), 160 => to_unsigned(98, 10), 161 => to_unsigned(574, 10), 162 => to_unsigned(931, 10), 163 => to_unsigned(734, 10), 164 => to_unsigned(123, 10), 165 => to_unsigned(963, 10), 166 => to_unsigned(594, 10), 167 => to_unsigned(942, 10), 168 => to_unsigned(739, 10), 169 => to_unsigned(148, 10), 170 => to_unsigned(209, 10), 171 => to_unsigned(562, 10), 172 => to_unsigned(411, 10), 173 => to_unsigned(782, 10), 174 => to_unsigned(41, 10), 175 => to_unsigned(58, 10), 176 => to_unsigned(705, 10), 177 => to_unsigned(36, 10), 178 => to_unsigned(778, 10), 179 => to_unsigned(86, 10), 180 => to_unsigned(43, 10), 181 => to_unsigned(872, 10), 182 => to_unsigned(11, 10), 183 => to_unsigned(770, 10), 184 => to_unsigned(307, 10), 185 => to_unsigned(80, 10), 186 => to_unsigned(32, 10), 187 => to_unsigned(182, 10), 188 => to_unsigned(128, 10), 189 => to_unsigned(806, 10), 190 => to_unsigned(275, 10), 191 => to_unsigned(174, 10), 192 => to_unsigned(554, 10), 193 => to_unsigned(371, 10), 194 => to_unsigned(184, 10), 195 => to_unsigned(444, 10), 196 => to_unsigned(488, 10), 197 => to_unsigned(589, 10), 198 => to_unsigned(286, 10), 199 => to_unsigned(280, 10), 200 => to_unsigned(637, 10), 201 => to_unsigned(770, 10), 202 => to_unsigned(515, 10), 203 => to_unsigned(94, 10), 204 => to_unsigned(226, 10), 205 => to_unsigned(875, 10), 206 => to_unsigned(269, 10), 207 => to_unsigned(880, 10), 208 => to_unsigned(296, 10), 209 => to_unsigned(328, 10), 210 => to_unsigned(19, 10), 211 => to_unsigned(607, 10), 212 => to_unsigned(840, 10), 213 => to_unsigned(410, 10), 214 => to_unsigned(450, 10), 215 => to_unsigned(248, 10), 216 => to_unsigned(180, 10), 217 => to_unsigned(323, 10), 218 => to_unsigned(1004, 10), 219 => to_unsigned(829, 10), 220 => to_unsigned(782, 10), 221 => to_unsigned(864, 10), 222 => to_unsigned(260, 10), 223 => to_unsigned(963, 10), 224 => to_unsigned(749, 10), 225 => to_unsigned(139, 10), 226 => to_unsigned(1020, 10), 227 => to_unsigned(598, 10), 228 => to_unsigned(461, 10), 229 => to_unsigned(889, 10), 230 => to_unsigned(621, 10), 231 => to_unsigned(843, 10), 232 => to_unsigned(696, 10), 233 => to_unsigned(528, 10), 234 => to_unsigned(152, 10), 235 => to_unsigned(925, 10), 236 => to_unsigned(149, 10), 237 => to_unsigned(110, 10), 238 => to_unsigned(25, 10), 239 => to_unsigned(464, 10), 240 => to_unsigned(956, 10), 241 => to_unsigned(889, 10), 242 => to_unsigned(886, 10), 243 => to_unsigned(117, 10), 244 => to_unsigned(445, 10), 245 => to_unsigned(595, 10), 246 => to_unsigned(673, 10), 247 => to_unsigned(872, 10), 248 => to_unsigned(928, 10), 249 => to_unsigned(228, 10), 250 => to_unsigned(507, 10), 251 => to_unsigned(763, 10), 252 => to_unsigned(121, 10), 253 => to_unsigned(326, 10), 254 => to_unsigned(469, 10), 255 => to_unsigned(287, 10), 256 => to_unsigned(525, 10), 257 => to_unsigned(839, 10), 258 => to_unsigned(696, 10), 259 => to_unsigned(152, 10), 260 => to_unsigned(591, 10), 261 => to_unsigned(41, 10), 262 => to_unsigned(274, 10), 263 => to_unsigned(552, 10), 264 => to_unsigned(438, 10), 265 => to_unsigned(207, 10), 266 => to_unsigned(779, 10), 267 => to_unsigned(166, 10), 268 => to_unsigned(111, 10), 269 => to_unsigned(349, 10), 270 => to_unsigned(1017, 10), 271 => to_unsigned(129, 10), 272 => to_unsigned(735, 10), 273 => to_unsigned(886, 10), 274 => to_unsigned(812, 10), 275 => to_unsigned(216, 10), 276 => to_unsigned(381, 10), 277 => to_unsigned(24, 10), 278 => to_unsigned(67, 10), 279 => to_unsigned(978, 10), 280 => to_unsigned(1007, 10), 281 => to_unsigned(771, 10), 282 => to_unsigned(234, 10), 283 => to_unsigned(716, 10), 284 => to_unsigned(998, 10), 285 => to_unsigned(291, 10), 286 => to_unsigned(726, 10), 287 => to_unsigned(1022, 10), 288 => to_unsigned(701, 10), 289 => to_unsigned(709, 10), 290 => to_unsigned(727, 10), 291 => to_unsigned(555, 10), 292 => to_unsigned(32, 10), 293 => to_unsigned(11, 10), 294 => to_unsigned(616, 10), 295 => to_unsigned(212, 10), 296 => to_unsigned(138, 10), 297 => to_unsigned(694, 10), 298 => to_unsigned(1003, 10), 299 => to_unsigned(421, 10), 300 => to_unsigned(637, 10), 301 => to_unsigned(668, 10), 302 => to_unsigned(623, 10), 303 => to_unsigned(488, 10), 304 => to_unsigned(770, 10), 305 => to_unsigned(539, 10), 306 => to_unsigned(979, 10), 307 => to_unsigned(217, 10), 308 => to_unsigned(663, 10), 309 => to_unsigned(821, 10), 310 => to_unsigned(307, 10), 311 => to_unsigned(174, 10), 312 => to_unsigned(148, 10), 313 => to_unsigned(949, 10), 314 => to_unsigned(541, 10), 315 => to_unsigned(579, 10), 316 => to_unsigned(547, 10), 317 => to_unsigned(807, 10), 318 => to_unsigned(393, 10), 319 => to_unsigned(73, 10), 320 => to_unsigned(297, 10), 321 => to_unsigned(919, 10), 322 => to_unsigned(899, 10), 323 => to_unsigned(814, 10), 324 => to_unsigned(730, 10), 325 => to_unsigned(946, 10), 326 => to_unsigned(876, 10), 327 => to_unsigned(771, 10), 328 => to_unsigned(799, 10), 329 => to_unsigned(777, 10), 330 => to_unsigned(394, 10), 331 => to_unsigned(539, 10), 332 => to_unsigned(429, 10), 333 => to_unsigned(199, 10), 334 => to_unsigned(423, 10), 335 => to_unsigned(61, 10), 336 => to_unsigned(341, 10), 337 => to_unsigned(865, 10), 338 => to_unsigned(44, 10), 339 => to_unsigned(802, 10), 340 => to_unsigned(930, 10), 341 => to_unsigned(88, 10), 342 => to_unsigned(33, 10), 343 => to_unsigned(645, 10), 344 => to_unsigned(232, 10), 345 => to_unsigned(767, 10), 346 => to_unsigned(36, 10), 347 => to_unsigned(768, 10), 348 => to_unsigned(459, 10), 349 => to_unsigned(290, 10), 350 => to_unsigned(197, 10), 351 => to_unsigned(894, 10), 352 => to_unsigned(949, 10), 353 => to_unsigned(254, 10), 354 => to_unsigned(80, 10), 355 => to_unsigned(446, 10), 356 => to_unsigned(136, 10), 357 => to_unsigned(189, 10), 358 => to_unsigned(129, 10), 359 => to_unsigned(209, 10), 360 => to_unsigned(368, 10), 361 => to_unsigned(291, 10), 362 => to_unsigned(376, 10), 363 => to_unsigned(347, 10), 364 => to_unsigned(168, 10), 365 => to_unsigned(884, 10), 366 => to_unsigned(804, 10), 367 => to_unsigned(176, 10), 368 => to_unsigned(537, 10), 369 => to_unsigned(323, 10), 370 => to_unsigned(871, 10), 371 => to_unsigned(508, 10), 372 => to_unsigned(803, 10), 373 => to_unsigned(114, 10), 374 => to_unsigned(798, 10), 375 => to_unsigned(29, 10), 376 => to_unsigned(753, 10), 377 => to_unsigned(289, 10), 378 => to_unsigned(146, 10), 379 => to_unsigned(273, 10), 380 => to_unsigned(221, 10), 381 => to_unsigned(340, 10), 382 => to_unsigned(509, 10), 383 => to_unsigned(514, 10), 384 => to_unsigned(69, 10), 385 => to_unsigned(357, 10), 386 => to_unsigned(908, 10), 387 => to_unsigned(556, 10), 388 => to_unsigned(885, 10), 389 => to_unsigned(765, 10), 390 => to_unsigned(322, 10), 391 => to_unsigned(623, 10), 392 => to_unsigned(91, 10), 393 => to_unsigned(341, 10), 394 => to_unsigned(423, 10), 395 => to_unsigned(551, 10), 396 => to_unsigned(971, 10), 397 => to_unsigned(662, 10), 398 => to_unsigned(414, 10), 399 => to_unsigned(657, 10), 400 => to_unsigned(710, 10), 401 => to_unsigned(967, 10), 402 => to_unsigned(274, 10), 403 => to_unsigned(860, 10), 404 => to_unsigned(43, 10), 405 => to_unsigned(83, 10), 406 => to_unsigned(433, 10), 407 => to_unsigned(809, 10), 408 => to_unsigned(93, 10), 409 => to_unsigned(174, 10), 410 => to_unsigned(405, 10), 411 => to_unsigned(201, 10), 412 => to_unsigned(857, 10), 413 => to_unsigned(498, 10), 414 => to_unsigned(480, 10), 415 => to_unsigned(987, 10), 416 => to_unsigned(329, 10), 417 => to_unsigned(540, 10), 418 => to_unsigned(1003, 10), 419 => to_unsigned(209, 10), 420 => to_unsigned(617, 10), 421 => to_unsigned(954, 10), 422 => to_unsigned(896, 10), 423 => to_unsigned(982, 10), 424 => to_unsigned(575, 10), 425 => to_unsigned(16, 10), 426 => to_unsigned(106, 10), 427 => to_unsigned(164, 10), 428 => to_unsigned(606, 10), 429 => to_unsigned(536, 10), 430 => to_unsigned(628, 10), 431 => to_unsigned(191, 10), 432 => to_unsigned(195, 10), 433 => to_unsigned(307, 10), 434 => to_unsigned(136, 10), 435 => to_unsigned(952, 10), 436 => to_unsigned(859, 10), 437 => to_unsigned(93, 10), 438 => to_unsigned(891, 10), 439 => to_unsigned(750, 10), 440 => to_unsigned(87, 10), 441 => to_unsigned(160, 10), 442 => to_unsigned(147, 10), 443 => to_unsigned(584, 10), 444 => to_unsigned(455, 10), 445 => to_unsigned(87, 10), 446 => to_unsigned(13, 10), 447 => to_unsigned(314, 10), 448 => to_unsigned(593, 10), 449 => to_unsigned(120, 10), 450 => to_unsigned(884, 10), 451 => to_unsigned(951, 10), 452 => to_unsigned(832, 10), 453 => to_unsigned(715, 10), 454 => to_unsigned(732, 10), 455 => to_unsigned(932, 10), 456 => to_unsigned(281, 10), 457 => to_unsigned(800, 10), 458 => to_unsigned(426, 10), 459 => to_unsigned(782, 10), 460 => to_unsigned(470, 10), 461 => to_unsigned(284, 10), 462 => to_unsigned(276, 10), 463 => to_unsigned(978, 10), 464 => to_unsigned(324, 10), 465 => to_unsigned(534, 10), 466 => to_unsigned(227, 10), 467 => to_unsigned(890, 10), 468 => to_unsigned(595, 10), 469 => to_unsigned(647, 10), 470 => to_unsigned(968, 10), 471 => to_unsigned(573, 10), 472 => to_unsigned(653, 10), 473 => to_unsigned(517, 10), 474 => to_unsigned(256, 10), 475 => to_unsigned(136, 10), 476 => to_unsigned(207, 10), 477 => to_unsigned(463, 10), 478 => to_unsigned(949, 10), 479 => to_unsigned(139, 10), 480 => to_unsigned(4, 10), 481 => to_unsigned(423, 10), 482 => to_unsigned(348, 10), 483 => to_unsigned(941, 10), 484 => to_unsigned(282, 10), 485 => to_unsigned(586, 10), 486 => to_unsigned(820, 10), 487 => to_unsigned(1006, 10), 488 => to_unsigned(433, 10), 489 => to_unsigned(219, 10), 490 => to_unsigned(819, 10), 491 => to_unsigned(739, 10), 492 => to_unsigned(873, 10), 493 => to_unsigned(786, 10), 494 => to_unsigned(373, 10), 495 => to_unsigned(290, 10), 496 => to_unsigned(563, 10), 497 => to_unsigned(670, 10), 498 => to_unsigned(437, 10), 499 => to_unsigned(826, 10), 500 => to_unsigned(939, 10), 501 => to_unsigned(823, 10), 502 => to_unsigned(508, 10), 503 => to_unsigned(1020, 10), 504 => to_unsigned(786, 10), 505 => to_unsigned(941, 10), 506 => to_unsigned(855, 10), 507 => to_unsigned(449, 10), 508 => to_unsigned(326, 10), 509 => to_unsigned(490, 10), 510 => to_unsigned(53, 10), 511 => to_unsigned(816, 10), 512 => to_unsigned(94, 10), 513 => to_unsigned(59, 10), 514 => to_unsigned(336, 10), 515 => to_unsigned(666, 10), 516 => to_unsigned(636, 10), 517 => to_unsigned(163, 10), 518 => to_unsigned(570, 10), 519 => to_unsigned(945, 10), 520 => to_unsigned(106, 10), 521 => to_unsigned(201, 10), 522 => to_unsigned(300, 10), 523 => to_unsigned(781, 10), 524 => to_unsigned(889, 10), 525 => to_unsigned(838, 10), 526 => to_unsigned(550, 10), 527 => to_unsigned(679, 10), 528 => to_unsigned(648, 10), 529 => to_unsigned(13, 10), 530 => to_unsigned(1016, 10), 531 => to_unsigned(903, 10), 532 => to_unsigned(720, 10), 533 => to_unsigned(1016, 10), 534 => to_unsigned(534, 10), 535 => to_unsigned(504, 10), 536 => to_unsigned(847, 10), 537 => to_unsigned(985, 10), 538 => to_unsigned(776, 10), 539 => to_unsigned(739, 10), 540 => to_unsigned(774, 10), 541 => to_unsigned(209, 10), 542 => to_unsigned(455, 10), 543 => to_unsigned(468, 10), 544 => to_unsigned(473, 10), 545 => to_unsigned(962, 10), 546 => to_unsigned(572, 10), 547 => to_unsigned(400, 10), 548 => to_unsigned(56, 10), 549 => to_unsigned(882, 10), 550 => to_unsigned(749, 10), 551 => to_unsigned(663, 10), 552 => to_unsigned(280, 10), 553 => to_unsigned(4, 10), 554 => to_unsigned(612, 10), 555 => to_unsigned(1004, 10), 556 => to_unsigned(305, 10), 557 => to_unsigned(343, 10), 558 => to_unsigned(542, 10), 559 => to_unsigned(566, 10), 560 => to_unsigned(153, 10), 561 => to_unsigned(788, 10), 562 => to_unsigned(353, 10), 563 => to_unsigned(357, 10), 564 => to_unsigned(697, 10), 565 => to_unsigned(407, 10), 566 => to_unsigned(411, 10), 567 => to_unsigned(29, 10), 568 => to_unsigned(929, 10), 569 => to_unsigned(371, 10), 570 => to_unsigned(821, 10), 571 => to_unsigned(631, 10), 572 => to_unsigned(947, 10), 573 => to_unsigned(854, 10), 574 => to_unsigned(502, 10), 575 => to_unsigned(7, 10), 576 => to_unsigned(617, 10), 577 => to_unsigned(1009, 10), 578 => to_unsigned(137, 10), 579 => to_unsigned(694, 10), 580 => to_unsigned(896, 10), 581 => to_unsigned(851, 10), 582 => to_unsigned(376, 10), 583 => to_unsigned(932, 10), 584 => to_unsigned(721, 10), 585 => to_unsigned(148, 10), 586 => to_unsigned(885, 10), 587 => to_unsigned(1008, 10), 588 => to_unsigned(259, 10), 589 => to_unsigned(126, 10), 590 => to_unsigned(810, 10), 591 => to_unsigned(577, 10), 592 => to_unsigned(532, 10), 593 => to_unsigned(804, 10), 594 => to_unsigned(324, 10), 595 => to_unsigned(976, 10), 596 => to_unsigned(112, 10), 597 => to_unsigned(943, 10), 598 => to_unsigned(650, 10), 599 => to_unsigned(237, 10), 600 => to_unsigned(360, 10), 601 => to_unsigned(990, 10), 602 => to_unsigned(859, 10), 603 => to_unsigned(555, 10), 604 => to_unsigned(63, 10), 605 => to_unsigned(927, 10), 606 => to_unsigned(916, 10), 607 => to_unsigned(454, 10), 608 => to_unsigned(265, 10), 609 => to_unsigned(444, 10), 610 => to_unsigned(603, 10), 611 => to_unsigned(623, 10), 612 => to_unsigned(419, 10), 613 => to_unsigned(339, 10), 614 => to_unsigned(844, 10), 615 => to_unsigned(274, 10), 616 => to_unsigned(369, 10), 617 => to_unsigned(842, 10), 618 => to_unsigned(226, 10), 619 => to_unsigned(225, 10), 620 => to_unsigned(939, 10), 621 => to_unsigned(643, 10), 622 => to_unsigned(908, 10), 623 => to_unsigned(228, 10), 624 => to_unsigned(826, 10), 625 => to_unsigned(897, 10), 626 => to_unsigned(369, 10), 627 => to_unsigned(128, 10), 628 => to_unsigned(807, 10), 629 => to_unsigned(24, 10), 630 => to_unsigned(698, 10), 631 => to_unsigned(292, 10), 632 => to_unsigned(355, 10), 633 => to_unsigned(837, 10), 634 => to_unsigned(134, 10), 635 => to_unsigned(3, 10), 636 => to_unsigned(226, 10), 637 => to_unsigned(889, 10), 638 => to_unsigned(680, 10), 639 => to_unsigned(444, 10), 640 => to_unsigned(417, 10), 641 => to_unsigned(284, 10), 642 => to_unsigned(836, 10), 643 => to_unsigned(26, 10), 644 => to_unsigned(736, 10), 645 => to_unsigned(248, 10), 646 => to_unsigned(365, 10), 647 => to_unsigned(947, 10), 648 => to_unsigned(201, 10), 649 => to_unsigned(437, 10), 650 => to_unsigned(197, 10), 651 => to_unsigned(929, 10), 652 => to_unsigned(647, 10), 653 => to_unsigned(637, 10), 654 => to_unsigned(606, 10), 655 => to_unsigned(72, 10), 656 => to_unsigned(246, 10), 657 => to_unsigned(852, 10), 658 => to_unsigned(135, 10), 659 => to_unsigned(707, 10), 660 => to_unsigned(213, 10), 661 => to_unsigned(475, 10), 662 => to_unsigned(620, 10), 663 => to_unsigned(323, 10), 664 => to_unsigned(102, 10), 665 => to_unsigned(852, 10), 666 => to_unsigned(327, 10), 667 => to_unsigned(595, 10), 668 => to_unsigned(223, 10), 669 => to_unsigned(256, 10), 670 => to_unsigned(645, 10), 671 => to_unsigned(347, 10), 672 => to_unsigned(107, 10), 673 => to_unsigned(926, 10), 674 => to_unsigned(969, 10), 675 => to_unsigned(979, 10), 676 => to_unsigned(519, 10), 677 => to_unsigned(149, 10), 678 => to_unsigned(997, 10), 679 => to_unsigned(476, 10), 680 => to_unsigned(392, 10), 681 => to_unsigned(683, 10), 682 => to_unsigned(558, 10), 683 => to_unsigned(0, 10), 684 => to_unsigned(360, 10), 685 => to_unsigned(691, 10), 686 => to_unsigned(550, 10), 687 => to_unsigned(89, 10), 688 => to_unsigned(74, 10), 689 => to_unsigned(499, 10), 690 => to_unsigned(738, 10), 691 => to_unsigned(635, 10), 692 => to_unsigned(343, 10), 693 => to_unsigned(96, 10), 694 => to_unsigned(851, 10), 695 => to_unsigned(282, 10), 696 => to_unsigned(718, 10), 697 => to_unsigned(32, 10), 698 => to_unsigned(115, 10), 699 => to_unsigned(454, 10), 700 => to_unsigned(865, 10), 701 => to_unsigned(428, 10), 702 => to_unsigned(827, 10), 703 => to_unsigned(825, 10), 704 => to_unsigned(690, 10), 705 => to_unsigned(173, 10), 706 => to_unsigned(745, 10), 707 => to_unsigned(132, 10), 708 => to_unsigned(441, 10), 709 => to_unsigned(93, 10), 710 => to_unsigned(347, 10), 711 => to_unsigned(401, 10), 712 => to_unsigned(419, 10), 713 => to_unsigned(706, 10), 714 => to_unsigned(404, 10), 715 => to_unsigned(941, 10), 716 => to_unsigned(185, 10), 717 => to_unsigned(975, 10), 718 => to_unsigned(375, 10), 719 => to_unsigned(676, 10), 720 => to_unsigned(873, 10), 721 => to_unsigned(702, 10), 722 => to_unsigned(516, 10), 723 => to_unsigned(497, 10), 724 => to_unsigned(498, 10), 725 => to_unsigned(205, 10), 726 => to_unsigned(414, 10), 727 => to_unsigned(365, 10), 728 => to_unsigned(855, 10), 729 => to_unsigned(738, 10), 730 => to_unsigned(419, 10), 731 => to_unsigned(585, 10), 732 => to_unsigned(218, 10), 733 => to_unsigned(951, 10), 734 => to_unsigned(538, 10), 735 => to_unsigned(374, 10), 736 => to_unsigned(22, 10), 737 => to_unsigned(460, 10), 738 => to_unsigned(719, 10), 739 => to_unsigned(354, 10), 740 => to_unsigned(602, 10), 741 => to_unsigned(51, 10), 742 => to_unsigned(998, 10), 743 => to_unsigned(814, 10), 744 => to_unsigned(720, 10), 745 => to_unsigned(573, 10), 746 => to_unsigned(444, 10), 747 => to_unsigned(815, 10), 748 => to_unsigned(1018, 10), 749 => to_unsigned(104, 10), 750 => to_unsigned(640, 10), 751 => to_unsigned(394, 10), 752 => to_unsigned(971, 10), 753 => to_unsigned(909, 10), 754 => to_unsigned(327, 10), 755 => to_unsigned(606, 10), 756 => to_unsigned(518, 10), 757 => to_unsigned(685, 10), 758 => to_unsigned(245, 10), 759 => to_unsigned(414, 10), 760 => to_unsigned(527, 10), 761 => to_unsigned(169, 10), 762 => to_unsigned(166, 10), 763 => to_unsigned(309, 10), 764 => to_unsigned(939, 10), 765 => to_unsigned(594, 10), 766 => to_unsigned(391, 10), 767 => to_unsigned(220, 10), 768 => to_unsigned(833, 10), 769 => to_unsigned(681, 10), 770 => to_unsigned(834, 10), 771 => to_unsigned(114, 10), 772 => to_unsigned(860, 10), 773 => to_unsigned(334, 10), 774 => to_unsigned(741, 10), 775 => to_unsigned(219, 10), 776 => to_unsigned(246, 10), 777 => to_unsigned(100, 10), 778 => to_unsigned(415, 10), 779 => to_unsigned(221, 10), 780 => to_unsigned(178, 10), 781 => to_unsigned(508, 10), 782 => to_unsigned(174, 10), 783 => to_unsigned(605, 10), 784 => to_unsigned(626, 10), 785 => to_unsigned(673, 10), 786 => to_unsigned(780, 10), 787 => to_unsigned(736, 10), 788 => to_unsigned(745, 10), 789 => to_unsigned(848, 10), 790 => to_unsigned(66, 10), 791 => to_unsigned(456, 10), 792 => to_unsigned(1011, 10), 793 => to_unsigned(125, 10), 794 => to_unsigned(138, 10), 795 => to_unsigned(624, 10), 796 => to_unsigned(730, 10), 797 => to_unsigned(155, 10), 798 => to_unsigned(696, 10), 799 => to_unsigned(120, 10), 800 => to_unsigned(321, 10), 801 => to_unsigned(448, 10), 802 => to_unsigned(709, 10), 803 => to_unsigned(856, 10), 804 => to_unsigned(290, 10), 805 => to_unsigned(975, 10), 806 => to_unsigned(3, 10), 807 => to_unsigned(700, 10), 808 => to_unsigned(238, 10), 809 => to_unsigned(677, 10), 810 => to_unsigned(171, 10), 811 => to_unsigned(723, 10), 812 => to_unsigned(856, 10), 813 => to_unsigned(582, 10), 814 => to_unsigned(660, 10), 815 => to_unsigned(902, 10), 816 => to_unsigned(796, 10), 817 => to_unsigned(627, 10), 818 => to_unsigned(902, 10), 819 => to_unsigned(834, 10), 820 => to_unsigned(604, 10), 821 => to_unsigned(988, 10), 822 => to_unsigned(614, 10), 823 => to_unsigned(869, 10), 824 => to_unsigned(379, 10), 825 => to_unsigned(709, 10), 826 => to_unsigned(109, 10), 827 => to_unsigned(329, 10), 828 => to_unsigned(100, 10), 829 => to_unsigned(694, 10), 830 => to_unsigned(845, 10), 831 => to_unsigned(917, 10), 832 => to_unsigned(507, 10), 833 => to_unsigned(671, 10), 834 => to_unsigned(593, 10), 835 => to_unsigned(35, 10), 836 => to_unsigned(237, 10), 837 => to_unsigned(243, 10), 838 => to_unsigned(250, 10), 839 => to_unsigned(392, 10), 840 => to_unsigned(766, 10), 841 => to_unsigned(281, 10), 842 => to_unsigned(21, 10), 843 => to_unsigned(429, 10), 844 => to_unsigned(229, 10), 845 => to_unsigned(982, 10), 846 => to_unsigned(400, 10), 847 => to_unsigned(153, 10), 848 => to_unsigned(1006, 10), 849 => to_unsigned(119, 10), 850 => to_unsigned(677, 10), 851 => to_unsigned(895, 10), 852 => to_unsigned(385, 10), 853 => to_unsigned(389, 10), 854 => to_unsigned(710, 10), 855 => to_unsigned(396, 10), 856 => to_unsigned(346, 10), 857 => to_unsigned(586, 10), 858 => to_unsigned(1019, 10), 859 => to_unsigned(950, 10), 860 => to_unsigned(78, 10), 861 => to_unsigned(830, 10), 862 => to_unsigned(584, 10), 863 => to_unsigned(199, 10), 864 => to_unsigned(813, 10), 865 => to_unsigned(133, 10), 866 => to_unsigned(559, 10), 867 => to_unsigned(699, 10), 868 => to_unsigned(170, 10), 869 => to_unsigned(451, 10), 870 => to_unsigned(138, 10), 871 => to_unsigned(754, 10), 872 => to_unsigned(313, 10), 873 => to_unsigned(475, 10), 874 => to_unsigned(345, 10), 875 => to_unsigned(387, 10), 876 => to_unsigned(125, 10), 877 => to_unsigned(718, 10), 878 => to_unsigned(850, 10), 879 => to_unsigned(197, 10), 880 => to_unsigned(698, 10), 881 => to_unsigned(900, 10), 882 => to_unsigned(17, 10), 883 => to_unsigned(709, 10), 884 => to_unsigned(447, 10), 885 => to_unsigned(350, 10), 886 => to_unsigned(664, 10), 887 => to_unsigned(643, 10), 888 => to_unsigned(325, 10), 889 => to_unsigned(424, 10), 890 => to_unsigned(164, 10), 891 => to_unsigned(570, 10), 892 => to_unsigned(177, 10), 893 => to_unsigned(439, 10), 894 => to_unsigned(664, 10), 895 => to_unsigned(673, 10), 896 => to_unsigned(914, 10), 897 => to_unsigned(865, 10), 898 => to_unsigned(462, 10), 899 => to_unsigned(753, 10), 900 => to_unsigned(135, 10), 901 => to_unsigned(949, 10), 902 => to_unsigned(747, 10), 903 => to_unsigned(46, 10), 904 => to_unsigned(496, 10), 905 => to_unsigned(1012, 10), 906 => to_unsigned(639, 10), 907 => to_unsigned(929, 10), 908 => to_unsigned(337, 10), 909 => to_unsigned(157, 10), 910 => to_unsigned(524, 10), 911 => to_unsigned(630, 10), 912 => to_unsigned(814, 10), 913 => to_unsigned(886, 10), 914 => to_unsigned(288, 10), 915 => to_unsigned(802, 10), 916 => to_unsigned(115, 10), 917 => to_unsigned(599, 10), 918 => to_unsigned(636, 10), 919 => to_unsigned(409, 10), 920 => to_unsigned(174, 10), 921 => to_unsigned(498, 10), 922 => to_unsigned(875, 10), 923 => to_unsigned(564, 10), 924 => to_unsigned(1001, 10), 925 => to_unsigned(622, 10), 926 => to_unsigned(576, 10), 927 => to_unsigned(332, 10), 928 => to_unsigned(886, 10), 929 => to_unsigned(585, 10), 930 => to_unsigned(146, 10), 931 => to_unsigned(772, 10), 932 => to_unsigned(775, 10), 933 => to_unsigned(643, 10), 934 => to_unsigned(48, 10), 935 => to_unsigned(76, 10), 936 => to_unsigned(293, 10), 937 => to_unsigned(116, 10), 938 => to_unsigned(493, 10), 939 => to_unsigned(560, 10), 940 => to_unsigned(109, 10), 941 => to_unsigned(978, 10), 942 => to_unsigned(179, 10), 943 => to_unsigned(561, 10), 944 => to_unsigned(71, 10), 945 => to_unsigned(858, 10), 946 => to_unsigned(433, 10), 947 => to_unsigned(1006, 10), 948 => to_unsigned(285, 10), 949 => to_unsigned(515, 10), 950 => to_unsigned(74, 10), 951 => to_unsigned(596, 10), 952 => to_unsigned(490, 10), 953 => to_unsigned(321, 10), 954 => to_unsigned(887, 10), 955 => to_unsigned(532, 10), 956 => to_unsigned(208, 10), 957 => to_unsigned(42, 10), 958 => to_unsigned(498, 10), 959 => to_unsigned(28, 10), 960 => to_unsigned(410, 10), 961 => to_unsigned(855, 10), 962 => to_unsigned(180, 10), 963 => to_unsigned(304, 10), 964 => to_unsigned(962, 10), 965 => to_unsigned(614, 10), 966 => to_unsigned(777, 10), 967 => to_unsigned(258, 10), 968 => to_unsigned(372, 10), 969 => to_unsigned(876, 10), 970 => to_unsigned(745, 10), 971 => to_unsigned(857, 10), 972 => to_unsigned(380, 10), 973 => to_unsigned(885, 10), 974 => to_unsigned(612, 10), 975 => to_unsigned(90, 10), 976 => to_unsigned(68, 10), 977 => to_unsigned(617, 10), 978 => to_unsigned(522, 10), 979 => to_unsigned(12, 10), 980 => to_unsigned(616, 10), 981 => to_unsigned(225, 10), 982 => to_unsigned(421, 10), 983 => to_unsigned(167, 10), 984 => to_unsigned(928, 10), 985 => to_unsigned(378, 10), 986 => to_unsigned(289, 10), 987 => to_unsigned(922, 10), 988 => to_unsigned(99, 10), 989 => to_unsigned(217, 10), 990 => to_unsigned(306, 10), 991 => to_unsigned(344, 10), 992 => to_unsigned(210, 10), 993 => to_unsigned(788, 10), 994 => to_unsigned(734, 10), 995 => to_unsigned(668, 10), 996 => to_unsigned(584, 10), 997 => to_unsigned(274, 10), 998 => to_unsigned(409, 10), 999 => to_unsigned(920, 10), 1000 => to_unsigned(551, 10), 1001 => to_unsigned(234, 10), 1002 => to_unsigned(635, 10), 1003 => to_unsigned(284, 10), 1004 => to_unsigned(664, 10), 1005 => to_unsigned(658, 10), 1006 => to_unsigned(707, 10), 1007 => to_unsigned(172, 10), 1008 => to_unsigned(723, 10), 1009 => to_unsigned(301, 10), 1010 => to_unsigned(822, 10), 1011 => to_unsigned(0, 10), 1012 => to_unsigned(138, 10), 1013 => to_unsigned(707, 10), 1014 => to_unsigned(902, 10), 1015 => to_unsigned(731, 10), 1016 => to_unsigned(867, 10), 1017 => to_unsigned(441, 10), 1018 => to_unsigned(966, 10), 1019 => to_unsigned(915, 10), 1020 => to_unsigned(162, 10), 1021 => to_unsigned(50, 10), 1022 => to_unsigned(242, 10), 1023 => to_unsigned(870, 10), 1024 => to_unsigned(20, 10), 1025 => to_unsigned(683, 10), 1026 => to_unsigned(630, 10), 1027 => to_unsigned(128, 10), 1028 => to_unsigned(484, 10), 1029 => to_unsigned(365, 10), 1030 => to_unsigned(105, 10), 1031 => to_unsigned(706, 10), 1032 => to_unsigned(225, 10), 1033 => to_unsigned(652, 10), 1034 => to_unsigned(783, 10), 1035 => to_unsigned(118, 10), 1036 => to_unsigned(545, 10), 1037 => to_unsigned(151, 10), 1038 => to_unsigned(908, 10), 1039 => to_unsigned(901, 10), 1040 => to_unsigned(38, 10), 1041 => to_unsigned(769, 10), 1042 => to_unsigned(266, 10), 1043 => to_unsigned(6, 10), 1044 => to_unsigned(893, 10), 1045 => to_unsigned(262, 10), 1046 => to_unsigned(614, 10), 1047 => to_unsigned(934, 10), 1048 => to_unsigned(331, 10), 1049 => to_unsigned(370, 10), 1050 => to_unsigned(341, 10), 1051 => to_unsigned(382, 10), 1052 => to_unsigned(370, 10), 1053 => to_unsigned(690, 10), 1054 => to_unsigned(819, 10), 1055 => to_unsigned(258, 10), 1056 => to_unsigned(332, 10), 1057 => to_unsigned(669, 10), 1058 => to_unsigned(521, 10), 1059 => to_unsigned(627, 10), 1060 => to_unsigned(968, 10), 1061 => to_unsigned(389, 10), 1062 => to_unsigned(628, 10), 1063 => to_unsigned(181, 10), 1064 => to_unsigned(235, 10), 1065 => to_unsigned(193, 10), 1066 => to_unsigned(811, 10), 1067 => to_unsigned(591, 10), 1068 => to_unsigned(62, 10), 1069 => to_unsigned(332, 10), 1070 => to_unsigned(559, 10), 1071 => to_unsigned(588, 10), 1072 => to_unsigned(661, 10), 1073 => to_unsigned(120, 10), 1074 => to_unsigned(786, 10), 1075 => to_unsigned(345, 10), 1076 => to_unsigned(525, 10), 1077 => to_unsigned(222, 10), 1078 => to_unsigned(604, 10), 1079 => to_unsigned(236, 10), 1080 => to_unsigned(105, 10), 1081 => to_unsigned(213, 10), 1082 => to_unsigned(518, 10), 1083 => to_unsigned(612, 10), 1084 => to_unsigned(560, 10), 1085 => to_unsigned(552, 10), 1086 => to_unsigned(922, 10), 1087 => to_unsigned(158, 10), 1088 => to_unsigned(389, 10), 1089 => to_unsigned(143, 10), 1090 => to_unsigned(959, 10), 1091 => to_unsigned(485, 10), 1092 => to_unsigned(37, 10), 1093 => to_unsigned(571, 10), 1094 => to_unsigned(625, 10), 1095 => to_unsigned(95, 10), 1096 => to_unsigned(352, 10), 1097 => to_unsigned(496, 10), 1098 => to_unsigned(208, 10), 1099 => to_unsigned(288, 10), 1100 => to_unsigned(62, 10), 1101 => to_unsigned(394, 10), 1102 => to_unsigned(396, 10), 1103 => to_unsigned(605, 10), 1104 => to_unsigned(832, 10), 1105 => to_unsigned(413, 10), 1106 => to_unsigned(346, 10), 1107 => to_unsigned(999, 10), 1108 => to_unsigned(150, 10), 1109 => to_unsigned(403, 10), 1110 => to_unsigned(389, 10), 1111 => to_unsigned(804, 10), 1112 => to_unsigned(595, 10), 1113 => to_unsigned(127, 10), 1114 => to_unsigned(484, 10), 1115 => to_unsigned(773, 10), 1116 => to_unsigned(348, 10), 1117 => to_unsigned(460, 10), 1118 => to_unsigned(154, 10), 1119 => to_unsigned(753, 10), 1120 => to_unsigned(83, 10), 1121 => to_unsigned(908, 10), 1122 => to_unsigned(998, 10), 1123 => to_unsigned(135, 10), 1124 => to_unsigned(180, 10), 1125 => to_unsigned(592, 10), 1126 => to_unsigned(413, 10), 1127 => to_unsigned(0, 10), 1128 => to_unsigned(727, 10), 1129 => to_unsigned(719, 10), 1130 => to_unsigned(842, 10), 1131 => to_unsigned(764, 10), 1132 => to_unsigned(643, 10), 1133 => to_unsigned(573, 10), 1134 => to_unsigned(323, 10), 1135 => to_unsigned(144, 10), 1136 => to_unsigned(880, 10), 1137 => to_unsigned(457, 10), 1138 => to_unsigned(596, 10), 1139 => to_unsigned(116, 10), 1140 => to_unsigned(741, 10), 1141 => to_unsigned(767, 10), 1142 => to_unsigned(824, 10), 1143 => to_unsigned(318, 10), 1144 => to_unsigned(952, 10), 1145 => to_unsigned(560, 10), 1146 => to_unsigned(145, 10), 1147 => to_unsigned(885, 10), 1148 => to_unsigned(953, 10), 1149 => to_unsigned(521, 10), 1150 => to_unsigned(492, 10), 1151 => to_unsigned(190, 10), 1152 => to_unsigned(79, 10), 1153 => to_unsigned(742, 10), 1154 => to_unsigned(206, 10), 1155 => to_unsigned(417, 10), 1156 => to_unsigned(900, 10), 1157 => to_unsigned(912, 10), 1158 => to_unsigned(228, 10), 1159 => to_unsigned(839, 10), 1160 => to_unsigned(318, 10), 1161 => to_unsigned(791, 10), 1162 => to_unsigned(859, 10), 1163 => to_unsigned(366, 10), 1164 => to_unsigned(7, 10), 1165 => to_unsigned(509, 10), 1166 => to_unsigned(790, 10), 1167 => to_unsigned(866, 10), 1168 => to_unsigned(158, 10), 1169 => to_unsigned(758, 10), 1170 => to_unsigned(592, 10), 1171 => to_unsigned(155, 10), 1172 => to_unsigned(559, 10), 1173 => to_unsigned(495, 10), 1174 => to_unsigned(626, 10), 1175 => to_unsigned(523, 10), 1176 => to_unsigned(983, 10), 1177 => to_unsigned(846, 10), 1178 => to_unsigned(999, 10), 1179 => to_unsigned(798, 10), 1180 => to_unsigned(90, 10), 1181 => to_unsigned(290, 10), 1182 => to_unsigned(566, 10), 1183 => to_unsigned(849, 10), 1184 => to_unsigned(675, 10), 1185 => to_unsigned(71, 10), 1186 => to_unsigned(877, 10), 1187 => to_unsigned(827, 10), 1188 => to_unsigned(624, 10), 1189 => to_unsigned(421, 10), 1190 => to_unsigned(68, 10), 1191 => to_unsigned(437, 10), 1192 => to_unsigned(13, 10), 1193 => to_unsigned(101, 10), 1194 => to_unsigned(787, 10), 1195 => to_unsigned(875, 10), 1196 => to_unsigned(264, 10), 1197 => to_unsigned(864, 10), 1198 => to_unsigned(721, 10), 1199 => to_unsigned(197, 10), 1200 => to_unsigned(380, 10), 1201 => to_unsigned(100, 10), 1202 => to_unsigned(385, 10), 1203 => to_unsigned(765, 10), 1204 => to_unsigned(157, 10), 1205 => to_unsigned(901, 10), 1206 => to_unsigned(976, 10), 1207 => to_unsigned(230, 10), 1208 => to_unsigned(504, 10), 1209 => to_unsigned(936, 10), 1210 => to_unsigned(662, 10), 1211 => to_unsigned(30, 10), 1212 => to_unsigned(255, 10), 1213 => to_unsigned(531, 10), 1214 => to_unsigned(772, 10), 1215 => to_unsigned(660, 10), 1216 => to_unsigned(874, 10), 1217 => to_unsigned(586, 10), 1218 => to_unsigned(123, 10), 1219 => to_unsigned(451, 10), 1220 => to_unsigned(214, 10), 1221 => to_unsigned(316, 10), 1222 => to_unsigned(741, 10), 1223 => to_unsigned(250, 10), 1224 => to_unsigned(605, 10), 1225 => to_unsigned(681, 10), 1226 => to_unsigned(552, 10), 1227 => to_unsigned(188, 10), 1228 => to_unsigned(209, 10), 1229 => to_unsigned(691, 10), 1230 => to_unsigned(296, 10), 1231 => to_unsigned(59, 10), 1232 => to_unsigned(490, 10), 1233 => to_unsigned(478, 10), 1234 => to_unsigned(541, 10), 1235 => to_unsigned(225, 10), 1236 => to_unsigned(606, 10), 1237 => to_unsigned(238, 10), 1238 => to_unsigned(677, 10), 1239 => to_unsigned(382, 10), 1240 => to_unsigned(216, 10), 1241 => to_unsigned(272, 10), 1242 => to_unsigned(867, 10), 1243 => to_unsigned(167, 10), 1244 => to_unsigned(669, 10), 1245 => to_unsigned(508, 10), 1246 => to_unsigned(65, 10), 1247 => to_unsigned(791, 10), 1248 => to_unsigned(200, 10), 1249 => to_unsigned(384, 10), 1250 => to_unsigned(87, 10), 1251 => to_unsigned(805, 10), 1252 => to_unsigned(367, 10), 1253 => to_unsigned(447, 10), 1254 => to_unsigned(410, 10), 1255 => to_unsigned(729, 10), 1256 => to_unsigned(345, 10), 1257 => to_unsigned(134, 10), 1258 => to_unsigned(216, 10), 1259 => to_unsigned(503, 10), 1260 => to_unsigned(463, 10), 1261 => to_unsigned(101, 10), 1262 => to_unsigned(297, 10), 1263 => to_unsigned(913, 10), 1264 => to_unsigned(976, 10), 1265 => to_unsigned(880, 10), 1266 => to_unsigned(43, 10), 1267 => to_unsigned(110, 10), 1268 => to_unsigned(453, 10), 1269 => to_unsigned(374, 10), 1270 => to_unsigned(915, 10), 1271 => to_unsigned(751, 10), 1272 => to_unsigned(790, 10), 1273 => to_unsigned(365, 10), 1274 => to_unsigned(907, 10), 1275 => to_unsigned(523, 10), 1276 => to_unsigned(929, 10), 1277 => to_unsigned(903, 10), 1278 => to_unsigned(119, 10), 1279 => to_unsigned(282, 10), 1280 => to_unsigned(560, 10), 1281 => to_unsigned(199, 10), 1282 => to_unsigned(239, 10), 1283 => to_unsigned(694, 10), 1284 => to_unsigned(608, 10), 1285 => to_unsigned(356, 10), 1286 => to_unsigned(850, 10), 1287 => to_unsigned(599, 10), 1288 => to_unsigned(405, 10), 1289 => to_unsigned(510, 10), 1290 => to_unsigned(514, 10), 1291 => to_unsigned(264, 10), 1292 => to_unsigned(266, 10), 1293 => to_unsigned(261, 10), 1294 => to_unsigned(294, 10), 1295 => to_unsigned(934, 10), 1296 => to_unsigned(612, 10), 1297 => to_unsigned(449, 10), 1298 => to_unsigned(629, 10), 1299 => to_unsigned(571, 10), 1300 => to_unsigned(676, 10), 1301 => to_unsigned(901, 10), 1302 => to_unsigned(261, 10), 1303 => to_unsigned(38, 10), 1304 => to_unsigned(675, 10), 1305 => to_unsigned(88, 10), 1306 => to_unsigned(945, 10), 1307 => to_unsigned(719, 10), 1308 => to_unsigned(340, 10), 1309 => to_unsigned(370, 10), 1310 => to_unsigned(265, 10), 1311 => to_unsigned(1015, 10), 1312 => to_unsigned(132, 10), 1313 => to_unsigned(945, 10), 1314 => to_unsigned(24, 10), 1315 => to_unsigned(606, 10), 1316 => to_unsigned(386, 10), 1317 => to_unsigned(851, 10), 1318 => to_unsigned(899, 10), 1319 => to_unsigned(589, 10), 1320 => to_unsigned(267, 10), 1321 => to_unsigned(397, 10), 1322 => to_unsigned(484, 10), 1323 => to_unsigned(81, 10), 1324 => to_unsigned(154, 10), 1325 => to_unsigned(966, 10), 1326 => to_unsigned(687, 10), 1327 => to_unsigned(610, 10), 1328 => to_unsigned(533, 10), 1329 => to_unsigned(916, 10), 1330 => to_unsigned(682, 10), 1331 => to_unsigned(890, 10), 1332 => to_unsigned(441, 10), 1333 => to_unsigned(145, 10), 1334 => to_unsigned(613, 10), 1335 => to_unsigned(985, 10), 1336 => to_unsigned(244, 10), 1337 => to_unsigned(469, 10), 1338 => to_unsigned(183, 10), 1339 => to_unsigned(612, 10), 1340 => to_unsigned(196, 10), 1341 => to_unsigned(111, 10), 1342 => to_unsigned(226, 10), 1343 => to_unsigned(779, 10), 1344 => to_unsigned(994, 10), 1345 => to_unsigned(97, 10), 1346 => to_unsigned(238, 10), 1347 => to_unsigned(403, 10), 1348 => to_unsigned(880, 10), 1349 => to_unsigned(11, 10), 1350 => to_unsigned(993, 10), 1351 => to_unsigned(537, 10), 1352 => to_unsigned(97, 10), 1353 => to_unsigned(351, 10), 1354 => to_unsigned(301, 10), 1355 => to_unsigned(774, 10), 1356 => to_unsigned(601, 10), 1357 => to_unsigned(856, 10), 1358 => to_unsigned(493, 10), 1359 => to_unsigned(550, 10), 1360 => to_unsigned(51, 10), 1361 => to_unsigned(16, 10), 1362 => to_unsigned(919, 10), 1363 => to_unsigned(730, 10), 1364 => to_unsigned(771, 10), 1365 => to_unsigned(858, 10), 1366 => to_unsigned(430, 10), 1367 => to_unsigned(634, 10), 1368 => to_unsigned(413, 10), 1369 => to_unsigned(770, 10), 1370 => to_unsigned(645, 10), 1371 => to_unsigned(377, 10), 1372 => to_unsigned(967, 10), 1373 => to_unsigned(783, 10), 1374 => to_unsigned(846, 10), 1375 => to_unsigned(419, 10), 1376 => to_unsigned(180, 10), 1377 => to_unsigned(359, 10), 1378 => to_unsigned(886, 10), 1379 => to_unsigned(263, 10), 1380 => to_unsigned(691, 10), 1381 => to_unsigned(358, 10), 1382 => to_unsigned(761, 10), 1383 => to_unsigned(947, 10), 1384 => to_unsigned(925, 10), 1385 => to_unsigned(695, 10), 1386 => to_unsigned(625, 10), 1387 => to_unsigned(395, 10), 1388 => to_unsigned(451, 10), 1389 => to_unsigned(717, 10), 1390 => to_unsigned(890, 10), 1391 => to_unsigned(311, 10), 1392 => to_unsigned(600, 10), 1393 => to_unsigned(507, 10), 1394 => to_unsigned(252, 10), 1395 => to_unsigned(504, 10), 1396 => to_unsigned(836, 10), 1397 => to_unsigned(117, 10), 1398 => to_unsigned(371, 10), 1399 => to_unsigned(470, 10), 1400 => to_unsigned(185, 10), 1401 => to_unsigned(349, 10), 1402 => to_unsigned(614, 10), 1403 => to_unsigned(907, 10), 1404 => to_unsigned(718, 10), 1405 => to_unsigned(594, 10), 1406 => to_unsigned(985, 10), 1407 => to_unsigned(236, 10), 1408 => to_unsigned(3, 10), 1409 => to_unsigned(165, 10), 1410 => to_unsigned(391, 10), 1411 => to_unsigned(797, 10), 1412 => to_unsigned(78, 10), 1413 => to_unsigned(779, 10), 1414 => to_unsigned(969, 10), 1415 => to_unsigned(523, 10), 1416 => to_unsigned(784, 10), 1417 => to_unsigned(60, 10), 1418 => to_unsigned(635, 10), 1419 => to_unsigned(103, 10), 1420 => to_unsigned(703, 10), 1421 => to_unsigned(699, 10), 1422 => to_unsigned(129, 10), 1423 => to_unsigned(914, 10), 1424 => to_unsigned(693, 10), 1425 => to_unsigned(284, 10), 1426 => to_unsigned(448, 10), 1427 => to_unsigned(853, 10), 1428 => to_unsigned(728, 10), 1429 => to_unsigned(585, 10), 1430 => to_unsigned(904, 10), 1431 => to_unsigned(978, 10), 1432 => to_unsigned(395, 10), 1433 => to_unsigned(476, 10), 1434 => to_unsigned(373, 10), 1435 => to_unsigned(947, 10), 1436 => to_unsigned(849, 10), 1437 => to_unsigned(439, 10), 1438 => to_unsigned(15, 10), 1439 => to_unsigned(131, 10), 1440 => to_unsigned(106, 10), 1441 => to_unsigned(472, 10), 1442 => to_unsigned(213, 10), 1443 => to_unsigned(284, 10), 1444 => to_unsigned(826, 10), 1445 => to_unsigned(725, 10), 1446 => to_unsigned(590, 10), 1447 => to_unsigned(879, 10), 1448 => to_unsigned(833, 10), 1449 => to_unsigned(844, 10), 1450 => to_unsigned(267, 10), 1451 => to_unsigned(281, 10), 1452 => to_unsigned(359, 10), 1453 => to_unsigned(779, 10), 1454 => to_unsigned(858, 10), 1455 => to_unsigned(749, 10), 1456 => to_unsigned(418, 10), 1457 => to_unsigned(897, 10), 1458 => to_unsigned(1022, 10), 1459 => to_unsigned(656, 10), 1460 => to_unsigned(257, 10), 1461 => to_unsigned(528, 10), 1462 => to_unsigned(545, 10), 1463 => to_unsigned(33, 10), 1464 => to_unsigned(172, 10), 1465 => to_unsigned(486, 10), 1466 => to_unsigned(808, 10), 1467 => to_unsigned(328, 10), 1468 => to_unsigned(205, 10), 1469 => to_unsigned(106, 10), 1470 => to_unsigned(595, 10), 1471 => to_unsigned(754, 10), 1472 => to_unsigned(416, 10), 1473 => to_unsigned(919, 10), 1474 => to_unsigned(324, 10), 1475 => to_unsigned(415, 10), 1476 => to_unsigned(662, 10), 1477 => to_unsigned(64, 10), 1478 => to_unsigned(741, 10), 1479 => to_unsigned(287, 10), 1480 => to_unsigned(79, 10), 1481 => to_unsigned(83, 10), 1482 => to_unsigned(783, 10), 1483 => to_unsigned(819, 10), 1484 => to_unsigned(505, 10), 1485 => to_unsigned(396, 10), 1486 => to_unsigned(685, 10), 1487 => to_unsigned(10, 10), 1488 => to_unsigned(500, 10), 1489 => to_unsigned(617, 10), 1490 => to_unsigned(848, 10), 1491 => to_unsigned(70, 10), 1492 => to_unsigned(21, 10), 1493 => to_unsigned(734, 10), 1494 => to_unsigned(707, 10), 1495 => to_unsigned(336, 10), 1496 => to_unsigned(320, 10), 1497 => to_unsigned(129, 10), 1498 => to_unsigned(818, 10), 1499 => to_unsigned(864, 10), 1500 => to_unsigned(363, 10), 1501 => to_unsigned(1019, 10), 1502 => to_unsigned(466, 10), 1503 => to_unsigned(338, 10), 1504 => to_unsigned(697, 10), 1505 => to_unsigned(406, 10), 1506 => to_unsigned(783, 10), 1507 => to_unsigned(911, 10), 1508 => to_unsigned(540, 10), 1509 => to_unsigned(327, 10), 1510 => to_unsigned(283, 10), 1511 => to_unsigned(216, 10), 1512 => to_unsigned(313, 10), 1513 => to_unsigned(826, 10), 1514 => to_unsigned(216, 10), 1515 => to_unsigned(972, 10), 1516 => to_unsigned(269, 10), 1517 => to_unsigned(914, 10), 1518 => to_unsigned(78, 10), 1519 => to_unsigned(974, 10), 1520 => to_unsigned(788, 10), 1521 => to_unsigned(583, 10), 1522 => to_unsigned(695, 10), 1523 => to_unsigned(300, 10), 1524 => to_unsigned(235, 10), 1525 => to_unsigned(245, 10), 1526 => to_unsigned(91, 10), 1527 => to_unsigned(44, 10), 1528 => to_unsigned(783, 10), 1529 => to_unsigned(1021, 10), 1530 => to_unsigned(599, 10), 1531 => to_unsigned(971, 10), 1532 => to_unsigned(589, 10), 1533 => to_unsigned(510, 10), 1534 => to_unsigned(413, 10), 1535 => to_unsigned(607, 10), 1536 => to_unsigned(110, 10), 1537 => to_unsigned(722, 10), 1538 => to_unsigned(644, 10), 1539 => to_unsigned(540, 10), 1540 => to_unsigned(705, 10), 1541 => to_unsigned(49, 10), 1542 => to_unsigned(945, 10), 1543 => to_unsigned(343, 10), 1544 => to_unsigned(569, 10), 1545 => to_unsigned(720, 10), 1546 => to_unsigned(41, 10), 1547 => to_unsigned(474, 10), 1548 => to_unsigned(752, 10), 1549 => to_unsigned(194, 10), 1550 => to_unsigned(943, 10), 1551 => to_unsigned(273, 10), 1552 => to_unsigned(20, 10), 1553 => to_unsigned(678, 10), 1554 => to_unsigned(320, 10), 1555 => to_unsigned(646, 10), 1556 => to_unsigned(236, 10), 1557 => to_unsigned(662, 10), 1558 => to_unsigned(79, 10), 1559 => to_unsigned(74, 10), 1560 => to_unsigned(162, 10), 1561 => to_unsigned(680, 10), 1562 => to_unsigned(678, 10), 1563 => to_unsigned(1014, 10), 1564 => to_unsigned(661, 10), 1565 => to_unsigned(802, 10), 1566 => to_unsigned(373, 10), 1567 => to_unsigned(160, 10), 1568 => to_unsigned(426, 10), 1569 => to_unsigned(383, 10), 1570 => to_unsigned(300, 10), 1571 => to_unsigned(611, 10), 1572 => to_unsigned(809, 10), 1573 => to_unsigned(761, 10), 1574 => to_unsigned(871, 10), 1575 => to_unsigned(923, 10), 1576 => to_unsigned(763, 10), 1577 => to_unsigned(304, 10), 1578 => to_unsigned(383, 10), 1579 => to_unsigned(650, 10), 1580 => to_unsigned(324, 10), 1581 => to_unsigned(273, 10), 1582 => to_unsigned(771, 10), 1583 => to_unsigned(613, 10), 1584 => to_unsigned(606, 10), 1585 => to_unsigned(471, 10), 1586 => to_unsigned(285, 10), 1587 => to_unsigned(614, 10), 1588 => to_unsigned(635, 10), 1589 => to_unsigned(158, 10), 1590 => to_unsigned(203, 10), 1591 => to_unsigned(450, 10), 1592 => to_unsigned(477, 10), 1593 => to_unsigned(316, 10), 1594 => to_unsigned(647, 10), 1595 => to_unsigned(691, 10), 1596 => to_unsigned(244, 10), 1597 => to_unsigned(585, 10), 1598 => to_unsigned(471, 10), 1599 => to_unsigned(960, 10), 1600 => to_unsigned(1008, 10), 1601 => to_unsigned(401, 10), 1602 => to_unsigned(680, 10), 1603 => to_unsigned(243, 10), 1604 => to_unsigned(533, 10), 1605 => to_unsigned(606, 10), 1606 => to_unsigned(922, 10), 1607 => to_unsigned(143, 10), 1608 => to_unsigned(752, 10), 1609 => to_unsigned(785, 10), 1610 => to_unsigned(266, 10), 1611 => to_unsigned(657, 10), 1612 => to_unsigned(131, 10), 1613 => to_unsigned(999, 10), 1614 => to_unsigned(585, 10), 1615 => to_unsigned(797, 10), 1616 => to_unsigned(195, 10), 1617 => to_unsigned(455, 10), 1618 => to_unsigned(464, 10), 1619 => to_unsigned(226, 10), 1620 => to_unsigned(644, 10), 1621 => to_unsigned(445, 10), 1622 => to_unsigned(858, 10), 1623 => to_unsigned(100, 10), 1624 => to_unsigned(134, 10), 1625 => to_unsigned(32, 10), 1626 => to_unsigned(81, 10), 1627 => to_unsigned(631, 10), 1628 => to_unsigned(374, 10), 1629 => to_unsigned(757, 10), 1630 => to_unsigned(293, 10), 1631 => to_unsigned(631, 10), 1632 => to_unsigned(283, 10), 1633 => to_unsigned(51, 10), 1634 => to_unsigned(590, 10), 1635 => to_unsigned(955, 10), 1636 => to_unsigned(598, 10), 1637 => to_unsigned(607, 10), 1638 => to_unsigned(8, 10), 1639 => to_unsigned(312, 10), 1640 => to_unsigned(797, 10), 1641 => to_unsigned(668, 10), 1642 => to_unsigned(991, 10), 1643 => to_unsigned(418, 10), 1644 => to_unsigned(186, 10), 1645 => to_unsigned(895, 10), 1646 => to_unsigned(894, 10), 1647 => to_unsigned(977, 10), 1648 => to_unsigned(476, 10), 1649 => to_unsigned(111, 10), 1650 => to_unsigned(656, 10), 1651 => to_unsigned(968, 10), 1652 => to_unsigned(571, 10), 1653 => to_unsigned(247, 10), 1654 => to_unsigned(1004, 10), 1655 => to_unsigned(7, 10), 1656 => to_unsigned(908, 10), 1657 => to_unsigned(288, 10), 1658 => to_unsigned(724, 10), 1659 => to_unsigned(747, 10), 1660 => to_unsigned(75, 10), 1661 => to_unsigned(221, 10), 1662 => to_unsigned(40, 10), 1663 => to_unsigned(0, 10), 1664 => to_unsigned(212, 10), 1665 => to_unsigned(109, 10), 1666 => to_unsigned(604, 10), 1667 => to_unsigned(205, 10), 1668 => to_unsigned(165, 10), 1669 => to_unsigned(431, 10), 1670 => to_unsigned(573, 10), 1671 => to_unsigned(103, 10), 1672 => to_unsigned(946, 10), 1673 => to_unsigned(580, 10), 1674 => to_unsigned(494, 10), 1675 => to_unsigned(972, 10), 1676 => to_unsigned(697, 10), 1677 => to_unsigned(887, 10), 1678 => to_unsigned(997, 10), 1679 => to_unsigned(1008, 10), 1680 => to_unsigned(132, 10), 1681 => to_unsigned(617, 10), 1682 => to_unsigned(548, 10), 1683 => to_unsigned(336, 10), 1684 => to_unsigned(466, 10), 1685 => to_unsigned(165, 10), 1686 => to_unsigned(734, 10), 1687 => to_unsigned(373, 10), 1688 => to_unsigned(494, 10), 1689 => to_unsigned(291, 10), 1690 => to_unsigned(944, 10), 1691 => to_unsigned(640, 10), 1692 => to_unsigned(561, 10), 1693 => to_unsigned(185, 10), 1694 => to_unsigned(265, 10), 1695 => to_unsigned(50, 10), 1696 => to_unsigned(737, 10), 1697 => to_unsigned(176, 10), 1698 => to_unsigned(1009, 10), 1699 => to_unsigned(524, 10), 1700 => to_unsigned(710, 10), 1701 => to_unsigned(636, 10), 1702 => to_unsigned(499, 10), 1703 => to_unsigned(932, 10), 1704 => to_unsigned(99, 10), 1705 => to_unsigned(358, 10), 1706 => to_unsigned(36, 10), 1707 => to_unsigned(286, 10), 1708 => to_unsigned(626, 10), 1709 => to_unsigned(147, 10), 1710 => to_unsigned(422, 10), 1711 => to_unsigned(428, 10), 1712 => to_unsigned(35, 10), 1713 => to_unsigned(782, 10), 1714 => to_unsigned(29, 10), 1715 => to_unsigned(947, 10), 1716 => to_unsigned(60, 10), 1717 => to_unsigned(1016, 10), 1718 => to_unsigned(337, 10), 1719 => to_unsigned(835, 10), 1720 => to_unsigned(797, 10), 1721 => to_unsigned(155, 10), 1722 => to_unsigned(131, 10), 1723 => to_unsigned(33, 10), 1724 => to_unsigned(757, 10), 1725 => to_unsigned(435, 10), 1726 => to_unsigned(886, 10), 1727 => to_unsigned(411, 10), 1728 => to_unsigned(228, 10), 1729 => to_unsigned(56, 10), 1730 => to_unsigned(277, 10), 1731 => to_unsigned(679, 10), 1732 => to_unsigned(746, 10), 1733 => to_unsigned(330, 10), 1734 => to_unsigned(541, 10), 1735 => to_unsigned(241, 10), 1736 => to_unsigned(925, 10), 1737 => to_unsigned(957, 10), 1738 => to_unsigned(570, 10), 1739 => to_unsigned(792, 10), 1740 => to_unsigned(114, 10), 1741 => to_unsigned(272, 10), 1742 => to_unsigned(448, 10), 1743 => to_unsigned(868, 10), 1744 => to_unsigned(994, 10), 1745 => to_unsigned(635, 10), 1746 => to_unsigned(13, 10), 1747 => to_unsigned(769, 10), 1748 => to_unsigned(763, 10), 1749 => to_unsigned(258, 10), 1750 => to_unsigned(834, 10), 1751 => to_unsigned(147, 10), 1752 => to_unsigned(500, 10), 1753 => to_unsigned(762, 10), 1754 => to_unsigned(460, 10), 1755 => to_unsigned(670, 10), 1756 => to_unsigned(551, 10), 1757 => to_unsigned(469, 10), 1758 => to_unsigned(589, 10), 1759 => to_unsigned(945, 10), 1760 => to_unsigned(282, 10), 1761 => to_unsigned(371, 10), 1762 => to_unsigned(140, 10), 1763 => to_unsigned(241, 10), 1764 => to_unsigned(960, 10), 1765 => to_unsigned(257, 10), 1766 => to_unsigned(420, 10), 1767 => to_unsigned(778, 10), 1768 => to_unsigned(874, 10), 1769 => to_unsigned(288, 10), 1770 => to_unsigned(510, 10), 1771 => to_unsigned(284, 10), 1772 => to_unsigned(698, 10), 1773 => to_unsigned(706, 10), 1774 => to_unsigned(732, 10), 1775 => to_unsigned(65, 10), 1776 => to_unsigned(205, 10), 1777 => to_unsigned(339, 10), 1778 => to_unsigned(559, 10), 1779 => to_unsigned(593, 10), 1780 => to_unsigned(420, 10), 1781 => to_unsigned(199, 10), 1782 => to_unsigned(309, 10), 1783 => to_unsigned(710, 10), 1784 => to_unsigned(649, 10), 1785 => to_unsigned(527, 10), 1786 => to_unsigned(786, 10), 1787 => to_unsigned(157, 10), 1788 => to_unsigned(693, 10), 1789 => to_unsigned(956, 10), 1790 => to_unsigned(554, 10), 1791 => to_unsigned(466, 10), 1792 => to_unsigned(642, 10), 1793 => to_unsigned(797, 10), 1794 => to_unsigned(401, 10), 1795 => to_unsigned(35, 10), 1796 => to_unsigned(888, 10), 1797 => to_unsigned(275, 10), 1798 => to_unsigned(912, 10), 1799 => to_unsigned(535, 10), 1800 => to_unsigned(652, 10), 1801 => to_unsigned(355, 10), 1802 => to_unsigned(877, 10), 1803 => to_unsigned(696, 10), 1804 => to_unsigned(706, 10), 1805 => to_unsigned(788, 10), 1806 => to_unsigned(131, 10), 1807 => to_unsigned(81, 10), 1808 => to_unsigned(940, 10), 1809 => to_unsigned(38, 10), 1810 => to_unsigned(42, 10), 1811 => to_unsigned(970, 10), 1812 => to_unsigned(549, 10), 1813 => to_unsigned(362, 10), 1814 => to_unsigned(552, 10), 1815 => to_unsigned(879, 10), 1816 => to_unsigned(795, 10), 1817 => to_unsigned(644, 10), 1818 => to_unsigned(435, 10), 1819 => to_unsigned(406, 10), 1820 => to_unsigned(677, 10), 1821 => to_unsigned(803, 10), 1822 => to_unsigned(542, 10), 1823 => to_unsigned(775, 10), 1824 => to_unsigned(984, 10), 1825 => to_unsigned(600, 10), 1826 => to_unsigned(239, 10), 1827 => to_unsigned(911, 10), 1828 => to_unsigned(394, 10), 1829 => to_unsigned(147, 10), 1830 => to_unsigned(845, 10), 1831 => to_unsigned(999, 10), 1832 => to_unsigned(824, 10), 1833 => to_unsigned(997, 10), 1834 => to_unsigned(999, 10), 1835 => to_unsigned(914, 10), 1836 => to_unsigned(455, 10), 1837 => to_unsigned(60, 10), 1838 => to_unsigned(24, 10), 1839 => to_unsigned(160, 10), 1840 => to_unsigned(364, 10), 1841 => to_unsigned(295, 10), 1842 => to_unsigned(884, 10), 1843 => to_unsigned(104, 10), 1844 => to_unsigned(382, 10), 1845 => to_unsigned(367, 10), 1846 => to_unsigned(116, 10), 1847 => to_unsigned(996, 10), 1848 => to_unsigned(1002, 10), 1849 => to_unsigned(16, 10), 1850 => to_unsigned(948, 10), 1851 => to_unsigned(218, 10), 1852 => to_unsigned(1000, 10), 1853 => to_unsigned(208, 10), 1854 => to_unsigned(814, 10), 1855 => to_unsigned(224, 10), 1856 => to_unsigned(606, 10), 1857 => to_unsigned(852, 10), 1858 => to_unsigned(791, 10), 1859 => to_unsigned(655, 10), 1860 => to_unsigned(172, 10), 1861 => to_unsigned(595, 10), 1862 => to_unsigned(119, 10), 1863 => to_unsigned(567, 10), 1864 => to_unsigned(354, 10), 1865 => to_unsigned(411, 10), 1866 => to_unsigned(301, 10), 1867 => to_unsigned(994, 10), 1868 => to_unsigned(337, 10), 1869 => to_unsigned(727, 10), 1870 => to_unsigned(411, 10), 1871 => to_unsigned(589, 10), 1872 => to_unsigned(432, 10), 1873 => to_unsigned(983, 10), 1874 => to_unsigned(862, 10), 1875 => to_unsigned(389, 10), 1876 => to_unsigned(377, 10), 1877 => to_unsigned(231, 10), 1878 => to_unsigned(737, 10), 1879 => to_unsigned(881, 10), 1880 => to_unsigned(994, 10), 1881 => to_unsigned(796, 10), 1882 => to_unsigned(244, 10), 1883 => to_unsigned(65, 10), 1884 => to_unsigned(68, 10), 1885 => to_unsigned(725, 10), 1886 => to_unsigned(456, 10), 1887 => to_unsigned(764, 10), 1888 => to_unsigned(370, 10), 1889 => to_unsigned(929, 10), 1890 => to_unsigned(374, 10), 1891 => to_unsigned(483, 10), 1892 => to_unsigned(560, 10), 1893 => to_unsigned(99, 10), 1894 => to_unsigned(985, 10), 1895 => to_unsigned(581, 10), 1896 => to_unsigned(961, 10), 1897 => to_unsigned(611, 10), 1898 => to_unsigned(71, 10), 1899 => to_unsigned(513, 10), 1900 => to_unsigned(129, 10), 1901 => to_unsigned(199, 10), 1902 => to_unsigned(665, 10), 1903 => to_unsigned(100, 10), 1904 => to_unsigned(589, 10), 1905 => to_unsigned(620, 10), 1906 => to_unsigned(178, 10), 1907 => to_unsigned(411, 10), 1908 => to_unsigned(96, 10), 1909 => to_unsigned(555, 10), 1910 => to_unsigned(787, 10), 1911 => to_unsigned(354, 10), 1912 => to_unsigned(301, 10), 1913 => to_unsigned(100, 10), 1914 => to_unsigned(336, 10), 1915 => to_unsigned(112, 10), 1916 => to_unsigned(234, 10), 1917 => to_unsigned(889, 10), 1918 => to_unsigned(939, 10), 1919 => to_unsigned(451, 10), 1920 => to_unsigned(520, 10), 1921 => to_unsigned(211, 10), 1922 => to_unsigned(942, 10), 1923 => to_unsigned(576, 10), 1924 => to_unsigned(372, 10), 1925 => to_unsigned(916, 10), 1926 => to_unsigned(96, 10), 1927 => to_unsigned(482, 10), 1928 => to_unsigned(875, 10), 1929 => to_unsigned(389, 10), 1930 => to_unsigned(341, 10), 1931 => to_unsigned(280, 10), 1932 => to_unsigned(2, 10), 1933 => to_unsigned(509, 10), 1934 => to_unsigned(1021, 10), 1935 => to_unsigned(455, 10), 1936 => to_unsigned(108, 10), 1937 => to_unsigned(203, 10), 1938 => to_unsigned(243, 10), 1939 => to_unsigned(796, 10), 1940 => to_unsigned(374, 10), 1941 => to_unsigned(863, 10), 1942 => to_unsigned(65, 10), 1943 => to_unsigned(464, 10), 1944 => to_unsigned(370, 10), 1945 => to_unsigned(210, 10), 1946 => to_unsigned(398, 10), 1947 => to_unsigned(533, 10), 1948 => to_unsigned(111, 10), 1949 => to_unsigned(879, 10), 1950 => to_unsigned(197, 10), 1951 => to_unsigned(801, 10), 1952 => to_unsigned(618, 10), 1953 => to_unsigned(130, 10), 1954 => to_unsigned(539, 10), 1955 => to_unsigned(744, 10), 1956 => to_unsigned(375, 10), 1957 => to_unsigned(147, 10), 1958 => to_unsigned(911, 10), 1959 => to_unsigned(839, 10), 1960 => to_unsigned(1004, 10), 1961 => to_unsigned(797, 10), 1962 => to_unsigned(419, 10), 1963 => to_unsigned(737, 10), 1964 => to_unsigned(304, 10), 1965 => to_unsigned(945, 10), 1966 => to_unsigned(848, 10), 1967 => to_unsigned(184, 10), 1968 => to_unsigned(319, 10), 1969 => to_unsigned(472, 10), 1970 => to_unsigned(442, 10), 1971 => to_unsigned(901, 10), 1972 => to_unsigned(819, 10), 1973 => to_unsigned(250, 10), 1974 => to_unsigned(573, 10), 1975 => to_unsigned(106, 10), 1976 => to_unsigned(467, 10), 1977 => to_unsigned(273, 10), 1978 => to_unsigned(45, 10), 1979 => to_unsigned(992, 10), 1980 => to_unsigned(574, 10), 1981 => to_unsigned(22, 10), 1982 => to_unsigned(225, 10), 1983 => to_unsigned(614, 10), 1984 => to_unsigned(649, 10), 1985 => to_unsigned(773, 10), 1986 => to_unsigned(332, 10), 1987 => to_unsigned(573, 10), 1988 => to_unsigned(170, 10), 1989 => to_unsigned(759, 10), 1990 => to_unsigned(400, 10), 1991 => to_unsigned(315, 10), 1992 => to_unsigned(273, 10), 1993 => to_unsigned(196, 10), 1994 => to_unsigned(316, 10), 1995 => to_unsigned(665, 10), 1996 => to_unsigned(142, 10), 1997 => to_unsigned(877, 10), 1998 => to_unsigned(829, 10), 1999 => to_unsigned(181, 10), 2000 => to_unsigned(81, 10), 2001 => to_unsigned(541, 10), 2002 => to_unsigned(198, 10), 2003 => to_unsigned(28, 10), 2004 => to_unsigned(714, 10), 2005 => to_unsigned(645, 10), 2006 => to_unsigned(484, 10), 2007 => to_unsigned(484, 10), 2008 => to_unsigned(340, 10), 2009 => to_unsigned(951, 10), 2010 => to_unsigned(498, 10), 2011 => to_unsigned(178, 10), 2012 => to_unsigned(598, 10), 2013 => to_unsigned(181, 10), 2014 => to_unsigned(778, 10), 2015 => to_unsigned(555, 10), 2016 => to_unsigned(955, 10), 2017 => to_unsigned(414, 10), 2018 => to_unsigned(827, 10), 2019 => to_unsigned(142, 10), 2020 => to_unsigned(1011, 10), 2021 => to_unsigned(432, 10), 2022 => to_unsigned(632, 10), 2023 => to_unsigned(381, 10), 2024 => to_unsigned(56, 10), 2025 => to_unsigned(449, 10), 2026 => to_unsigned(872, 10), 2027 => to_unsigned(903, 10), 2028 => to_unsigned(965, 10), 2029 => to_unsigned(143, 10), 2030 => to_unsigned(631, 10), 2031 => to_unsigned(1001, 10), 2032 => to_unsigned(308, 10), 2033 => to_unsigned(288, 10), 2034 => to_unsigned(87, 10), 2035 => to_unsigned(974, 10), 2036 => to_unsigned(930, 10), 2037 => to_unsigned(541, 10), 2038 => to_unsigned(51, 10), 2039 => to_unsigned(473, 10), 2040 => to_unsigned(437, 10), 2041 => to_unsigned(772, 10), 2042 => to_unsigned(192, 10), 2043 => to_unsigned(891, 10), 2044 => to_unsigned(154, 10), 2045 => to_unsigned(468, 10), 2046 => to_unsigned(389, 10), 2047 => to_unsigned(378, 10)),
            1 => (0 => to_unsigned(856, 10), 1 => to_unsigned(273, 10), 2 => to_unsigned(964, 10), 3 => to_unsigned(312, 10), 4 => to_unsigned(160, 10), 5 => to_unsigned(241, 10), 6 => to_unsigned(337, 10), 7 => to_unsigned(584, 10), 8 => to_unsigned(73, 10), 9 => to_unsigned(740, 10), 10 => to_unsigned(415, 10), 11 => to_unsigned(350, 10), 12 => to_unsigned(329, 10), 13 => to_unsigned(364, 10), 14 => to_unsigned(176, 10), 15 => to_unsigned(739, 10), 16 => to_unsigned(416, 10), 17 => to_unsigned(270, 10), 18 => to_unsigned(573, 10), 19 => to_unsigned(343, 10), 20 => to_unsigned(416, 10), 21 => to_unsigned(312, 10), 22 => to_unsigned(412, 10), 23 => to_unsigned(171, 10), 24 => to_unsigned(97, 10), 25 => to_unsigned(178, 10), 26 => to_unsigned(814, 10), 27 => to_unsigned(108, 10), 28 => to_unsigned(840, 10), 29 => to_unsigned(421, 10), 30 => to_unsigned(632, 10), 31 => to_unsigned(2, 10), 32 => to_unsigned(785, 10), 33 => to_unsigned(143, 10), 34 => to_unsigned(707, 10), 35 => to_unsigned(341, 10), 36 => to_unsigned(496, 10), 37 => to_unsigned(754, 10), 38 => to_unsigned(93, 10), 39 => to_unsigned(869, 10), 40 => to_unsigned(120, 10), 41 => to_unsigned(662, 10), 42 => to_unsigned(210, 10), 43 => to_unsigned(519, 10), 44 => to_unsigned(823, 10), 45 => to_unsigned(177, 10), 46 => to_unsigned(26, 10), 47 => to_unsigned(760, 10), 48 => to_unsigned(644, 10), 49 => to_unsigned(109, 10), 50 => to_unsigned(89, 10), 51 => to_unsigned(26, 10), 52 => to_unsigned(700, 10), 53 => to_unsigned(243, 10), 54 => to_unsigned(623, 10), 55 => to_unsigned(595, 10), 56 => to_unsigned(590, 10), 57 => to_unsigned(658, 10), 58 => to_unsigned(121, 10), 59 => to_unsigned(608, 10), 60 => to_unsigned(347, 10), 61 => to_unsigned(804, 10), 62 => to_unsigned(358, 10), 63 => to_unsigned(404, 10), 64 => to_unsigned(383, 10), 65 => to_unsigned(492, 10), 66 => to_unsigned(387, 10), 67 => to_unsigned(658, 10), 68 => to_unsigned(205, 10), 69 => to_unsigned(51, 10), 70 => to_unsigned(561, 10), 71 => to_unsigned(543, 10), 72 => to_unsigned(481, 10), 73 => to_unsigned(658, 10), 74 => to_unsigned(268, 10), 75 => to_unsigned(623, 10), 76 => to_unsigned(987, 10), 77 => to_unsigned(231, 10), 78 => to_unsigned(866, 10), 79 => to_unsigned(839, 10), 80 => to_unsigned(606, 10), 81 => to_unsigned(813, 10), 82 => to_unsigned(720, 10), 83 => to_unsigned(65, 10), 84 => to_unsigned(88, 10), 85 => to_unsigned(272, 10), 86 => to_unsigned(301, 10), 87 => to_unsigned(383, 10), 88 => to_unsigned(219, 10), 89 => to_unsigned(165, 10), 90 => to_unsigned(434, 10), 91 => to_unsigned(408, 10), 92 => to_unsigned(944, 10), 93 => to_unsigned(204, 10), 94 => to_unsigned(4, 10), 95 => to_unsigned(1008, 10), 96 => to_unsigned(947, 10), 97 => to_unsigned(174, 10), 98 => to_unsigned(40, 10), 99 => to_unsigned(910, 10), 100 => to_unsigned(241, 10), 101 => to_unsigned(394, 10), 102 => to_unsigned(411, 10), 103 => to_unsigned(334, 10), 104 => to_unsigned(870, 10), 105 => to_unsigned(397, 10), 106 => to_unsigned(516, 10), 107 => to_unsigned(726, 10), 108 => to_unsigned(271, 10), 109 => to_unsigned(29, 10), 110 => to_unsigned(974, 10), 111 => to_unsigned(170, 10), 112 => to_unsigned(665, 10), 113 => to_unsigned(203, 10), 114 => to_unsigned(479, 10), 115 => to_unsigned(219, 10), 116 => to_unsigned(534, 10), 117 => to_unsigned(110, 10), 118 => to_unsigned(811, 10), 119 => to_unsigned(468, 10), 120 => to_unsigned(695, 10), 121 => to_unsigned(765, 10), 122 => to_unsigned(130, 10), 123 => to_unsigned(665, 10), 124 => to_unsigned(637, 10), 125 => to_unsigned(120, 10), 126 => to_unsigned(640, 10), 127 => to_unsigned(351, 10), 128 => to_unsigned(184, 10), 129 => to_unsigned(110, 10), 130 => to_unsigned(710, 10), 131 => to_unsigned(978, 10), 132 => to_unsigned(598, 10), 133 => to_unsigned(190, 10), 134 => to_unsigned(767, 10), 135 => to_unsigned(558, 10), 136 => to_unsigned(763, 10), 137 => to_unsigned(89, 10), 138 => to_unsigned(717, 10), 139 => to_unsigned(652, 10), 140 => to_unsigned(318, 10), 141 => to_unsigned(293, 10), 142 => to_unsigned(979, 10), 143 => to_unsigned(159, 10), 144 => to_unsigned(887, 10), 145 => to_unsigned(924, 10), 146 => to_unsigned(315, 10), 147 => to_unsigned(504, 10), 148 => to_unsigned(339, 10), 149 => to_unsigned(808, 10), 150 => to_unsigned(360, 10), 151 => to_unsigned(377, 10), 152 => to_unsigned(601, 10), 153 => to_unsigned(1007, 10), 154 => to_unsigned(797, 10), 155 => to_unsigned(796, 10), 156 => to_unsigned(52, 10), 157 => to_unsigned(298, 10), 158 => to_unsigned(650, 10), 159 => to_unsigned(724, 10), 160 => to_unsigned(273, 10), 161 => to_unsigned(640, 10), 162 => to_unsigned(679, 10), 163 => to_unsigned(38, 10), 164 => to_unsigned(482, 10), 165 => to_unsigned(193, 10), 166 => to_unsigned(560, 10), 167 => to_unsigned(214, 10), 168 => to_unsigned(45, 10), 169 => to_unsigned(122, 10), 170 => to_unsigned(689, 10), 171 => to_unsigned(534, 10), 172 => to_unsigned(231, 10), 173 => to_unsigned(510, 10), 174 => to_unsigned(348, 10), 175 => to_unsigned(321, 10), 176 => to_unsigned(341, 10), 177 => to_unsigned(834, 10), 178 => to_unsigned(544, 10), 179 => to_unsigned(434, 10), 180 => to_unsigned(326, 10), 181 => to_unsigned(614, 10), 182 => to_unsigned(931, 10), 183 => to_unsigned(1013, 10), 184 => to_unsigned(484, 10), 185 => to_unsigned(151, 10), 186 => to_unsigned(1011, 10), 187 => to_unsigned(122, 10), 188 => to_unsigned(82, 10), 189 => to_unsigned(102, 10), 190 => to_unsigned(89, 10), 191 => to_unsigned(750, 10), 192 => to_unsigned(79, 10), 193 => to_unsigned(113, 10), 194 => to_unsigned(155, 10), 195 => to_unsigned(853, 10), 196 => to_unsigned(513, 10), 197 => to_unsigned(265, 10), 198 => to_unsigned(115, 10), 199 => to_unsigned(849, 10), 200 => to_unsigned(395, 10), 201 => to_unsigned(64, 10), 202 => to_unsigned(247, 10), 203 => to_unsigned(835, 10), 204 => to_unsigned(505, 10), 205 => to_unsigned(189, 10), 206 => to_unsigned(54, 10), 207 => to_unsigned(292, 10), 208 => to_unsigned(468, 10), 209 => to_unsigned(126, 10), 210 => to_unsigned(19, 10), 211 => to_unsigned(1007, 10), 212 => to_unsigned(709, 10), 213 => to_unsigned(724, 10), 214 => to_unsigned(637, 10), 215 => to_unsigned(702, 10), 216 => to_unsigned(196, 10), 217 => to_unsigned(169, 10), 218 => to_unsigned(208, 10), 219 => to_unsigned(656, 10), 220 => to_unsigned(185, 10), 221 => to_unsigned(645, 10), 222 => to_unsigned(96, 10), 223 => to_unsigned(278, 10), 224 => to_unsigned(131, 10), 225 => to_unsigned(392, 10), 226 => to_unsigned(830, 10), 227 => to_unsigned(860, 10), 228 => to_unsigned(169, 10), 229 => to_unsigned(842, 10), 230 => to_unsigned(102, 10), 231 => to_unsigned(604, 10), 232 => to_unsigned(95, 10), 233 => to_unsigned(108, 10), 234 => to_unsigned(907, 10), 235 => to_unsigned(930, 10), 236 => to_unsigned(91, 10), 237 => to_unsigned(817, 10), 238 => to_unsigned(583, 10), 239 => to_unsigned(423, 10), 240 => to_unsigned(870, 10), 241 => to_unsigned(887, 10), 242 => to_unsigned(58, 10), 243 => to_unsigned(5, 10), 244 => to_unsigned(73, 10), 245 => to_unsigned(856, 10), 246 => to_unsigned(140, 10), 247 => to_unsigned(744, 10), 248 => to_unsigned(225, 10), 249 => to_unsigned(827, 10), 250 => to_unsigned(718, 10), 251 => to_unsigned(1005, 10), 252 => to_unsigned(527, 10), 253 => to_unsigned(4, 10), 254 => to_unsigned(918, 10), 255 => to_unsigned(692, 10), 256 => to_unsigned(66, 10), 257 => to_unsigned(839, 10), 258 => to_unsigned(365, 10), 259 => to_unsigned(328, 10), 260 => to_unsigned(261, 10), 261 => to_unsigned(551, 10), 262 => to_unsigned(335, 10), 263 => to_unsigned(847, 10), 264 => to_unsigned(809, 10), 265 => to_unsigned(985, 10), 266 => to_unsigned(662, 10), 267 => to_unsigned(473, 10), 268 => to_unsigned(217, 10), 269 => to_unsigned(915, 10), 270 => to_unsigned(830, 10), 271 => to_unsigned(797, 10), 272 => to_unsigned(777, 10), 273 => to_unsigned(395, 10), 274 => to_unsigned(893, 10), 275 => to_unsigned(99, 10), 276 => to_unsigned(538, 10), 277 => to_unsigned(871, 10), 278 => to_unsigned(255, 10), 279 => to_unsigned(722, 10), 280 => to_unsigned(584, 10), 281 => to_unsigned(255, 10), 282 => to_unsigned(641, 10), 283 => to_unsigned(867, 10), 284 => to_unsigned(626, 10), 285 => to_unsigned(241, 10), 286 => to_unsigned(686, 10), 287 => to_unsigned(311, 10), 288 => to_unsigned(522, 10), 289 => to_unsigned(714, 10), 290 => to_unsigned(280, 10), 291 => to_unsigned(511, 10), 292 => to_unsigned(351, 10), 293 => to_unsigned(43, 10), 294 => to_unsigned(987, 10), 295 => to_unsigned(653, 10), 296 => to_unsigned(974, 10), 297 => to_unsigned(55, 10), 298 => to_unsigned(5, 10), 299 => to_unsigned(407, 10), 300 => to_unsigned(42, 10), 301 => to_unsigned(615, 10), 302 => to_unsigned(49, 10), 303 => to_unsigned(357, 10), 304 => to_unsigned(870, 10), 305 => to_unsigned(587, 10), 306 => to_unsigned(885, 10), 307 => to_unsigned(952, 10), 308 => to_unsigned(427, 10), 309 => to_unsigned(152, 10), 310 => to_unsigned(337, 10), 311 => to_unsigned(533, 10), 312 => to_unsigned(990, 10), 313 => to_unsigned(146, 10), 314 => to_unsigned(63, 10), 315 => to_unsigned(345, 10), 316 => to_unsigned(541, 10), 317 => to_unsigned(293, 10), 318 => to_unsigned(945, 10), 319 => to_unsigned(168, 10), 320 => to_unsigned(497, 10), 321 => to_unsigned(362, 10), 322 => to_unsigned(223, 10), 323 => to_unsigned(103, 10), 324 => to_unsigned(267, 10), 325 => to_unsigned(312, 10), 326 => to_unsigned(1013, 10), 327 => to_unsigned(447, 10), 328 => to_unsigned(142, 10), 329 => to_unsigned(288, 10), 330 => to_unsigned(193, 10), 331 => to_unsigned(121, 10), 332 => to_unsigned(373, 10), 333 => to_unsigned(833, 10), 334 => to_unsigned(36, 10), 335 => to_unsigned(762, 10), 336 => to_unsigned(25, 10), 337 => to_unsigned(972, 10), 338 => to_unsigned(72, 10), 339 => to_unsigned(50, 10), 340 => to_unsigned(524, 10), 341 => to_unsigned(920, 10), 342 => to_unsigned(147, 10), 343 => to_unsigned(707, 10), 344 => to_unsigned(394, 10), 345 => to_unsigned(519, 10), 346 => to_unsigned(948, 10), 347 => to_unsigned(92, 10), 348 => to_unsigned(526, 10), 349 => to_unsigned(456, 10), 350 => to_unsigned(46, 10), 351 => to_unsigned(227, 10), 352 => to_unsigned(35, 10), 353 => to_unsigned(209, 10), 354 => to_unsigned(151, 10), 355 => to_unsigned(61, 10), 356 => to_unsigned(629, 10), 357 => to_unsigned(181, 10), 358 => to_unsigned(524, 10), 359 => to_unsigned(429, 10), 360 => to_unsigned(519, 10), 361 => to_unsigned(506, 10), 362 => to_unsigned(431, 10), 363 => to_unsigned(110, 10), 364 => to_unsigned(679, 10), 365 => to_unsigned(862, 10), 366 => to_unsigned(659, 10), 367 => to_unsigned(234, 10), 368 => to_unsigned(877, 10), 369 => to_unsigned(946, 10), 370 => to_unsigned(577, 10), 371 => to_unsigned(939, 10), 372 => to_unsigned(594, 10), 373 => to_unsigned(462, 10), 374 => to_unsigned(1019, 10), 375 => to_unsigned(89, 10), 376 => to_unsigned(101, 10), 377 => to_unsigned(376, 10), 378 => to_unsigned(184, 10), 379 => to_unsigned(584, 10), 380 => to_unsigned(690, 10), 381 => to_unsigned(34, 10), 382 => to_unsigned(986, 10), 383 => to_unsigned(523, 10), 384 => to_unsigned(620, 10), 385 => to_unsigned(139, 10), 386 => to_unsigned(360, 10), 387 => to_unsigned(420, 10), 388 => to_unsigned(894, 10), 389 => to_unsigned(177, 10), 390 => to_unsigned(972, 10), 391 => to_unsigned(977, 10), 392 => to_unsigned(223, 10), 393 => to_unsigned(970, 10), 394 => to_unsigned(816, 10), 395 => to_unsigned(586, 10), 396 => to_unsigned(139, 10), 397 => to_unsigned(605, 10), 398 => to_unsigned(546, 10), 399 => to_unsigned(714, 10), 400 => to_unsigned(460, 10), 401 => to_unsigned(753, 10), 402 => to_unsigned(295, 10), 403 => to_unsigned(368, 10), 404 => to_unsigned(522, 10), 405 => to_unsigned(770, 10), 406 => to_unsigned(377, 10), 407 => to_unsigned(1007, 10), 408 => to_unsigned(75, 10), 409 => to_unsigned(942, 10), 410 => to_unsigned(51, 10), 411 => to_unsigned(500, 10), 412 => to_unsigned(937, 10), 413 => to_unsigned(1018, 10), 414 => to_unsigned(91, 10), 415 => to_unsigned(643, 10), 416 => to_unsigned(272, 10), 417 => to_unsigned(319, 10), 418 => to_unsigned(832, 10), 419 => to_unsigned(781, 10), 420 => to_unsigned(806, 10), 421 => to_unsigned(260, 10), 422 => to_unsigned(515, 10), 423 => to_unsigned(915, 10), 424 => to_unsigned(593, 10), 425 => to_unsigned(144, 10), 426 => to_unsigned(382, 10), 427 => to_unsigned(839, 10), 428 => to_unsigned(664, 10), 429 => to_unsigned(267, 10), 430 => to_unsigned(150, 10), 431 => to_unsigned(572, 10), 432 => to_unsigned(219, 10), 433 => to_unsigned(642, 10), 434 => to_unsigned(904, 10), 435 => to_unsigned(72, 10), 436 => to_unsigned(729, 10), 437 => to_unsigned(294, 10), 438 => to_unsigned(564, 10), 439 => to_unsigned(737, 10), 440 => to_unsigned(344, 10), 441 => to_unsigned(319, 10), 442 => to_unsigned(917, 10), 443 => to_unsigned(516, 10), 444 => to_unsigned(415, 10), 445 => to_unsigned(755, 10), 446 => to_unsigned(203, 10), 447 => to_unsigned(677, 10), 448 => to_unsigned(775, 10), 449 => to_unsigned(662, 10), 450 => to_unsigned(636, 10), 451 => to_unsigned(298, 10), 452 => to_unsigned(187, 10), 453 => to_unsigned(735, 10), 454 => to_unsigned(310, 10), 455 => to_unsigned(969, 10), 456 => to_unsigned(883, 10), 457 => to_unsigned(435, 10), 458 => to_unsigned(594, 10), 459 => to_unsigned(791, 10), 460 => to_unsigned(83, 10), 461 => to_unsigned(793, 10), 462 => to_unsigned(825, 10), 463 => to_unsigned(197, 10), 464 => to_unsigned(345, 10), 465 => to_unsigned(301, 10), 466 => to_unsigned(367, 10), 467 => to_unsigned(600, 10), 468 => to_unsigned(947, 10), 469 => to_unsigned(315, 10), 470 => to_unsigned(940, 10), 471 => to_unsigned(154, 10), 472 => to_unsigned(632, 10), 473 => to_unsigned(629, 10), 474 => to_unsigned(939, 10), 475 => to_unsigned(633, 10), 476 => to_unsigned(416, 10), 477 => to_unsigned(798, 10), 478 => to_unsigned(654, 10), 479 => to_unsigned(327, 10), 480 => to_unsigned(96, 10), 481 => to_unsigned(701, 10), 482 => to_unsigned(513, 10), 483 => to_unsigned(502, 10), 484 => to_unsigned(431, 10), 485 => to_unsigned(380, 10), 486 => to_unsigned(365, 10), 487 => to_unsigned(118, 10), 488 => to_unsigned(171, 10), 489 => to_unsigned(474, 10), 490 => to_unsigned(15, 10), 491 => to_unsigned(836, 10), 492 => to_unsigned(202, 10), 493 => to_unsigned(85, 10), 494 => to_unsigned(679, 10), 495 => to_unsigned(106, 10), 496 => to_unsigned(491, 10), 497 => to_unsigned(606, 10), 498 => to_unsigned(470, 10), 499 => to_unsigned(256, 10), 500 => to_unsigned(593, 10), 501 => to_unsigned(186, 10), 502 => to_unsigned(12, 10), 503 => to_unsigned(219, 10), 504 => to_unsigned(811, 10), 505 => to_unsigned(950, 10), 506 => to_unsigned(381, 10), 507 => to_unsigned(431, 10), 508 => to_unsigned(790, 10), 509 => to_unsigned(799, 10), 510 => to_unsigned(372, 10), 511 => to_unsigned(34, 10), 512 => to_unsigned(994, 10), 513 => to_unsigned(810, 10), 514 => to_unsigned(324, 10), 515 => to_unsigned(890, 10), 516 => to_unsigned(830, 10), 517 => to_unsigned(804, 10), 518 => to_unsigned(851, 10), 519 => to_unsigned(172, 10), 520 => to_unsigned(721, 10), 521 => to_unsigned(240, 10), 522 => to_unsigned(367, 10), 523 => to_unsigned(198, 10), 524 => to_unsigned(262, 10), 525 => to_unsigned(432, 10), 526 => to_unsigned(393, 10), 527 => to_unsigned(540, 10), 528 => to_unsigned(77, 10), 529 => to_unsigned(696, 10), 530 => to_unsigned(393, 10), 531 => to_unsigned(469, 10), 532 => to_unsigned(834, 10), 533 => to_unsigned(521, 10), 534 => to_unsigned(110, 10), 535 => to_unsigned(1016, 10), 536 => to_unsigned(164, 10), 537 => to_unsigned(284, 10), 538 => to_unsigned(500, 10), 539 => to_unsigned(64, 10), 540 => to_unsigned(970, 10), 541 => to_unsigned(892, 10), 542 => to_unsigned(141, 10), 543 => to_unsigned(235, 10), 544 => to_unsigned(514, 10), 545 => to_unsigned(421, 10), 546 => to_unsigned(967, 10), 547 => to_unsigned(87, 10), 548 => to_unsigned(734, 10), 549 => to_unsigned(977, 10), 550 => to_unsigned(515, 10), 551 => to_unsigned(111, 10), 552 => to_unsigned(994, 10), 553 => to_unsigned(848, 10), 554 => to_unsigned(755, 10), 555 => to_unsigned(594, 10), 556 => to_unsigned(818, 10), 557 => to_unsigned(957, 10), 558 => to_unsigned(490, 10), 559 => to_unsigned(978, 10), 560 => to_unsigned(28, 10), 561 => to_unsigned(803, 10), 562 => to_unsigned(309, 10), 563 => to_unsigned(794, 10), 564 => to_unsigned(369, 10), 565 => to_unsigned(359, 10), 566 => to_unsigned(554, 10), 567 => to_unsigned(814, 10), 568 => to_unsigned(197, 10), 569 => to_unsigned(540, 10), 570 => to_unsigned(127, 10), 571 => to_unsigned(171, 10), 572 => to_unsigned(83, 10), 573 => to_unsigned(62, 10), 574 => to_unsigned(842, 10), 575 => to_unsigned(202, 10), 576 => to_unsigned(649, 10), 577 => to_unsigned(219, 10), 578 => to_unsigned(739, 10), 579 => to_unsigned(843, 10), 580 => to_unsigned(864, 10), 581 => to_unsigned(166, 10), 582 => to_unsigned(31, 10), 583 => to_unsigned(755, 10), 584 => to_unsigned(918, 10), 585 => to_unsigned(382, 10), 586 => to_unsigned(859, 10), 587 => to_unsigned(825, 10), 588 => to_unsigned(21, 10), 589 => to_unsigned(737, 10), 590 => to_unsigned(829, 10), 591 => to_unsigned(492, 10), 592 => to_unsigned(809, 10), 593 => to_unsigned(371, 10), 594 => to_unsigned(875, 10), 595 => to_unsigned(355, 10), 596 => to_unsigned(169, 10), 597 => to_unsigned(250, 10), 598 => to_unsigned(663, 10), 599 => to_unsigned(253, 10), 600 => to_unsigned(744, 10), 601 => to_unsigned(820, 10), 602 => to_unsigned(279, 10), 603 => to_unsigned(122, 10), 604 => to_unsigned(840, 10), 605 => to_unsigned(553, 10), 606 => to_unsigned(237, 10), 607 => to_unsigned(828, 10), 608 => to_unsigned(815, 10), 609 => to_unsigned(655, 10), 610 => to_unsigned(36, 10), 611 => to_unsigned(961, 10), 612 => to_unsigned(606, 10), 613 => to_unsigned(997, 10), 614 => to_unsigned(810, 10), 615 => to_unsigned(766, 10), 616 => to_unsigned(512, 10), 617 => to_unsigned(979, 10), 618 => to_unsigned(902, 10), 619 => to_unsigned(733, 10), 620 => to_unsigned(67, 10), 621 => to_unsigned(287, 10), 622 => to_unsigned(797, 10), 623 => to_unsigned(16, 10), 624 => to_unsigned(963, 10), 625 => to_unsigned(282, 10), 626 => to_unsigned(1021, 10), 627 => to_unsigned(262, 10), 628 => to_unsigned(233, 10), 629 => to_unsigned(485, 10), 630 => to_unsigned(267, 10), 631 => to_unsigned(337, 10), 632 => to_unsigned(823, 10), 633 => to_unsigned(893, 10), 634 => to_unsigned(299, 10), 635 => to_unsigned(323, 10), 636 => to_unsigned(532, 10), 637 => to_unsigned(475, 10), 638 => to_unsigned(511, 10), 639 => to_unsigned(631, 10), 640 => to_unsigned(476, 10), 641 => to_unsigned(270, 10), 642 => to_unsigned(270, 10), 643 => to_unsigned(80, 10), 644 => to_unsigned(483, 10), 645 => to_unsigned(447, 10), 646 => to_unsigned(373, 10), 647 => to_unsigned(742, 10), 648 => to_unsigned(43, 10), 649 => to_unsigned(155, 10), 650 => to_unsigned(358, 10), 651 => to_unsigned(727, 10), 652 => to_unsigned(916, 10), 653 => to_unsigned(1019, 10), 654 => to_unsigned(535, 10), 655 => to_unsigned(290, 10), 656 => to_unsigned(288, 10), 657 => to_unsigned(833, 10), 658 => to_unsigned(278, 10), 659 => to_unsigned(789, 10), 660 => to_unsigned(441, 10), 661 => to_unsigned(580, 10), 662 => to_unsigned(813, 10), 663 => to_unsigned(1000, 10), 664 => to_unsigned(935, 10), 665 => to_unsigned(792, 10), 666 => to_unsigned(342, 10), 667 => to_unsigned(273, 10), 668 => to_unsigned(948, 10), 669 => to_unsigned(474, 10), 670 => to_unsigned(648, 10), 671 => to_unsigned(773, 10), 672 => to_unsigned(225, 10), 673 => to_unsigned(342, 10), 674 => to_unsigned(250, 10), 675 => to_unsigned(594, 10), 676 => to_unsigned(778, 10), 677 => to_unsigned(574, 10), 678 => to_unsigned(541, 10), 679 => to_unsigned(139, 10), 680 => to_unsigned(158, 10), 681 => to_unsigned(327, 10), 682 => to_unsigned(570, 10), 683 => to_unsigned(990, 10), 684 => to_unsigned(42, 10), 685 => to_unsigned(981, 10), 686 => to_unsigned(327, 10), 687 => to_unsigned(665, 10), 688 => to_unsigned(492, 10), 689 => to_unsigned(822, 10), 690 => to_unsigned(118, 10), 691 => to_unsigned(339, 10), 692 => to_unsigned(25, 10), 693 => to_unsigned(173, 10), 694 => to_unsigned(377, 10), 695 => to_unsigned(490, 10), 696 => to_unsigned(131, 10), 697 => to_unsigned(884, 10), 698 => to_unsigned(980, 10), 699 => to_unsigned(1009, 10), 700 => to_unsigned(851, 10), 701 => to_unsigned(249, 10), 702 => to_unsigned(549, 10), 703 => to_unsigned(161, 10), 704 => to_unsigned(444, 10), 705 => to_unsigned(876, 10), 706 => to_unsigned(729, 10), 707 => to_unsigned(519, 10), 708 => to_unsigned(956, 10), 709 => to_unsigned(165, 10), 710 => to_unsigned(596, 10), 711 => to_unsigned(1018, 10), 712 => to_unsigned(354, 10), 713 => to_unsigned(272, 10), 714 => to_unsigned(685, 10), 715 => to_unsigned(488, 10), 716 => to_unsigned(167, 10), 717 => to_unsigned(545, 10), 718 => to_unsigned(865, 10), 719 => to_unsigned(833, 10), 720 => to_unsigned(201, 10), 721 => to_unsigned(87, 10), 722 => to_unsigned(324, 10), 723 => to_unsigned(280, 10), 724 => to_unsigned(6, 10), 725 => to_unsigned(865, 10), 726 => to_unsigned(370, 10), 727 => to_unsigned(767, 10), 728 => to_unsigned(572, 10), 729 => to_unsigned(216, 10), 730 => to_unsigned(61, 10), 731 => to_unsigned(1012, 10), 732 => to_unsigned(187, 10), 733 => to_unsigned(503, 10), 734 => to_unsigned(633, 10), 735 => to_unsigned(458, 10), 736 => to_unsigned(797, 10), 737 => to_unsigned(239, 10), 738 => to_unsigned(1016, 10), 739 => to_unsigned(28, 10), 740 => to_unsigned(152, 10), 741 => to_unsigned(387, 10), 742 => to_unsigned(466, 10), 743 => to_unsigned(661, 10), 744 => to_unsigned(262, 10), 745 => to_unsigned(84, 10), 746 => to_unsigned(277, 10), 747 => to_unsigned(631, 10), 748 => to_unsigned(283, 10), 749 => to_unsigned(922, 10), 750 => to_unsigned(985, 10), 751 => to_unsigned(448, 10), 752 => to_unsigned(366, 10), 753 => to_unsigned(387, 10), 754 => to_unsigned(821, 10), 755 => to_unsigned(805, 10), 756 => to_unsigned(7, 10), 757 => to_unsigned(376, 10), 758 => to_unsigned(336, 10), 759 => to_unsigned(459, 10), 760 => to_unsigned(651, 10), 761 => to_unsigned(1004, 10), 762 => to_unsigned(386, 10), 763 => to_unsigned(310, 10), 764 => to_unsigned(517, 10), 765 => to_unsigned(785, 10), 766 => to_unsigned(762, 10), 767 => to_unsigned(893, 10), 768 => to_unsigned(590, 10), 769 => to_unsigned(901, 10), 770 => to_unsigned(846, 10), 771 => to_unsigned(81, 10), 772 => to_unsigned(233, 10), 773 => to_unsigned(110, 10), 774 => to_unsigned(620, 10), 775 => to_unsigned(30, 10), 776 => to_unsigned(866, 10), 777 => to_unsigned(771, 10), 778 => to_unsigned(128, 10), 779 => to_unsigned(861, 10), 780 => to_unsigned(300, 10), 781 => to_unsigned(684, 10), 782 => to_unsigned(236, 10), 783 => to_unsigned(895, 10), 784 => to_unsigned(627, 10), 785 => to_unsigned(957, 10), 786 => to_unsigned(254, 10), 787 => to_unsigned(0, 10), 788 => to_unsigned(785, 10), 789 => to_unsigned(413, 10), 790 => to_unsigned(603, 10), 791 => to_unsigned(930, 10), 792 => to_unsigned(1010, 10), 793 => to_unsigned(1011, 10), 794 => to_unsigned(228, 10), 795 => to_unsigned(187, 10), 796 => to_unsigned(21, 10), 797 => to_unsigned(63, 10), 798 => to_unsigned(734, 10), 799 => to_unsigned(504, 10), 800 => to_unsigned(613, 10), 801 => to_unsigned(657, 10), 802 => to_unsigned(38, 10), 803 => to_unsigned(719, 10), 804 => to_unsigned(897, 10), 805 => to_unsigned(143, 10), 806 => to_unsigned(1001, 10), 807 => to_unsigned(726, 10), 808 => to_unsigned(749, 10), 809 => to_unsigned(529, 10), 810 => to_unsigned(236, 10), 811 => to_unsigned(949, 10), 812 => to_unsigned(406, 10), 813 => to_unsigned(461, 10), 814 => to_unsigned(626, 10), 815 => to_unsigned(175, 10), 816 => to_unsigned(706, 10), 817 => to_unsigned(267, 10), 818 => to_unsigned(905, 10), 819 => to_unsigned(498, 10), 820 => to_unsigned(808, 10), 821 => to_unsigned(950, 10), 822 => to_unsigned(947, 10), 823 => to_unsigned(47, 10), 824 => to_unsigned(772, 10), 825 => to_unsigned(906, 10), 826 => to_unsigned(497, 10), 827 => to_unsigned(254, 10), 828 => to_unsigned(646, 10), 829 => to_unsigned(374, 10), 830 => to_unsigned(428, 10), 831 => to_unsigned(328, 10), 832 => to_unsigned(392, 10), 833 => to_unsigned(200, 10), 834 => to_unsigned(492, 10), 835 => to_unsigned(741, 10), 836 => to_unsigned(18, 10), 837 => to_unsigned(2, 10), 838 => to_unsigned(197, 10), 839 => to_unsigned(221, 10), 840 => to_unsigned(505, 10), 841 => to_unsigned(229, 10), 842 => to_unsigned(612, 10), 843 => to_unsigned(362, 10), 844 => to_unsigned(157, 10), 845 => to_unsigned(155, 10), 846 => to_unsigned(657, 10), 847 => to_unsigned(442, 10), 848 => to_unsigned(395, 10), 849 => to_unsigned(305, 10), 850 => to_unsigned(328, 10), 851 => to_unsigned(344, 10), 852 => to_unsigned(515, 10), 853 => to_unsigned(624, 10), 854 => to_unsigned(11, 10), 855 => to_unsigned(825, 10), 856 => to_unsigned(434, 10), 857 => to_unsigned(655, 10), 858 => to_unsigned(953, 10), 859 => to_unsigned(131, 10), 860 => to_unsigned(886, 10), 861 => to_unsigned(996, 10), 862 => to_unsigned(956, 10), 863 => to_unsigned(935, 10), 864 => to_unsigned(510, 10), 865 => to_unsigned(981, 10), 866 => to_unsigned(157, 10), 867 => to_unsigned(949, 10), 868 => to_unsigned(67, 10), 869 => to_unsigned(568, 10), 870 => to_unsigned(203, 10), 871 => to_unsigned(375, 10), 872 => to_unsigned(79, 10), 873 => to_unsigned(301, 10), 874 => to_unsigned(602, 10), 875 => to_unsigned(79, 10), 876 => to_unsigned(225, 10), 877 => to_unsigned(11, 10), 878 => to_unsigned(503, 10), 879 => to_unsigned(133, 10), 880 => to_unsigned(926, 10), 881 => to_unsigned(186, 10), 882 => to_unsigned(580, 10), 883 => to_unsigned(315, 10), 884 => to_unsigned(544, 10), 885 => to_unsigned(805, 10), 886 => to_unsigned(171, 10), 887 => to_unsigned(637, 10), 888 => to_unsigned(316, 10), 889 => to_unsigned(557, 10), 890 => to_unsigned(285, 10), 891 => to_unsigned(250, 10), 892 => to_unsigned(155, 10), 893 => to_unsigned(743, 10), 894 => to_unsigned(795, 10), 895 => to_unsigned(29, 10), 896 => to_unsigned(126, 10), 897 => to_unsigned(72, 10), 898 => to_unsigned(75, 10), 899 => to_unsigned(97, 10), 900 => to_unsigned(206, 10), 901 => to_unsigned(550, 10), 902 => to_unsigned(267, 10), 903 => to_unsigned(458, 10), 904 => to_unsigned(758, 10), 905 => to_unsigned(857, 10), 906 => to_unsigned(32, 10), 907 => to_unsigned(690, 10), 908 => to_unsigned(40, 10), 909 => to_unsigned(198, 10), 910 => to_unsigned(286, 10), 911 => to_unsigned(662, 10), 912 => to_unsigned(123, 10), 913 => to_unsigned(587, 10), 914 => to_unsigned(291, 10), 915 => to_unsigned(468, 10), 916 => to_unsigned(964, 10), 917 => to_unsigned(575, 10), 918 => to_unsigned(772, 10), 919 => to_unsigned(689, 10), 920 => to_unsigned(884, 10), 921 => to_unsigned(157, 10), 922 => to_unsigned(703, 10), 923 => to_unsigned(829, 10), 924 => to_unsigned(603, 10), 925 => to_unsigned(623, 10), 926 => to_unsigned(211, 10), 927 => to_unsigned(360, 10), 928 => to_unsigned(90, 10), 929 => to_unsigned(538, 10), 930 => to_unsigned(585, 10), 931 => to_unsigned(946, 10), 932 => to_unsigned(223, 10), 933 => to_unsigned(862, 10), 934 => to_unsigned(785, 10), 935 => to_unsigned(711, 10), 936 => to_unsigned(824, 10), 937 => to_unsigned(1011, 10), 938 => to_unsigned(803, 10), 939 => to_unsigned(201, 10), 940 => to_unsigned(732, 10), 941 => to_unsigned(815, 10), 942 => to_unsigned(48, 10), 943 => to_unsigned(375, 10), 944 => to_unsigned(967, 10), 945 => to_unsigned(629, 10), 946 => to_unsigned(579, 10), 947 => to_unsigned(635, 10), 948 => to_unsigned(711, 10), 949 => to_unsigned(318, 10), 950 => to_unsigned(968, 10), 951 => to_unsigned(293, 10), 952 => to_unsigned(5, 10), 953 => to_unsigned(609, 10), 954 => to_unsigned(55, 10), 955 => to_unsigned(476, 10), 956 => to_unsigned(430, 10), 957 => to_unsigned(38, 10), 958 => to_unsigned(561, 10), 959 => to_unsigned(264, 10), 960 => to_unsigned(634, 10), 961 => to_unsigned(193, 10), 962 => to_unsigned(322, 10), 963 => to_unsigned(62, 10), 964 => to_unsigned(16, 10), 965 => to_unsigned(189, 10), 966 => to_unsigned(194, 10), 967 => to_unsigned(267, 10), 968 => to_unsigned(415, 10), 969 => to_unsigned(394, 10), 970 => to_unsigned(20, 10), 971 => to_unsigned(100, 10), 972 => to_unsigned(782, 10), 973 => to_unsigned(632, 10), 974 => to_unsigned(52, 10), 975 => to_unsigned(455, 10), 976 => to_unsigned(669, 10), 977 => to_unsigned(901, 10), 978 => to_unsigned(270, 10), 979 => to_unsigned(626, 10), 980 => to_unsigned(750, 10), 981 => to_unsigned(975, 10), 982 => to_unsigned(819, 10), 983 => to_unsigned(32, 10), 984 => to_unsigned(407, 10), 985 => to_unsigned(761, 10), 986 => to_unsigned(859, 10), 987 => to_unsigned(774, 10), 988 => to_unsigned(713, 10), 989 => to_unsigned(120, 10), 990 => to_unsigned(65, 10), 991 => to_unsigned(75, 10), 992 => to_unsigned(855, 10), 993 => to_unsigned(508, 10), 994 => to_unsigned(710, 10), 995 => to_unsigned(808, 10), 996 => to_unsigned(700, 10), 997 => to_unsigned(36, 10), 998 => to_unsigned(908, 10), 999 => to_unsigned(931, 10), 1000 => to_unsigned(62, 10), 1001 => to_unsigned(453, 10), 1002 => to_unsigned(830, 10), 1003 => to_unsigned(442, 10), 1004 => to_unsigned(588, 10), 1005 => to_unsigned(530, 10), 1006 => to_unsigned(384, 10), 1007 => to_unsigned(1, 10), 1008 => to_unsigned(724, 10), 1009 => to_unsigned(717, 10), 1010 => to_unsigned(602, 10), 1011 => to_unsigned(112, 10), 1012 => to_unsigned(107, 10), 1013 => to_unsigned(149, 10), 1014 => to_unsigned(590, 10), 1015 => to_unsigned(269, 10), 1016 => to_unsigned(1000, 10), 1017 => to_unsigned(67, 10), 1018 => to_unsigned(873, 10), 1019 => to_unsigned(401, 10), 1020 => to_unsigned(261, 10), 1021 => to_unsigned(26, 10), 1022 => to_unsigned(703, 10), 1023 => to_unsigned(411, 10), 1024 => to_unsigned(1003, 10), 1025 => to_unsigned(749, 10), 1026 => to_unsigned(937, 10), 1027 => to_unsigned(525, 10), 1028 => to_unsigned(813, 10), 1029 => to_unsigned(432, 10), 1030 => to_unsigned(568, 10), 1031 => to_unsigned(58, 10), 1032 => to_unsigned(17, 10), 1033 => to_unsigned(214, 10), 1034 => to_unsigned(863, 10), 1035 => to_unsigned(985, 10), 1036 => to_unsigned(220, 10), 1037 => to_unsigned(205, 10), 1038 => to_unsigned(391, 10), 1039 => to_unsigned(282, 10), 1040 => to_unsigned(273, 10), 1041 => to_unsigned(708, 10), 1042 => to_unsigned(555, 10), 1043 => to_unsigned(431, 10), 1044 => to_unsigned(734, 10), 1045 => to_unsigned(125, 10), 1046 => to_unsigned(348, 10), 1047 => to_unsigned(505, 10), 1048 => to_unsigned(840, 10), 1049 => to_unsigned(698, 10), 1050 => to_unsigned(795, 10), 1051 => to_unsigned(6, 10), 1052 => to_unsigned(903, 10), 1053 => to_unsigned(693, 10), 1054 => to_unsigned(887, 10), 1055 => to_unsigned(504, 10), 1056 => to_unsigned(26, 10), 1057 => to_unsigned(635, 10), 1058 => to_unsigned(715, 10), 1059 => to_unsigned(805, 10), 1060 => to_unsigned(93, 10), 1061 => to_unsigned(433, 10), 1062 => to_unsigned(532, 10), 1063 => to_unsigned(477, 10), 1064 => to_unsigned(887, 10), 1065 => to_unsigned(440, 10), 1066 => to_unsigned(957, 10), 1067 => to_unsigned(439, 10), 1068 => to_unsigned(732, 10), 1069 => to_unsigned(151, 10), 1070 => to_unsigned(697, 10), 1071 => to_unsigned(649, 10), 1072 => to_unsigned(640, 10), 1073 => to_unsigned(614, 10), 1074 => to_unsigned(403, 10), 1075 => to_unsigned(455, 10), 1076 => to_unsigned(50, 10), 1077 => to_unsigned(550, 10), 1078 => to_unsigned(963, 10), 1079 => to_unsigned(764, 10), 1080 => to_unsigned(414, 10), 1081 => to_unsigned(549, 10), 1082 => to_unsigned(952, 10), 1083 => to_unsigned(894, 10), 1084 => to_unsigned(1001, 10), 1085 => to_unsigned(645, 10), 1086 => to_unsigned(59, 10), 1087 => to_unsigned(976, 10), 1088 => to_unsigned(474, 10), 1089 => to_unsigned(445, 10), 1090 => to_unsigned(799, 10), 1091 => to_unsigned(966, 10), 1092 => to_unsigned(345, 10), 1093 => to_unsigned(203, 10), 1094 => to_unsigned(657, 10), 1095 => to_unsigned(31, 10), 1096 => to_unsigned(671, 10), 1097 => to_unsigned(84, 10), 1098 => to_unsigned(90, 10), 1099 => to_unsigned(39, 10), 1100 => to_unsigned(757, 10), 1101 => to_unsigned(178, 10), 1102 => to_unsigned(586, 10), 1103 => to_unsigned(294, 10), 1104 => to_unsigned(580, 10), 1105 => to_unsigned(379, 10), 1106 => to_unsigned(551, 10), 1107 => to_unsigned(127, 10), 1108 => to_unsigned(207, 10), 1109 => to_unsigned(13, 10), 1110 => to_unsigned(163, 10), 1111 => to_unsigned(486, 10), 1112 => to_unsigned(891, 10), 1113 => to_unsigned(395, 10), 1114 => to_unsigned(359, 10), 1115 => to_unsigned(331, 10), 1116 => to_unsigned(1008, 10), 1117 => to_unsigned(822, 10), 1118 => to_unsigned(420, 10), 1119 => to_unsigned(82, 10), 1120 => to_unsigned(203, 10), 1121 => to_unsigned(691, 10), 1122 => to_unsigned(162, 10), 1123 => to_unsigned(954, 10), 1124 => to_unsigned(80, 10), 1125 => to_unsigned(540, 10), 1126 => to_unsigned(393, 10), 1127 => to_unsigned(869, 10), 1128 => to_unsigned(8, 10), 1129 => to_unsigned(145, 10), 1130 => to_unsigned(752, 10), 1131 => to_unsigned(236, 10), 1132 => to_unsigned(220, 10), 1133 => to_unsigned(665, 10), 1134 => to_unsigned(350, 10), 1135 => to_unsigned(123, 10), 1136 => to_unsigned(101, 10), 1137 => to_unsigned(699, 10), 1138 => to_unsigned(379, 10), 1139 => to_unsigned(990, 10), 1140 => to_unsigned(1017, 10), 1141 => to_unsigned(59, 10), 1142 => to_unsigned(186, 10), 1143 => to_unsigned(274, 10), 1144 => to_unsigned(524, 10), 1145 => to_unsigned(897, 10), 1146 => to_unsigned(283, 10), 1147 => to_unsigned(522, 10), 1148 => to_unsigned(963, 10), 1149 => to_unsigned(957, 10), 1150 => to_unsigned(784, 10), 1151 => to_unsigned(283, 10), 1152 => to_unsigned(636, 10), 1153 => to_unsigned(774, 10), 1154 => to_unsigned(512, 10), 1155 => to_unsigned(7, 10), 1156 => to_unsigned(665, 10), 1157 => to_unsigned(67, 10), 1158 => to_unsigned(827, 10), 1159 => to_unsigned(760, 10), 1160 => to_unsigned(372, 10), 1161 => to_unsigned(511, 10), 1162 => to_unsigned(420, 10), 1163 => to_unsigned(428, 10), 1164 => to_unsigned(725, 10), 1165 => to_unsigned(625, 10), 1166 => to_unsigned(758, 10), 1167 => to_unsigned(511, 10), 1168 => to_unsigned(200, 10), 1169 => to_unsigned(623, 10), 1170 => to_unsigned(166, 10), 1171 => to_unsigned(938, 10), 1172 => to_unsigned(993, 10), 1173 => to_unsigned(676, 10), 1174 => to_unsigned(68, 10), 1175 => to_unsigned(91, 10), 1176 => to_unsigned(781, 10), 1177 => to_unsigned(653, 10), 1178 => to_unsigned(937, 10), 1179 => to_unsigned(328, 10), 1180 => to_unsigned(646, 10), 1181 => to_unsigned(350, 10), 1182 => to_unsigned(140, 10), 1183 => to_unsigned(610, 10), 1184 => to_unsigned(899, 10), 1185 => to_unsigned(232, 10), 1186 => to_unsigned(528, 10), 1187 => to_unsigned(261, 10), 1188 => to_unsigned(552, 10), 1189 => to_unsigned(439, 10), 1190 => to_unsigned(925, 10), 1191 => to_unsigned(693, 10), 1192 => to_unsigned(278, 10), 1193 => to_unsigned(357, 10), 1194 => to_unsigned(535, 10), 1195 => to_unsigned(251, 10), 1196 => to_unsigned(890, 10), 1197 => to_unsigned(932, 10), 1198 => to_unsigned(747, 10), 1199 => to_unsigned(187, 10), 1200 => to_unsigned(34, 10), 1201 => to_unsigned(966, 10), 1202 => to_unsigned(390, 10), 1203 => to_unsigned(344, 10), 1204 => to_unsigned(588, 10), 1205 => to_unsigned(17, 10), 1206 => to_unsigned(607, 10), 1207 => to_unsigned(560, 10), 1208 => to_unsigned(805, 10), 1209 => to_unsigned(0, 10), 1210 => to_unsigned(458, 10), 1211 => to_unsigned(625, 10), 1212 => to_unsigned(876, 10), 1213 => to_unsigned(4, 10), 1214 => to_unsigned(607, 10), 1215 => to_unsigned(956, 10), 1216 => to_unsigned(639, 10), 1217 => to_unsigned(522, 10), 1218 => to_unsigned(797, 10), 1219 => to_unsigned(865, 10), 1220 => to_unsigned(873, 10), 1221 => to_unsigned(240, 10), 1222 => to_unsigned(525, 10), 1223 => to_unsigned(275, 10), 1224 => to_unsigned(41, 10), 1225 => to_unsigned(204, 10), 1226 => to_unsigned(428, 10), 1227 => to_unsigned(51, 10), 1228 => to_unsigned(107, 10), 1229 => to_unsigned(144, 10), 1230 => to_unsigned(504, 10), 1231 => to_unsigned(1022, 10), 1232 => to_unsigned(754, 10), 1233 => to_unsigned(933, 10), 1234 => to_unsigned(526, 10), 1235 => to_unsigned(676, 10), 1236 => to_unsigned(114, 10), 1237 => to_unsigned(132, 10), 1238 => to_unsigned(1010, 10), 1239 => to_unsigned(303, 10), 1240 => to_unsigned(896, 10), 1241 => to_unsigned(817, 10), 1242 => to_unsigned(933, 10), 1243 => to_unsigned(254, 10), 1244 => to_unsigned(459, 10), 1245 => to_unsigned(812, 10), 1246 => to_unsigned(581, 10), 1247 => to_unsigned(360, 10), 1248 => to_unsigned(494, 10), 1249 => to_unsigned(784, 10), 1250 => to_unsigned(272, 10), 1251 => to_unsigned(778, 10), 1252 => to_unsigned(517, 10), 1253 => to_unsigned(919, 10), 1254 => to_unsigned(943, 10), 1255 => to_unsigned(579, 10), 1256 => to_unsigned(166, 10), 1257 => to_unsigned(1008, 10), 1258 => to_unsigned(274, 10), 1259 => to_unsigned(94, 10), 1260 => to_unsigned(464, 10), 1261 => to_unsigned(799, 10), 1262 => to_unsigned(426, 10), 1263 => to_unsigned(47, 10), 1264 => to_unsigned(277, 10), 1265 => to_unsigned(993, 10), 1266 => to_unsigned(55, 10), 1267 => to_unsigned(330, 10), 1268 => to_unsigned(108, 10), 1269 => to_unsigned(31, 10), 1270 => to_unsigned(595, 10), 1271 => to_unsigned(66, 10), 1272 => to_unsigned(147, 10), 1273 => to_unsigned(159, 10), 1274 => to_unsigned(882, 10), 1275 => to_unsigned(787, 10), 1276 => to_unsigned(807, 10), 1277 => to_unsigned(935, 10), 1278 => to_unsigned(573, 10), 1279 => to_unsigned(609, 10), 1280 => to_unsigned(940, 10), 1281 => to_unsigned(244, 10), 1282 => to_unsigned(748, 10), 1283 => to_unsigned(438, 10), 1284 => to_unsigned(734, 10), 1285 => to_unsigned(122, 10), 1286 => to_unsigned(487, 10), 1287 => to_unsigned(190, 10), 1288 => to_unsigned(204, 10), 1289 => to_unsigned(912, 10), 1290 => to_unsigned(80, 10), 1291 => to_unsigned(510, 10), 1292 => to_unsigned(134, 10), 1293 => to_unsigned(452, 10), 1294 => to_unsigned(813, 10), 1295 => to_unsigned(980, 10), 1296 => to_unsigned(506, 10), 1297 => to_unsigned(670, 10), 1298 => to_unsigned(588, 10), 1299 => to_unsigned(891, 10), 1300 => to_unsigned(693, 10), 1301 => to_unsigned(417, 10), 1302 => to_unsigned(602, 10), 1303 => to_unsigned(402, 10), 1304 => to_unsigned(134, 10), 1305 => to_unsigned(632, 10), 1306 => to_unsigned(130, 10), 1307 => to_unsigned(154, 10), 1308 => to_unsigned(238, 10), 1309 => to_unsigned(281, 10), 1310 => to_unsigned(525, 10), 1311 => to_unsigned(959, 10), 1312 => to_unsigned(731, 10), 1313 => to_unsigned(574, 10), 1314 => to_unsigned(57, 10), 1315 => to_unsigned(293, 10), 1316 => to_unsigned(941, 10), 1317 => to_unsigned(405, 10), 1318 => to_unsigned(107, 10), 1319 => to_unsigned(504, 10), 1320 => to_unsigned(837, 10), 1321 => to_unsigned(1017, 10), 1322 => to_unsigned(817, 10), 1323 => to_unsigned(25, 10), 1324 => to_unsigned(268, 10), 1325 => to_unsigned(564, 10), 1326 => to_unsigned(838, 10), 1327 => to_unsigned(943, 10), 1328 => to_unsigned(765, 10), 1329 => to_unsigned(73, 10), 1330 => to_unsigned(906, 10), 1331 => to_unsigned(584, 10), 1332 => to_unsigned(474, 10), 1333 => to_unsigned(144, 10), 1334 => to_unsigned(351, 10), 1335 => to_unsigned(862, 10), 1336 => to_unsigned(766, 10), 1337 => to_unsigned(229, 10), 1338 => to_unsigned(294, 10), 1339 => to_unsigned(176, 10), 1340 => to_unsigned(700, 10), 1341 => to_unsigned(518, 10), 1342 => to_unsigned(1008, 10), 1343 => to_unsigned(966, 10), 1344 => to_unsigned(631, 10), 1345 => to_unsigned(513, 10), 1346 => to_unsigned(367, 10), 1347 => to_unsigned(191, 10), 1348 => to_unsigned(193, 10), 1349 => to_unsigned(637, 10), 1350 => to_unsigned(277, 10), 1351 => to_unsigned(814, 10), 1352 => to_unsigned(768, 10), 1353 => to_unsigned(726, 10), 1354 => to_unsigned(164, 10), 1355 => to_unsigned(666, 10), 1356 => to_unsigned(660, 10), 1357 => to_unsigned(340, 10), 1358 => to_unsigned(231, 10), 1359 => to_unsigned(546, 10), 1360 => to_unsigned(241, 10), 1361 => to_unsigned(878, 10), 1362 => to_unsigned(61, 10), 1363 => to_unsigned(926, 10), 1364 => to_unsigned(667, 10), 1365 => to_unsigned(740, 10), 1366 => to_unsigned(585, 10), 1367 => to_unsigned(328, 10), 1368 => to_unsigned(564, 10), 1369 => to_unsigned(596, 10), 1370 => to_unsigned(919, 10), 1371 => to_unsigned(318, 10), 1372 => to_unsigned(48, 10), 1373 => to_unsigned(999, 10), 1374 => to_unsigned(443, 10), 1375 => to_unsigned(299, 10), 1376 => to_unsigned(938, 10), 1377 => to_unsigned(653, 10), 1378 => to_unsigned(504, 10), 1379 => to_unsigned(367, 10), 1380 => to_unsigned(1017, 10), 1381 => to_unsigned(777, 10), 1382 => to_unsigned(155, 10), 1383 => to_unsigned(602, 10), 1384 => to_unsigned(997, 10), 1385 => to_unsigned(546, 10), 1386 => to_unsigned(838, 10), 1387 => to_unsigned(425, 10), 1388 => to_unsigned(1005, 10), 1389 => to_unsigned(37, 10), 1390 => to_unsigned(6, 10), 1391 => to_unsigned(314, 10), 1392 => to_unsigned(597, 10), 1393 => to_unsigned(3, 10), 1394 => to_unsigned(75, 10), 1395 => to_unsigned(746, 10), 1396 => to_unsigned(267, 10), 1397 => to_unsigned(413, 10), 1398 => to_unsigned(78, 10), 1399 => to_unsigned(723, 10), 1400 => to_unsigned(282, 10), 1401 => to_unsigned(363, 10), 1402 => to_unsigned(767, 10), 1403 => to_unsigned(80, 10), 1404 => to_unsigned(163, 10), 1405 => to_unsigned(564, 10), 1406 => to_unsigned(913, 10), 1407 => to_unsigned(592, 10), 1408 => to_unsigned(394, 10), 1409 => to_unsigned(1017, 10), 1410 => to_unsigned(188, 10), 1411 => to_unsigned(969, 10), 1412 => to_unsigned(99, 10), 1413 => to_unsigned(921, 10), 1414 => to_unsigned(639, 10), 1415 => to_unsigned(154, 10), 1416 => to_unsigned(563, 10), 1417 => to_unsigned(335, 10), 1418 => to_unsigned(283, 10), 1419 => to_unsigned(132, 10), 1420 => to_unsigned(358, 10), 1421 => to_unsigned(725, 10), 1422 => to_unsigned(103, 10), 1423 => to_unsigned(241, 10), 1424 => to_unsigned(437, 10), 1425 => to_unsigned(791, 10), 1426 => to_unsigned(1004, 10), 1427 => to_unsigned(998, 10), 1428 => to_unsigned(363, 10), 1429 => to_unsigned(619, 10), 1430 => to_unsigned(534, 10), 1431 => to_unsigned(348, 10), 1432 => to_unsigned(1006, 10), 1433 => to_unsigned(43, 10), 1434 => to_unsigned(6, 10), 1435 => to_unsigned(909, 10), 1436 => to_unsigned(205, 10), 1437 => to_unsigned(145, 10), 1438 => to_unsigned(424, 10), 1439 => to_unsigned(637, 10), 1440 => to_unsigned(478, 10), 1441 => to_unsigned(452, 10), 1442 => to_unsigned(786, 10), 1443 => to_unsigned(752, 10), 1444 => to_unsigned(130, 10), 1445 => to_unsigned(27, 10), 1446 => to_unsigned(392, 10), 1447 => to_unsigned(747, 10), 1448 => to_unsigned(207, 10), 1449 => to_unsigned(563, 10), 1450 => to_unsigned(215, 10), 1451 => to_unsigned(943, 10), 1452 => to_unsigned(831, 10), 1453 => to_unsigned(158, 10), 1454 => to_unsigned(525, 10), 1455 => to_unsigned(860, 10), 1456 => to_unsigned(942, 10), 1457 => to_unsigned(910, 10), 1458 => to_unsigned(754, 10), 1459 => to_unsigned(174, 10), 1460 => to_unsigned(173, 10), 1461 => to_unsigned(609, 10), 1462 => to_unsigned(260, 10), 1463 => to_unsigned(884, 10), 1464 => to_unsigned(650, 10), 1465 => to_unsigned(372, 10), 1466 => to_unsigned(63, 10), 1467 => to_unsigned(274, 10), 1468 => to_unsigned(484, 10), 1469 => to_unsigned(200, 10), 1470 => to_unsigned(119, 10), 1471 => to_unsigned(314, 10), 1472 => to_unsigned(713, 10), 1473 => to_unsigned(750, 10), 1474 => to_unsigned(397, 10), 1475 => to_unsigned(524, 10), 1476 => to_unsigned(669, 10), 1477 => to_unsigned(590, 10), 1478 => to_unsigned(360, 10), 1479 => to_unsigned(77, 10), 1480 => to_unsigned(649, 10), 1481 => to_unsigned(942, 10), 1482 => to_unsigned(700, 10), 1483 => to_unsigned(588, 10), 1484 => to_unsigned(229, 10), 1485 => to_unsigned(669, 10), 1486 => to_unsigned(109, 10), 1487 => to_unsigned(75, 10), 1488 => to_unsigned(492, 10), 1489 => to_unsigned(1001, 10), 1490 => to_unsigned(881, 10), 1491 => to_unsigned(920, 10), 1492 => to_unsigned(827, 10), 1493 => to_unsigned(968, 10), 1494 => to_unsigned(655, 10), 1495 => to_unsigned(438, 10), 1496 => to_unsigned(672, 10), 1497 => to_unsigned(492, 10), 1498 => to_unsigned(254, 10), 1499 => to_unsigned(720, 10), 1500 => to_unsigned(1010, 10), 1501 => to_unsigned(371, 10), 1502 => to_unsigned(620, 10), 1503 => to_unsigned(114, 10), 1504 => to_unsigned(369, 10), 1505 => to_unsigned(11, 10), 1506 => to_unsigned(271, 10), 1507 => to_unsigned(281, 10), 1508 => to_unsigned(789, 10), 1509 => to_unsigned(150, 10), 1510 => to_unsigned(977, 10), 1511 => to_unsigned(988, 10), 1512 => to_unsigned(762, 10), 1513 => to_unsigned(859, 10), 1514 => to_unsigned(108, 10), 1515 => to_unsigned(456, 10), 1516 => to_unsigned(859, 10), 1517 => to_unsigned(476, 10), 1518 => to_unsigned(743, 10), 1519 => to_unsigned(619, 10), 1520 => to_unsigned(103, 10), 1521 => to_unsigned(99, 10), 1522 => to_unsigned(414, 10), 1523 => to_unsigned(756, 10), 1524 => to_unsigned(937, 10), 1525 => to_unsigned(758, 10), 1526 => to_unsigned(393, 10), 1527 => to_unsigned(886, 10), 1528 => to_unsigned(820, 10), 1529 => to_unsigned(299, 10), 1530 => to_unsigned(849, 10), 1531 => to_unsigned(946, 10), 1532 => to_unsigned(400, 10), 1533 => to_unsigned(64, 10), 1534 => to_unsigned(794, 10), 1535 => to_unsigned(135, 10), 1536 => to_unsigned(438, 10), 1537 => to_unsigned(850, 10), 1538 => to_unsigned(954, 10), 1539 => to_unsigned(331, 10), 1540 => to_unsigned(313, 10), 1541 => to_unsigned(698, 10), 1542 => to_unsigned(972, 10), 1543 => to_unsigned(269, 10), 1544 => to_unsigned(968, 10), 1545 => to_unsigned(232, 10), 1546 => to_unsigned(786, 10), 1547 => to_unsigned(145, 10), 1548 => to_unsigned(170, 10), 1549 => to_unsigned(300, 10), 1550 => to_unsigned(226, 10), 1551 => to_unsigned(715, 10), 1552 => to_unsigned(855, 10), 1553 => to_unsigned(838, 10), 1554 => to_unsigned(206, 10), 1555 => to_unsigned(558, 10), 1556 => to_unsigned(566, 10), 1557 => to_unsigned(690, 10), 1558 => to_unsigned(43, 10), 1559 => to_unsigned(577, 10), 1560 => to_unsigned(974, 10), 1561 => to_unsigned(357, 10), 1562 => to_unsigned(262, 10), 1563 => to_unsigned(121, 10), 1564 => to_unsigned(175, 10), 1565 => to_unsigned(172, 10), 1566 => to_unsigned(777, 10), 1567 => to_unsigned(515, 10), 1568 => to_unsigned(393, 10), 1569 => to_unsigned(123, 10), 1570 => to_unsigned(756, 10), 1571 => to_unsigned(507, 10), 1572 => to_unsigned(34, 10), 1573 => to_unsigned(478, 10), 1574 => to_unsigned(513, 10), 1575 => to_unsigned(294, 10), 1576 => to_unsigned(206, 10), 1577 => to_unsigned(976, 10), 1578 => to_unsigned(862, 10), 1579 => to_unsigned(434, 10), 1580 => to_unsigned(141, 10), 1581 => to_unsigned(854, 10), 1582 => to_unsigned(46, 10), 1583 => to_unsigned(995, 10), 1584 => to_unsigned(855, 10), 1585 => to_unsigned(805, 10), 1586 => to_unsigned(861, 10), 1587 => to_unsigned(749, 10), 1588 => to_unsigned(746, 10), 1589 => to_unsigned(346, 10), 1590 => to_unsigned(82, 10), 1591 => to_unsigned(982, 10), 1592 => to_unsigned(518, 10), 1593 => to_unsigned(586, 10), 1594 => to_unsigned(427, 10), 1595 => to_unsigned(513, 10), 1596 => to_unsigned(457, 10), 1597 => to_unsigned(474, 10), 1598 => to_unsigned(176, 10), 1599 => to_unsigned(847, 10), 1600 => to_unsigned(401, 10), 1601 => to_unsigned(275, 10), 1602 => to_unsigned(254, 10), 1603 => to_unsigned(147, 10), 1604 => to_unsigned(833, 10), 1605 => to_unsigned(411, 10), 1606 => to_unsigned(1011, 10), 1607 => to_unsigned(740, 10), 1608 => to_unsigned(931, 10), 1609 => to_unsigned(265, 10), 1610 => to_unsigned(745, 10), 1611 => to_unsigned(13, 10), 1612 => to_unsigned(437, 10), 1613 => to_unsigned(326, 10), 1614 => to_unsigned(984, 10), 1615 => to_unsigned(778, 10), 1616 => to_unsigned(121, 10), 1617 => to_unsigned(299, 10), 1618 => to_unsigned(613, 10), 1619 => to_unsigned(389, 10), 1620 => to_unsigned(168, 10), 1621 => to_unsigned(244, 10), 1622 => to_unsigned(783, 10), 1623 => to_unsigned(14, 10), 1624 => to_unsigned(469, 10), 1625 => to_unsigned(0, 10), 1626 => to_unsigned(291, 10), 1627 => to_unsigned(609, 10), 1628 => to_unsigned(398, 10), 1629 => to_unsigned(774, 10), 1630 => to_unsigned(600, 10), 1631 => to_unsigned(502, 10), 1632 => to_unsigned(3, 10), 1633 => to_unsigned(324, 10), 1634 => to_unsigned(101, 10), 1635 => to_unsigned(488, 10), 1636 => to_unsigned(863, 10), 1637 => to_unsigned(923, 10), 1638 => to_unsigned(626, 10), 1639 => to_unsigned(1001, 10), 1640 => to_unsigned(579, 10), 1641 => to_unsigned(802, 10), 1642 => to_unsigned(425, 10), 1643 => to_unsigned(781, 10), 1644 => to_unsigned(895, 10), 1645 => to_unsigned(113, 10), 1646 => to_unsigned(401, 10), 1647 => to_unsigned(362, 10), 1648 => to_unsigned(680, 10), 1649 => to_unsigned(493, 10), 1650 => to_unsigned(970, 10), 1651 => to_unsigned(806, 10), 1652 => to_unsigned(554, 10), 1653 => to_unsigned(323, 10), 1654 => to_unsigned(283, 10), 1655 => to_unsigned(956, 10), 1656 => to_unsigned(655, 10), 1657 => to_unsigned(754, 10), 1658 => to_unsigned(930, 10), 1659 => to_unsigned(484, 10), 1660 => to_unsigned(746, 10), 1661 => to_unsigned(615, 10), 1662 => to_unsigned(690, 10), 1663 => to_unsigned(44, 10), 1664 => to_unsigned(340, 10), 1665 => to_unsigned(564, 10), 1666 => to_unsigned(921, 10), 1667 => to_unsigned(715, 10), 1668 => to_unsigned(172, 10), 1669 => to_unsigned(81, 10), 1670 => to_unsigned(1023, 10), 1671 => to_unsigned(645, 10), 1672 => to_unsigned(595, 10), 1673 => to_unsigned(711, 10), 1674 => to_unsigned(255, 10), 1675 => to_unsigned(836, 10), 1676 => to_unsigned(607, 10), 1677 => to_unsigned(349, 10), 1678 => to_unsigned(106, 10), 1679 => to_unsigned(754, 10), 1680 => to_unsigned(603, 10), 1681 => to_unsigned(160, 10), 1682 => to_unsigned(491, 10), 1683 => to_unsigned(937, 10), 1684 => to_unsigned(210, 10), 1685 => to_unsigned(413, 10), 1686 => to_unsigned(909, 10), 1687 => to_unsigned(1010, 10), 1688 => to_unsigned(364, 10), 1689 => to_unsigned(649, 10), 1690 => to_unsigned(54, 10), 1691 => to_unsigned(904, 10), 1692 => to_unsigned(25, 10), 1693 => to_unsigned(161, 10), 1694 => to_unsigned(529, 10), 1695 => to_unsigned(497, 10), 1696 => to_unsigned(431, 10), 1697 => to_unsigned(528, 10), 1698 => to_unsigned(561, 10), 1699 => to_unsigned(62, 10), 1700 => to_unsigned(839, 10), 1701 => to_unsigned(862, 10), 1702 => to_unsigned(1022, 10), 1703 => to_unsigned(976, 10), 1704 => to_unsigned(86, 10), 1705 => to_unsigned(507, 10), 1706 => to_unsigned(165, 10), 1707 => to_unsigned(265, 10), 1708 => to_unsigned(942, 10), 1709 => to_unsigned(652, 10), 1710 => to_unsigned(88, 10), 1711 => to_unsigned(381, 10), 1712 => to_unsigned(373, 10), 1713 => to_unsigned(406, 10), 1714 => to_unsigned(184, 10), 1715 => to_unsigned(590, 10), 1716 => to_unsigned(557, 10), 1717 => to_unsigned(801, 10), 1718 => to_unsigned(702, 10), 1719 => to_unsigned(516, 10), 1720 => to_unsigned(837, 10), 1721 => to_unsigned(637, 10), 1722 => to_unsigned(76, 10), 1723 => to_unsigned(681, 10), 1724 => to_unsigned(396, 10), 1725 => to_unsigned(768, 10), 1726 => to_unsigned(709, 10), 1727 => to_unsigned(150, 10), 1728 => to_unsigned(745, 10), 1729 => to_unsigned(353, 10), 1730 => to_unsigned(689, 10), 1731 => to_unsigned(627, 10), 1732 => to_unsigned(833, 10), 1733 => to_unsigned(394, 10), 1734 => to_unsigned(198, 10), 1735 => to_unsigned(122, 10), 1736 => to_unsigned(16, 10), 1737 => to_unsigned(711, 10), 1738 => to_unsigned(411, 10), 1739 => to_unsigned(294, 10), 1740 => to_unsigned(107, 10), 1741 => to_unsigned(84, 10), 1742 => to_unsigned(425, 10), 1743 => to_unsigned(722, 10), 1744 => to_unsigned(627, 10), 1745 => to_unsigned(1002, 10), 1746 => to_unsigned(454, 10), 1747 => to_unsigned(934, 10), 1748 => to_unsigned(674, 10), 1749 => to_unsigned(113, 10), 1750 => to_unsigned(714, 10), 1751 => to_unsigned(767, 10), 1752 => to_unsigned(359, 10), 1753 => to_unsigned(808, 10), 1754 => to_unsigned(40, 10), 1755 => to_unsigned(923, 10), 1756 => to_unsigned(94, 10), 1757 => to_unsigned(1019, 10), 1758 => to_unsigned(164, 10), 1759 => to_unsigned(98, 10), 1760 => to_unsigned(571, 10), 1761 => to_unsigned(601, 10), 1762 => to_unsigned(923, 10), 1763 => to_unsigned(696, 10), 1764 => to_unsigned(127, 10), 1765 => to_unsigned(954, 10), 1766 => to_unsigned(287, 10), 1767 => to_unsigned(816, 10), 1768 => to_unsigned(1003, 10), 1769 => to_unsigned(126, 10), 1770 => to_unsigned(387, 10), 1771 => to_unsigned(320, 10), 1772 => to_unsigned(549, 10), 1773 => to_unsigned(503, 10), 1774 => to_unsigned(679, 10), 1775 => to_unsigned(12, 10), 1776 => to_unsigned(852, 10), 1777 => to_unsigned(459, 10), 1778 => to_unsigned(332, 10), 1779 => to_unsigned(632, 10), 1780 => to_unsigned(370, 10), 1781 => to_unsigned(987, 10), 1782 => to_unsigned(943, 10), 1783 => to_unsigned(313, 10), 1784 => to_unsigned(149, 10), 1785 => to_unsigned(876, 10), 1786 => to_unsigned(524, 10), 1787 => to_unsigned(1007, 10), 1788 => to_unsigned(657, 10), 1789 => to_unsigned(423, 10), 1790 => to_unsigned(927, 10), 1791 => to_unsigned(623, 10), 1792 => to_unsigned(669, 10), 1793 => to_unsigned(439, 10), 1794 => to_unsigned(449, 10), 1795 => to_unsigned(293, 10), 1796 => to_unsigned(512, 10), 1797 => to_unsigned(791, 10), 1798 => to_unsigned(909, 10), 1799 => to_unsigned(136, 10), 1800 => to_unsigned(468, 10), 1801 => to_unsigned(53, 10), 1802 => to_unsigned(210, 10), 1803 => to_unsigned(336, 10), 1804 => to_unsigned(781, 10), 1805 => to_unsigned(392, 10), 1806 => to_unsigned(390, 10), 1807 => to_unsigned(411, 10), 1808 => to_unsigned(165, 10), 1809 => to_unsigned(419, 10), 1810 => to_unsigned(552, 10), 1811 => to_unsigned(666, 10), 1812 => to_unsigned(350, 10), 1813 => to_unsigned(972, 10), 1814 => to_unsigned(441, 10), 1815 => to_unsigned(301, 10), 1816 => to_unsigned(848, 10), 1817 => to_unsigned(314, 10), 1818 => to_unsigned(151, 10), 1819 => to_unsigned(766, 10), 1820 => to_unsigned(242, 10), 1821 => to_unsigned(746, 10), 1822 => to_unsigned(968, 10), 1823 => to_unsigned(1015, 10), 1824 => to_unsigned(1014, 10), 1825 => to_unsigned(464, 10), 1826 => to_unsigned(245, 10), 1827 => to_unsigned(893, 10), 1828 => to_unsigned(530, 10), 1829 => to_unsigned(970, 10), 1830 => to_unsigned(911, 10), 1831 => to_unsigned(486, 10), 1832 => to_unsigned(893, 10), 1833 => to_unsigned(856, 10), 1834 => to_unsigned(996, 10), 1835 => to_unsigned(751, 10), 1836 => to_unsigned(832, 10), 1837 => to_unsigned(387, 10), 1838 => to_unsigned(986, 10), 1839 => to_unsigned(916, 10), 1840 => to_unsigned(1007, 10), 1841 => to_unsigned(175, 10), 1842 => to_unsigned(446, 10), 1843 => to_unsigned(353, 10), 1844 => to_unsigned(24, 10), 1845 => to_unsigned(722, 10), 1846 => to_unsigned(808, 10), 1847 => to_unsigned(137, 10), 1848 => to_unsigned(328, 10), 1849 => to_unsigned(199, 10), 1850 => to_unsigned(476, 10), 1851 => to_unsigned(1007, 10), 1852 => to_unsigned(297, 10), 1853 => to_unsigned(787, 10), 1854 => to_unsigned(726, 10), 1855 => to_unsigned(323, 10), 1856 => to_unsigned(1015, 10), 1857 => to_unsigned(974, 10), 1858 => to_unsigned(127, 10), 1859 => to_unsigned(631, 10), 1860 => to_unsigned(834, 10), 1861 => to_unsigned(727, 10), 1862 => to_unsigned(235, 10), 1863 => to_unsigned(24, 10), 1864 => to_unsigned(596, 10), 1865 => to_unsigned(675, 10), 1866 => to_unsigned(890, 10), 1867 => to_unsigned(430, 10), 1868 => to_unsigned(544, 10), 1869 => to_unsigned(802, 10), 1870 => to_unsigned(554, 10), 1871 => to_unsigned(860, 10), 1872 => to_unsigned(37, 10), 1873 => to_unsigned(228, 10), 1874 => to_unsigned(850, 10), 1875 => to_unsigned(55, 10), 1876 => to_unsigned(874, 10), 1877 => to_unsigned(547, 10), 1878 => to_unsigned(999, 10), 1879 => to_unsigned(355, 10), 1880 => to_unsigned(65, 10), 1881 => to_unsigned(349, 10), 1882 => to_unsigned(660, 10), 1883 => to_unsigned(229, 10), 1884 => to_unsigned(355, 10), 1885 => to_unsigned(814, 10), 1886 => to_unsigned(354, 10), 1887 => to_unsigned(91, 10), 1888 => to_unsigned(62, 10), 1889 => to_unsigned(62, 10), 1890 => to_unsigned(497, 10), 1891 => to_unsigned(251, 10), 1892 => to_unsigned(590, 10), 1893 => to_unsigned(874, 10), 1894 => to_unsigned(158, 10), 1895 => to_unsigned(347, 10), 1896 => to_unsigned(51, 10), 1897 => to_unsigned(516, 10), 1898 => to_unsigned(708, 10), 1899 => to_unsigned(902, 10), 1900 => to_unsigned(745, 10), 1901 => to_unsigned(809, 10), 1902 => to_unsigned(259, 10), 1903 => to_unsigned(679, 10), 1904 => to_unsigned(492, 10), 1905 => to_unsigned(100, 10), 1906 => to_unsigned(411, 10), 1907 => to_unsigned(653, 10), 1908 => to_unsigned(300, 10), 1909 => to_unsigned(256, 10), 1910 => to_unsigned(842, 10), 1911 => to_unsigned(733, 10), 1912 => to_unsigned(846, 10), 1913 => to_unsigned(128, 10), 1914 => to_unsigned(256, 10), 1915 => to_unsigned(96, 10), 1916 => to_unsigned(884, 10), 1917 => to_unsigned(779, 10), 1918 => to_unsigned(29, 10), 1919 => to_unsigned(389, 10), 1920 => to_unsigned(69, 10), 1921 => to_unsigned(697, 10), 1922 => to_unsigned(286, 10), 1923 => to_unsigned(786, 10), 1924 => to_unsigned(618, 10), 1925 => to_unsigned(16, 10), 1926 => to_unsigned(887, 10), 1927 => to_unsigned(337, 10), 1928 => to_unsigned(203, 10), 1929 => to_unsigned(9, 10), 1930 => to_unsigned(905, 10), 1931 => to_unsigned(730, 10), 1932 => to_unsigned(76, 10), 1933 => to_unsigned(704, 10), 1934 => to_unsigned(231, 10), 1935 => to_unsigned(924, 10), 1936 => to_unsigned(758, 10), 1937 => to_unsigned(845, 10), 1938 => to_unsigned(855, 10), 1939 => to_unsigned(954, 10), 1940 => to_unsigned(633, 10), 1941 => to_unsigned(432, 10), 1942 => to_unsigned(411, 10), 1943 => to_unsigned(875, 10), 1944 => to_unsigned(153, 10), 1945 => to_unsigned(980, 10), 1946 => to_unsigned(111, 10), 1947 => to_unsigned(588, 10), 1948 => to_unsigned(536, 10), 1949 => to_unsigned(773, 10), 1950 => to_unsigned(34, 10), 1951 => to_unsigned(76, 10), 1952 => to_unsigned(187, 10), 1953 => to_unsigned(555, 10), 1954 => to_unsigned(975, 10), 1955 => to_unsigned(827, 10), 1956 => to_unsigned(277, 10), 1957 => to_unsigned(484, 10), 1958 => to_unsigned(497, 10), 1959 => to_unsigned(510, 10), 1960 => to_unsigned(364, 10), 1961 => to_unsigned(524, 10), 1962 => to_unsigned(880, 10), 1963 => to_unsigned(98, 10), 1964 => to_unsigned(645, 10), 1965 => to_unsigned(788, 10), 1966 => to_unsigned(636, 10), 1967 => to_unsigned(671, 10), 1968 => to_unsigned(866, 10), 1969 => to_unsigned(279, 10), 1970 => to_unsigned(531, 10), 1971 => to_unsigned(597, 10), 1972 => to_unsigned(815, 10), 1973 => to_unsigned(1018, 10), 1974 => to_unsigned(774, 10), 1975 => to_unsigned(68, 10), 1976 => to_unsigned(201, 10), 1977 => to_unsigned(536, 10), 1978 => to_unsigned(943, 10), 1979 => to_unsigned(928, 10), 1980 => to_unsigned(970, 10), 1981 => to_unsigned(730, 10), 1982 => to_unsigned(475, 10), 1983 => to_unsigned(272, 10), 1984 => to_unsigned(738, 10), 1985 => to_unsigned(150, 10), 1986 => to_unsigned(125, 10), 1987 => to_unsigned(28, 10), 1988 => to_unsigned(284, 10), 1989 => to_unsigned(625, 10), 1990 => to_unsigned(974, 10), 1991 => to_unsigned(869, 10), 1992 => to_unsigned(601, 10), 1993 => to_unsigned(133, 10), 1994 => to_unsigned(578, 10), 1995 => to_unsigned(419, 10), 1996 => to_unsigned(715, 10), 1997 => to_unsigned(947, 10), 1998 => to_unsigned(589, 10), 1999 => to_unsigned(995, 10), 2000 => to_unsigned(696, 10), 2001 => to_unsigned(479, 10), 2002 => to_unsigned(478, 10), 2003 => to_unsigned(261, 10), 2004 => to_unsigned(29, 10), 2005 => to_unsigned(91, 10), 2006 => to_unsigned(1017, 10), 2007 => to_unsigned(949, 10), 2008 => to_unsigned(449, 10), 2009 => to_unsigned(317, 10), 2010 => to_unsigned(488, 10), 2011 => to_unsigned(154, 10), 2012 => to_unsigned(284, 10), 2013 => to_unsigned(999, 10), 2014 => to_unsigned(423, 10), 2015 => to_unsigned(609, 10), 2016 => to_unsigned(105, 10), 2017 => to_unsigned(687, 10), 2018 => to_unsigned(109, 10), 2019 => to_unsigned(928, 10), 2020 => to_unsigned(377, 10), 2021 => to_unsigned(260, 10), 2022 => to_unsigned(438, 10), 2023 => to_unsigned(384, 10), 2024 => to_unsigned(267, 10), 2025 => to_unsigned(179, 10), 2026 => to_unsigned(611, 10), 2027 => to_unsigned(964, 10), 2028 => to_unsigned(794, 10), 2029 => to_unsigned(527, 10), 2030 => to_unsigned(497, 10), 2031 => to_unsigned(732, 10), 2032 => to_unsigned(874, 10), 2033 => to_unsigned(912, 10), 2034 => to_unsigned(884, 10), 2035 => to_unsigned(70, 10), 2036 => to_unsigned(760, 10), 2037 => to_unsigned(95, 10), 2038 => to_unsigned(2, 10), 2039 => to_unsigned(508, 10), 2040 => to_unsigned(273, 10), 2041 => to_unsigned(242, 10), 2042 => to_unsigned(833, 10), 2043 => to_unsigned(160, 10), 2044 => to_unsigned(225, 10), 2045 => to_unsigned(422, 10), 2046 => to_unsigned(580, 10), 2047 => to_unsigned(862, 10)),
            2 => (0 => to_unsigned(260, 10), 1 => to_unsigned(1019, 10), 2 => to_unsigned(335, 10), 3 => to_unsigned(127, 10), 4 => to_unsigned(277, 10), 5 => to_unsigned(889, 10), 6 => to_unsigned(371, 10), 7 => to_unsigned(102, 10), 8 => to_unsigned(778, 10), 9 => to_unsigned(272, 10), 10 => to_unsigned(2, 10), 11 => to_unsigned(814, 10), 12 => to_unsigned(701, 10), 13 => to_unsigned(174, 10), 14 => to_unsigned(110, 10), 15 => to_unsigned(288, 10), 16 => to_unsigned(231, 10), 17 => to_unsigned(919, 10), 18 => to_unsigned(701, 10), 19 => to_unsigned(385, 10), 20 => to_unsigned(292, 10), 21 => to_unsigned(857, 10), 22 => to_unsigned(264, 10), 23 => to_unsigned(559, 10), 24 => to_unsigned(859, 10), 25 => to_unsigned(0, 10), 26 => to_unsigned(163, 10), 27 => to_unsigned(26, 10), 28 => to_unsigned(190, 10), 29 => to_unsigned(879, 10), 30 => to_unsigned(948, 10), 31 => to_unsigned(1002, 10), 32 => to_unsigned(662, 10), 33 => to_unsigned(671, 10), 34 => to_unsigned(641, 10), 35 => to_unsigned(861, 10), 36 => to_unsigned(259, 10), 37 => to_unsigned(259, 10), 38 => to_unsigned(354, 10), 39 => to_unsigned(116, 10), 40 => to_unsigned(164, 10), 41 => to_unsigned(426, 10), 42 => to_unsigned(366, 10), 43 => to_unsigned(20, 10), 44 => to_unsigned(233, 10), 45 => to_unsigned(133, 10), 46 => to_unsigned(728, 10), 47 => to_unsigned(1023, 10), 48 => to_unsigned(83, 10), 49 => to_unsigned(694, 10), 50 => to_unsigned(741, 10), 51 => to_unsigned(259, 10), 52 => to_unsigned(851, 10), 53 => to_unsigned(151, 10), 54 => to_unsigned(48, 10), 55 => to_unsigned(862, 10), 56 => to_unsigned(670, 10), 57 => to_unsigned(217, 10), 58 => to_unsigned(903, 10), 59 => to_unsigned(938, 10), 60 => to_unsigned(652, 10), 61 => to_unsigned(516, 10), 62 => to_unsigned(240, 10), 63 => to_unsigned(923, 10), 64 => to_unsigned(204, 10), 65 => to_unsigned(623, 10), 66 => to_unsigned(714, 10), 67 => to_unsigned(764, 10), 68 => to_unsigned(427, 10), 69 => to_unsigned(693, 10), 70 => to_unsigned(238, 10), 71 => to_unsigned(650, 10), 72 => to_unsigned(755, 10), 73 => to_unsigned(43, 10), 74 => to_unsigned(774, 10), 75 => to_unsigned(711, 10), 76 => to_unsigned(512, 10), 77 => to_unsigned(563, 10), 78 => to_unsigned(674, 10), 79 => to_unsigned(864, 10), 80 => to_unsigned(23, 10), 81 => to_unsigned(448, 10), 82 => to_unsigned(711, 10), 83 => to_unsigned(926, 10), 84 => to_unsigned(786, 10), 85 => to_unsigned(800, 10), 86 => to_unsigned(2, 10), 87 => to_unsigned(678, 10), 88 => to_unsigned(268, 10), 89 => to_unsigned(576, 10), 90 => to_unsigned(894, 10), 91 => to_unsigned(764, 10), 92 => to_unsigned(72, 10), 93 => to_unsigned(771, 10), 94 => to_unsigned(397, 10), 95 => to_unsigned(894, 10), 96 => to_unsigned(986, 10), 97 => to_unsigned(131, 10), 98 => to_unsigned(230, 10), 99 => to_unsigned(454, 10), 100 => to_unsigned(646, 10), 101 => to_unsigned(404, 10), 102 => to_unsigned(826, 10), 103 => to_unsigned(2, 10), 104 => to_unsigned(981, 10), 105 => to_unsigned(175, 10), 106 => to_unsigned(511, 10), 107 => to_unsigned(692, 10), 108 => to_unsigned(570, 10), 109 => to_unsigned(110, 10), 110 => to_unsigned(594, 10), 111 => to_unsigned(254, 10), 112 => to_unsigned(592, 10), 113 => to_unsigned(313, 10), 114 => to_unsigned(683, 10), 115 => to_unsigned(289, 10), 116 => to_unsigned(490, 10), 117 => to_unsigned(69, 10), 118 => to_unsigned(221, 10), 119 => to_unsigned(79, 10), 120 => to_unsigned(89, 10), 121 => to_unsigned(493, 10), 122 => to_unsigned(1013, 10), 123 => to_unsigned(280, 10), 124 => to_unsigned(356, 10), 125 => to_unsigned(700, 10), 126 => to_unsigned(889, 10), 127 => to_unsigned(832, 10), 128 => to_unsigned(445, 10), 129 => to_unsigned(77, 10), 130 => to_unsigned(524, 10), 131 => to_unsigned(710, 10), 132 => to_unsigned(113, 10), 133 => to_unsigned(561, 10), 134 => to_unsigned(131, 10), 135 => to_unsigned(928, 10), 136 => to_unsigned(115, 10), 137 => to_unsigned(689, 10), 138 => to_unsigned(739, 10), 139 => to_unsigned(397, 10), 140 => to_unsigned(75, 10), 141 => to_unsigned(17, 10), 142 => to_unsigned(68, 10), 143 => to_unsigned(471, 10), 144 => to_unsigned(303, 10), 145 => to_unsigned(330, 10), 146 => to_unsigned(422, 10), 147 => to_unsigned(628, 10), 148 => to_unsigned(245, 10), 149 => to_unsigned(870, 10), 150 => to_unsigned(432, 10), 151 => to_unsigned(548, 10), 152 => to_unsigned(477, 10), 153 => to_unsigned(793, 10), 154 => to_unsigned(547, 10), 155 => to_unsigned(455, 10), 156 => to_unsigned(960, 10), 157 => to_unsigned(832, 10), 158 => to_unsigned(8, 10), 159 => to_unsigned(963, 10), 160 => to_unsigned(774, 10), 161 => to_unsigned(101, 10), 162 => to_unsigned(1020, 10), 163 => to_unsigned(391, 10), 164 => to_unsigned(947, 10), 165 => to_unsigned(461, 10), 166 => to_unsigned(82, 10), 167 => to_unsigned(376, 10), 168 => to_unsigned(529, 10), 169 => to_unsigned(771, 10), 170 => to_unsigned(126, 10), 171 => to_unsigned(264, 10), 172 => to_unsigned(47, 10), 173 => to_unsigned(555, 10), 174 => to_unsigned(701, 10), 175 => to_unsigned(771, 10), 176 => to_unsigned(300, 10), 177 => to_unsigned(75, 10), 178 => to_unsigned(1013, 10), 179 => to_unsigned(305, 10), 180 => to_unsigned(50, 10), 181 => to_unsigned(138, 10), 182 => to_unsigned(171, 10), 183 => to_unsigned(719, 10), 184 => to_unsigned(987, 10), 185 => to_unsigned(102, 10), 186 => to_unsigned(574, 10), 187 => to_unsigned(483, 10), 188 => to_unsigned(338, 10), 189 => to_unsigned(765, 10), 190 => to_unsigned(318, 10), 191 => to_unsigned(373, 10), 192 => to_unsigned(419, 10), 193 => to_unsigned(341, 10), 194 => to_unsigned(924, 10), 195 => to_unsigned(955, 10), 196 => to_unsigned(225, 10), 197 => to_unsigned(89, 10), 198 => to_unsigned(458, 10), 199 => to_unsigned(513, 10), 200 => to_unsigned(506, 10), 201 => to_unsigned(405, 10), 202 => to_unsigned(921, 10), 203 => to_unsigned(650, 10), 204 => to_unsigned(632, 10), 205 => to_unsigned(425, 10), 206 => to_unsigned(13, 10), 207 => to_unsigned(691, 10), 208 => to_unsigned(322, 10), 209 => to_unsigned(210, 10), 210 => to_unsigned(212, 10), 211 => to_unsigned(647, 10), 212 => to_unsigned(808, 10), 213 => to_unsigned(312, 10), 214 => to_unsigned(341, 10), 215 => to_unsigned(37, 10), 216 => to_unsigned(430, 10), 217 => to_unsigned(211, 10), 218 => to_unsigned(474, 10), 219 => to_unsigned(695, 10), 220 => to_unsigned(390, 10), 221 => to_unsigned(512, 10), 222 => to_unsigned(392, 10), 223 => to_unsigned(1020, 10), 224 => to_unsigned(725, 10), 225 => to_unsigned(379, 10), 226 => to_unsigned(239, 10), 227 => to_unsigned(677, 10), 228 => to_unsigned(963, 10), 229 => to_unsigned(686, 10), 230 => to_unsigned(744, 10), 231 => to_unsigned(425, 10), 232 => to_unsigned(860, 10), 233 => to_unsigned(63, 10), 234 => to_unsigned(57, 10), 235 => to_unsigned(1015, 10), 236 => to_unsigned(612, 10), 237 => to_unsigned(551, 10), 238 => to_unsigned(705, 10), 239 => to_unsigned(435, 10), 240 => to_unsigned(701, 10), 241 => to_unsigned(365, 10), 242 => to_unsigned(709, 10), 243 => to_unsigned(954, 10), 244 => to_unsigned(859, 10), 245 => to_unsigned(351, 10), 246 => to_unsigned(936, 10), 247 => to_unsigned(73, 10), 248 => to_unsigned(693, 10), 249 => to_unsigned(888, 10), 250 => to_unsigned(519, 10), 251 => to_unsigned(355, 10), 252 => to_unsigned(943, 10), 253 => to_unsigned(709, 10), 254 => to_unsigned(681, 10), 255 => to_unsigned(796, 10), 256 => to_unsigned(246, 10), 257 => to_unsigned(890, 10), 258 => to_unsigned(853, 10), 259 => to_unsigned(779, 10), 260 => to_unsigned(515, 10), 261 => to_unsigned(274, 10), 262 => to_unsigned(931, 10), 263 => to_unsigned(46, 10), 264 => to_unsigned(361, 10), 265 => to_unsigned(145, 10), 266 => to_unsigned(111, 10), 267 => to_unsigned(155, 10), 268 => to_unsigned(54, 10), 269 => to_unsigned(623, 10), 270 => to_unsigned(713, 10), 271 => to_unsigned(403, 10), 272 => to_unsigned(199, 10), 273 => to_unsigned(583, 10), 274 => to_unsigned(869, 10), 275 => to_unsigned(427, 10), 276 => to_unsigned(1022, 10), 277 => to_unsigned(940, 10), 278 => to_unsigned(622, 10), 279 => to_unsigned(686, 10), 280 => to_unsigned(674, 10), 281 => to_unsigned(673, 10), 282 => to_unsigned(74, 10), 283 => to_unsigned(375, 10), 284 => to_unsigned(837, 10), 285 => to_unsigned(476, 10), 286 => to_unsigned(814, 10), 287 => to_unsigned(928, 10), 288 => to_unsigned(211, 10), 289 => to_unsigned(423, 10), 290 => to_unsigned(414, 10), 291 => to_unsigned(223, 10), 292 => to_unsigned(879, 10), 293 => to_unsigned(175, 10), 294 => to_unsigned(897, 10), 295 => to_unsigned(928, 10), 296 => to_unsigned(894, 10), 297 => to_unsigned(104, 10), 298 => to_unsigned(369, 10), 299 => to_unsigned(703, 10), 300 => to_unsigned(119, 10), 301 => to_unsigned(301, 10), 302 => to_unsigned(183, 10), 303 => to_unsigned(110, 10), 304 => to_unsigned(886, 10), 305 => to_unsigned(320, 10), 306 => to_unsigned(869, 10), 307 => to_unsigned(469, 10), 308 => to_unsigned(662, 10), 309 => to_unsigned(411, 10), 310 => to_unsigned(5, 10), 311 => to_unsigned(877, 10), 312 => to_unsigned(35, 10), 313 => to_unsigned(877, 10), 314 => to_unsigned(803, 10), 315 => to_unsigned(636, 10), 316 => to_unsigned(616, 10), 317 => to_unsigned(195, 10), 318 => to_unsigned(156, 10), 319 => to_unsigned(603, 10), 320 => to_unsigned(763, 10), 321 => to_unsigned(137, 10), 322 => to_unsigned(299, 10), 323 => to_unsigned(643, 10), 324 => to_unsigned(107, 10), 325 => to_unsigned(907, 10), 326 => to_unsigned(947, 10), 327 => to_unsigned(470, 10), 328 => to_unsigned(618, 10), 329 => to_unsigned(746, 10), 330 => to_unsigned(132, 10), 331 => to_unsigned(669, 10), 332 => to_unsigned(316, 10), 333 => to_unsigned(428, 10), 334 => to_unsigned(2, 10), 335 => to_unsigned(990, 10), 336 => to_unsigned(69, 10), 337 => to_unsigned(559, 10), 338 => to_unsigned(204, 10), 339 => to_unsigned(657, 10), 340 => to_unsigned(79, 10), 341 => to_unsigned(696, 10), 342 => to_unsigned(553, 10), 343 => to_unsigned(920, 10), 344 => to_unsigned(725, 10), 345 => to_unsigned(616, 10), 346 => to_unsigned(515, 10), 347 => to_unsigned(700, 10), 348 => to_unsigned(814, 10), 349 => to_unsigned(368, 10), 350 => to_unsigned(159, 10), 351 => to_unsigned(454, 10), 352 => to_unsigned(1023, 10), 353 => to_unsigned(819, 10), 354 => to_unsigned(97, 10), 355 => to_unsigned(175, 10), 356 => to_unsigned(267, 10), 357 => to_unsigned(871, 10), 358 => to_unsigned(318, 10), 359 => to_unsigned(648, 10), 360 => to_unsigned(190, 10), 361 => to_unsigned(131, 10), 362 => to_unsigned(951, 10), 363 => to_unsigned(107, 10), 364 => to_unsigned(822, 10), 365 => to_unsigned(743, 10), 366 => to_unsigned(169, 10), 367 => to_unsigned(310, 10), 368 => to_unsigned(281, 10), 369 => to_unsigned(877, 10), 370 => to_unsigned(390, 10), 371 => to_unsigned(71, 10), 372 => to_unsigned(744, 10), 373 => to_unsigned(959, 10), 374 => to_unsigned(349, 10), 375 => to_unsigned(766, 10), 376 => to_unsigned(965, 10), 377 => to_unsigned(550, 10), 378 => to_unsigned(963, 10), 379 => to_unsigned(263, 10), 380 => to_unsigned(370, 10), 381 => to_unsigned(939, 10), 382 => to_unsigned(919, 10), 383 => to_unsigned(216, 10), 384 => to_unsigned(1010, 10), 385 => to_unsigned(797, 10), 386 => to_unsigned(307, 10), 387 => to_unsigned(913, 10), 388 => to_unsigned(696, 10), 389 => to_unsigned(299, 10), 390 => to_unsigned(929, 10), 391 => to_unsigned(816, 10), 392 => to_unsigned(718, 10), 393 => to_unsigned(874, 10), 394 => to_unsigned(426, 10), 395 => to_unsigned(720, 10), 396 => to_unsigned(239, 10), 397 => to_unsigned(1013, 10), 398 => to_unsigned(129, 10), 399 => to_unsigned(362, 10), 400 => to_unsigned(565, 10), 401 => to_unsigned(448, 10), 402 => to_unsigned(755, 10), 403 => to_unsigned(383, 10), 404 => to_unsigned(56, 10), 405 => to_unsigned(143, 10), 406 => to_unsigned(336, 10), 407 => to_unsigned(200, 10), 408 => to_unsigned(361, 10), 409 => to_unsigned(660, 10), 410 => to_unsigned(701, 10), 411 => to_unsigned(191, 10), 412 => to_unsigned(822, 10), 413 => to_unsigned(427, 10), 414 => to_unsigned(409, 10), 415 => to_unsigned(128, 10), 416 => to_unsigned(123, 10), 417 => to_unsigned(305, 10), 418 => to_unsigned(423, 10), 419 => to_unsigned(386, 10), 420 => to_unsigned(198, 10), 421 => to_unsigned(899, 10), 422 => to_unsigned(798, 10), 423 => to_unsigned(781, 10), 424 => to_unsigned(788, 10), 425 => to_unsigned(884, 10), 426 => to_unsigned(331, 10), 427 => to_unsigned(267, 10), 428 => to_unsigned(645, 10), 429 => to_unsigned(880, 10), 430 => to_unsigned(656, 10), 431 => to_unsigned(461, 10), 432 => to_unsigned(190, 10), 433 => to_unsigned(392, 10), 434 => to_unsigned(27, 10), 435 => to_unsigned(902, 10), 436 => to_unsigned(364, 10), 437 => to_unsigned(758, 10), 438 => to_unsigned(554, 10), 439 => to_unsigned(644, 10), 440 => to_unsigned(1000, 10), 441 => to_unsigned(745, 10), 442 => to_unsigned(399, 10), 443 => to_unsigned(956, 10), 444 => to_unsigned(384, 10), 445 => to_unsigned(167, 10), 446 => to_unsigned(549, 10), 447 => to_unsigned(518, 10), 448 => to_unsigned(755, 10), 449 => to_unsigned(605, 10), 450 => to_unsigned(826, 10), 451 => to_unsigned(879, 10), 452 => to_unsigned(921, 10), 453 => to_unsigned(588, 10), 454 => to_unsigned(64, 10), 455 => to_unsigned(958, 10), 456 => to_unsigned(948, 10), 457 => to_unsigned(50, 10), 458 => to_unsigned(177, 10), 459 => to_unsigned(412, 10), 460 => to_unsigned(1018, 10), 461 => to_unsigned(967, 10), 462 => to_unsigned(449, 10), 463 => to_unsigned(620, 10), 464 => to_unsigned(752, 10), 465 => to_unsigned(50, 10), 466 => to_unsigned(391, 10), 467 => to_unsigned(1000, 10), 468 => to_unsigned(794, 10), 469 => to_unsigned(680, 10), 470 => to_unsigned(317, 10), 471 => to_unsigned(688, 10), 472 => to_unsigned(494, 10), 473 => to_unsigned(150, 10), 474 => to_unsigned(782, 10), 475 => to_unsigned(319, 10), 476 => to_unsigned(479, 10), 477 => to_unsigned(853, 10), 478 => to_unsigned(564, 10), 479 => to_unsigned(391, 10), 480 => to_unsigned(36, 10), 481 => to_unsigned(464, 10), 482 => to_unsigned(710, 10), 483 => to_unsigned(234, 10), 484 => to_unsigned(404, 10), 485 => to_unsigned(550, 10), 486 => to_unsigned(388, 10), 487 => to_unsigned(144, 10), 488 => to_unsigned(738, 10), 489 => to_unsigned(111, 10), 490 => to_unsigned(184, 10), 491 => to_unsigned(251, 10), 492 => to_unsigned(879, 10), 493 => to_unsigned(782, 10), 494 => to_unsigned(1007, 10), 495 => to_unsigned(743, 10), 496 => to_unsigned(127, 10), 497 => to_unsigned(15, 10), 498 => to_unsigned(472, 10), 499 => to_unsigned(654, 10), 500 => to_unsigned(906, 10), 501 => to_unsigned(758, 10), 502 => to_unsigned(260, 10), 503 => to_unsigned(596, 10), 504 => to_unsigned(105, 10), 505 => to_unsigned(744, 10), 506 => to_unsigned(564, 10), 507 => to_unsigned(715, 10), 508 => to_unsigned(252, 10), 509 => to_unsigned(821, 10), 510 => to_unsigned(477, 10), 511 => to_unsigned(835, 10), 512 => to_unsigned(244, 10), 513 => to_unsigned(812, 10), 514 => to_unsigned(218, 10), 515 => to_unsigned(380, 10), 516 => to_unsigned(219, 10), 517 => to_unsigned(770, 10), 518 => to_unsigned(188, 10), 519 => to_unsigned(66, 10), 520 => to_unsigned(509, 10), 521 => to_unsigned(535, 10), 522 => to_unsigned(749, 10), 523 => to_unsigned(28, 10), 524 => to_unsigned(249, 10), 525 => to_unsigned(821, 10), 526 => to_unsigned(914, 10), 527 => to_unsigned(879, 10), 528 => to_unsigned(955, 10), 529 => to_unsigned(577, 10), 530 => to_unsigned(68, 10), 531 => to_unsigned(36, 10), 532 => to_unsigned(849, 10), 533 => to_unsigned(24, 10), 534 => to_unsigned(729, 10), 535 => to_unsigned(875, 10), 536 => to_unsigned(332, 10), 537 => to_unsigned(290, 10), 538 => to_unsigned(341, 10), 539 => to_unsigned(824, 10), 540 => to_unsigned(1010, 10), 541 => to_unsigned(575, 10), 542 => to_unsigned(969, 10), 543 => to_unsigned(292, 10), 544 => to_unsigned(875, 10), 545 => to_unsigned(425, 10), 546 => to_unsigned(262, 10), 547 => to_unsigned(913, 10), 548 => to_unsigned(287, 10), 549 => to_unsigned(506, 10), 550 => to_unsigned(626, 10), 551 => to_unsigned(239, 10), 552 => to_unsigned(1004, 10), 553 => to_unsigned(518, 10), 554 => to_unsigned(178, 10), 555 => to_unsigned(784, 10), 556 => to_unsigned(798, 10), 557 => to_unsigned(796, 10), 558 => to_unsigned(127, 10), 559 => to_unsigned(459, 10), 560 => to_unsigned(160, 10), 561 => to_unsigned(870, 10), 562 => to_unsigned(473, 10), 563 => to_unsigned(550, 10), 564 => to_unsigned(285, 10), 565 => to_unsigned(258, 10), 566 => to_unsigned(595, 10), 567 => to_unsigned(332, 10), 568 => to_unsigned(914, 10), 569 => to_unsigned(64, 10), 570 => to_unsigned(425, 10), 571 => to_unsigned(150, 10), 572 => to_unsigned(529, 10), 573 => to_unsigned(682, 10), 574 => to_unsigned(4, 10), 575 => to_unsigned(132, 10), 576 => to_unsigned(402, 10), 577 => to_unsigned(709, 10), 578 => to_unsigned(14, 10), 579 => to_unsigned(10, 10), 580 => to_unsigned(306, 10), 581 => to_unsigned(989, 10), 582 => to_unsigned(723, 10), 583 => to_unsigned(802, 10), 584 => to_unsigned(3, 10), 585 => to_unsigned(8, 10), 586 => to_unsigned(986, 10), 587 => to_unsigned(594, 10), 588 => to_unsigned(580, 10), 589 => to_unsigned(647, 10), 590 => to_unsigned(362, 10), 591 => to_unsigned(349, 10), 592 => to_unsigned(35, 10), 593 => to_unsigned(719, 10), 594 => to_unsigned(46, 10), 595 => to_unsigned(173, 10), 596 => to_unsigned(451, 10), 597 => to_unsigned(570, 10), 598 => to_unsigned(643, 10), 599 => to_unsigned(198, 10), 600 => to_unsigned(66, 10), 601 => to_unsigned(997, 10), 602 => to_unsigned(664, 10), 603 => to_unsigned(695, 10), 604 => to_unsigned(443, 10), 605 => to_unsigned(675, 10), 606 => to_unsigned(259, 10), 607 => to_unsigned(583, 10), 608 => to_unsigned(923, 10), 609 => to_unsigned(1010, 10), 610 => to_unsigned(834, 10), 611 => to_unsigned(510, 10), 612 => to_unsigned(368, 10), 613 => to_unsigned(583, 10), 614 => to_unsigned(10, 10), 615 => to_unsigned(109, 10), 616 => to_unsigned(191, 10), 617 => to_unsigned(379, 10), 618 => to_unsigned(112, 10), 619 => to_unsigned(377, 10), 620 => to_unsigned(5, 10), 621 => to_unsigned(500, 10), 622 => to_unsigned(296, 10), 623 => to_unsigned(982, 10), 624 => to_unsigned(436, 10), 625 => to_unsigned(939, 10), 626 => to_unsigned(449, 10), 627 => to_unsigned(902, 10), 628 => to_unsigned(796, 10), 629 => to_unsigned(389, 10), 630 => to_unsigned(232, 10), 631 => to_unsigned(586, 10), 632 => to_unsigned(647, 10), 633 => to_unsigned(797, 10), 634 => to_unsigned(868, 10), 635 => to_unsigned(338, 10), 636 => to_unsigned(47, 10), 637 => to_unsigned(444, 10), 638 => to_unsigned(319, 10), 639 => to_unsigned(635, 10), 640 => to_unsigned(450, 10), 641 => to_unsigned(297, 10), 642 => to_unsigned(541, 10), 643 => to_unsigned(96, 10), 644 => to_unsigned(561, 10), 645 => to_unsigned(700, 10), 646 => to_unsigned(820, 10), 647 => to_unsigned(537, 10), 648 => to_unsigned(548, 10), 649 => to_unsigned(659, 10), 650 => to_unsigned(864, 10), 651 => to_unsigned(245, 10), 652 => to_unsigned(603, 10), 653 => to_unsigned(154, 10), 654 => to_unsigned(568, 10), 655 => to_unsigned(312, 10), 656 => to_unsigned(796, 10), 657 => to_unsigned(941, 10), 658 => to_unsigned(983, 10), 659 => to_unsigned(466, 10), 660 => to_unsigned(261, 10), 661 => to_unsigned(961, 10), 662 => to_unsigned(597, 10), 663 => to_unsigned(290, 10), 664 => to_unsigned(897, 10), 665 => to_unsigned(605, 10), 666 => to_unsigned(749, 10), 667 => to_unsigned(994, 10), 668 => to_unsigned(270, 10), 669 => to_unsigned(234, 10), 670 => to_unsigned(542, 10), 671 => to_unsigned(905, 10), 672 => to_unsigned(438, 10), 673 => to_unsigned(795, 10), 674 => to_unsigned(391, 10), 675 => to_unsigned(972, 10), 676 => to_unsigned(349, 10), 677 => to_unsigned(676, 10), 678 => to_unsigned(166, 10), 679 => to_unsigned(92, 10), 680 => to_unsigned(625, 10), 681 => to_unsigned(597, 10), 682 => to_unsigned(215, 10), 683 => to_unsigned(421, 10), 684 => to_unsigned(916, 10), 685 => to_unsigned(781, 10), 686 => to_unsigned(109, 10), 687 => to_unsigned(680, 10), 688 => to_unsigned(434, 10), 689 => to_unsigned(489, 10), 690 => to_unsigned(310, 10), 691 => to_unsigned(126, 10), 692 => to_unsigned(449, 10), 693 => to_unsigned(840, 10), 694 => to_unsigned(58, 10), 695 => to_unsigned(103, 10), 696 => to_unsigned(876, 10), 697 => to_unsigned(73, 10), 698 => to_unsigned(561, 10), 699 => to_unsigned(273, 10), 700 => to_unsigned(305, 10), 701 => to_unsigned(89, 10), 702 => to_unsigned(471, 10), 703 => to_unsigned(953, 10), 704 => to_unsigned(1000, 10), 705 => to_unsigned(249, 10), 706 => to_unsigned(115, 10), 707 => to_unsigned(714, 10), 708 => to_unsigned(858, 10), 709 => to_unsigned(269, 10), 710 => to_unsigned(287, 10), 711 => to_unsigned(124, 10), 712 => to_unsigned(533, 10), 713 => to_unsigned(865, 10), 714 => to_unsigned(493, 10), 715 => to_unsigned(257, 10), 716 => to_unsigned(480, 10), 717 => to_unsigned(171, 10), 718 => to_unsigned(695, 10), 719 => to_unsigned(838, 10), 720 => to_unsigned(290, 10), 721 => to_unsigned(990, 10), 722 => to_unsigned(558, 10), 723 => to_unsigned(346, 10), 724 => to_unsigned(486, 10), 725 => to_unsigned(996, 10), 726 => to_unsigned(657, 10), 727 => to_unsigned(880, 10), 728 => to_unsigned(268, 10), 729 => to_unsigned(564, 10), 730 => to_unsigned(815, 10), 731 => to_unsigned(372, 10), 732 => to_unsigned(935, 10), 733 => to_unsigned(880, 10), 734 => to_unsigned(944, 10), 735 => to_unsigned(951, 10), 736 => to_unsigned(665, 10), 737 => to_unsigned(832, 10), 738 => to_unsigned(316, 10), 739 => to_unsigned(998, 10), 740 => to_unsigned(158, 10), 741 => to_unsigned(233, 10), 742 => to_unsigned(751, 10), 743 => to_unsigned(100, 10), 744 => to_unsigned(614, 10), 745 => to_unsigned(860, 10), 746 => to_unsigned(490, 10), 747 => to_unsigned(727, 10), 748 => to_unsigned(591, 10), 749 => to_unsigned(422, 10), 750 => to_unsigned(358, 10), 751 => to_unsigned(982, 10), 752 => to_unsigned(816, 10), 753 => to_unsigned(263, 10), 754 => to_unsigned(549, 10), 755 => to_unsigned(242, 10), 756 => to_unsigned(834, 10), 757 => to_unsigned(77, 10), 758 => to_unsigned(276, 10), 759 => to_unsigned(814, 10), 760 => to_unsigned(477, 10), 761 => to_unsigned(288, 10), 762 => to_unsigned(820, 10), 763 => to_unsigned(439, 10), 764 => to_unsigned(403, 10), 765 => to_unsigned(1004, 10), 766 => to_unsigned(1004, 10), 767 => to_unsigned(440, 10), 768 => to_unsigned(534, 10), 769 => to_unsigned(86, 10), 770 => to_unsigned(492, 10), 771 => to_unsigned(229, 10), 772 => to_unsigned(572, 10), 773 => to_unsigned(674, 10), 774 => to_unsigned(573, 10), 775 => to_unsigned(950, 10), 776 => to_unsigned(38, 10), 777 => to_unsigned(725, 10), 778 => to_unsigned(988, 10), 779 => to_unsigned(688, 10), 780 => to_unsigned(418, 10), 781 => to_unsigned(957, 10), 782 => to_unsigned(705, 10), 783 => to_unsigned(182, 10), 784 => to_unsigned(877, 10), 785 => to_unsigned(238, 10), 786 => to_unsigned(145, 10), 787 => to_unsigned(564, 10), 788 => to_unsigned(290, 10), 789 => to_unsigned(939, 10), 790 => to_unsigned(141, 10), 791 => to_unsigned(17, 10), 792 => to_unsigned(799, 10), 793 => to_unsigned(533, 10), 794 => to_unsigned(226, 10), 795 => to_unsigned(621, 10), 796 => to_unsigned(641, 10), 797 => to_unsigned(581, 10), 798 => to_unsigned(943, 10), 799 => to_unsigned(242, 10), 800 => to_unsigned(166, 10), 801 => to_unsigned(831, 10), 802 => to_unsigned(159, 10), 803 => to_unsigned(860, 10), 804 => to_unsigned(102, 10), 805 => to_unsigned(762, 10), 806 => to_unsigned(114, 10), 807 => to_unsigned(240, 10), 808 => to_unsigned(836, 10), 809 => to_unsigned(421, 10), 810 => to_unsigned(903, 10), 811 => to_unsigned(579, 10), 812 => to_unsigned(54, 10), 813 => to_unsigned(21, 10), 814 => to_unsigned(149, 10), 815 => to_unsigned(313, 10), 816 => to_unsigned(986, 10), 817 => to_unsigned(322, 10), 818 => to_unsigned(732, 10), 819 => to_unsigned(815, 10), 820 => to_unsigned(32, 10), 821 => to_unsigned(229, 10), 822 => to_unsigned(673, 10), 823 => to_unsigned(227, 10), 824 => to_unsigned(954, 10), 825 => to_unsigned(928, 10), 826 => to_unsigned(615, 10), 827 => to_unsigned(145, 10), 828 => to_unsigned(905, 10), 829 => to_unsigned(611, 10), 830 => to_unsigned(940, 10), 831 => to_unsigned(598, 10), 832 => to_unsigned(261, 10), 833 => to_unsigned(982, 10), 834 => to_unsigned(649, 10), 835 => to_unsigned(118, 10), 836 => to_unsigned(321, 10), 837 => to_unsigned(701, 10), 838 => to_unsigned(235, 10), 839 => to_unsigned(133, 10), 840 => to_unsigned(234, 10), 841 => to_unsigned(196, 10), 842 => to_unsigned(647, 10), 843 => to_unsigned(950, 10), 844 => to_unsigned(19, 10), 845 => to_unsigned(1010, 10), 846 => to_unsigned(819, 10), 847 => to_unsigned(934, 10), 848 => to_unsigned(1013, 10), 849 => to_unsigned(759, 10), 850 => to_unsigned(653, 10), 851 => to_unsigned(11, 10), 852 => to_unsigned(855, 10), 853 => to_unsigned(358, 10), 854 => to_unsigned(566, 10), 855 => to_unsigned(181, 10), 856 => to_unsigned(587, 10), 857 => to_unsigned(296, 10), 858 => to_unsigned(1013, 10), 859 => to_unsigned(607, 10), 860 => to_unsigned(515, 10), 861 => to_unsigned(503, 10), 862 => to_unsigned(701, 10), 863 => to_unsigned(130, 10), 864 => to_unsigned(967, 10), 865 => to_unsigned(258, 10), 866 => to_unsigned(281, 10), 867 => to_unsigned(814, 10), 868 => to_unsigned(389, 10), 869 => to_unsigned(16, 10), 870 => to_unsigned(114, 10), 871 => to_unsigned(136, 10), 872 => to_unsigned(721, 10), 873 => to_unsigned(120, 10), 874 => to_unsigned(370, 10), 875 => to_unsigned(604, 10), 876 => to_unsigned(590, 10), 877 => to_unsigned(440, 10), 878 => to_unsigned(518, 10), 879 => to_unsigned(589, 10), 880 => to_unsigned(568, 10), 881 => to_unsigned(988, 10), 882 => to_unsigned(771, 10), 883 => to_unsigned(492, 10), 884 => to_unsigned(315, 10), 885 => to_unsigned(614, 10), 886 => to_unsigned(367, 10), 887 => to_unsigned(4, 10), 888 => to_unsigned(0, 10), 889 => to_unsigned(715, 10), 890 => to_unsigned(934, 10), 891 => to_unsigned(134, 10), 892 => to_unsigned(883, 10), 893 => to_unsigned(660, 10), 894 => to_unsigned(504, 10), 895 => to_unsigned(710, 10), 896 => to_unsigned(912, 10), 897 => to_unsigned(832, 10), 898 => to_unsigned(323, 10), 899 => to_unsigned(123, 10), 900 => to_unsigned(69, 10), 901 => to_unsigned(367, 10), 902 => to_unsigned(61, 10), 903 => to_unsigned(295, 10), 904 => to_unsigned(315, 10), 905 => to_unsigned(208, 10), 906 => to_unsigned(473, 10), 907 => to_unsigned(505, 10), 908 => to_unsigned(990, 10), 909 => to_unsigned(283, 10), 910 => to_unsigned(203, 10), 911 => to_unsigned(1000, 10), 912 => to_unsigned(960, 10), 913 => to_unsigned(289, 10), 914 => to_unsigned(281, 10), 915 => to_unsigned(692, 10), 916 => to_unsigned(910, 10), 917 => to_unsigned(688, 10), 918 => to_unsigned(418, 10), 919 => to_unsigned(628, 10), 920 => to_unsigned(552, 10), 921 => to_unsigned(946, 10), 922 => to_unsigned(702, 10), 923 => to_unsigned(114, 10), 924 => to_unsigned(299, 10), 925 => to_unsigned(631, 10), 926 => to_unsigned(38, 10), 927 => to_unsigned(147, 10), 928 => to_unsigned(810, 10), 929 => to_unsigned(482, 10), 930 => to_unsigned(742, 10), 931 => to_unsigned(149, 10), 932 => to_unsigned(916, 10), 933 => to_unsigned(346, 10), 934 => to_unsigned(419, 10), 935 => to_unsigned(923, 10), 936 => to_unsigned(643, 10), 937 => to_unsigned(985, 10), 938 => to_unsigned(892, 10), 939 => to_unsigned(391, 10), 940 => to_unsigned(260, 10), 941 => to_unsigned(516, 10), 942 => to_unsigned(53, 10), 943 => to_unsigned(393, 10), 944 => to_unsigned(964, 10), 945 => to_unsigned(673, 10), 946 => to_unsigned(945, 10), 947 => to_unsigned(714, 10), 948 => to_unsigned(919, 10), 949 => to_unsigned(953, 10), 950 => to_unsigned(752, 10), 951 => to_unsigned(992, 10), 952 => to_unsigned(845, 10), 953 => to_unsigned(405, 10), 954 => to_unsigned(92, 10), 955 => to_unsigned(23, 10), 956 => to_unsigned(112, 10), 957 => to_unsigned(389, 10), 958 => to_unsigned(957, 10), 959 => to_unsigned(2, 10), 960 => to_unsigned(256, 10), 961 => to_unsigned(777, 10), 962 => to_unsigned(839, 10), 963 => to_unsigned(925, 10), 964 => to_unsigned(149, 10), 965 => to_unsigned(464, 10), 966 => to_unsigned(590, 10), 967 => to_unsigned(979, 10), 968 => to_unsigned(549, 10), 969 => to_unsigned(602, 10), 970 => to_unsigned(76, 10), 971 => to_unsigned(335, 10), 972 => to_unsigned(723, 10), 973 => to_unsigned(146, 10), 974 => to_unsigned(490, 10), 975 => to_unsigned(578, 10), 976 => to_unsigned(784, 10), 977 => to_unsigned(1016, 10), 978 => to_unsigned(331, 10), 979 => to_unsigned(995, 10), 980 => to_unsigned(521, 10), 981 => to_unsigned(377, 10), 982 => to_unsigned(329, 10), 983 => to_unsigned(798, 10), 984 => to_unsigned(22, 10), 985 => to_unsigned(618, 10), 986 => to_unsigned(276, 10), 987 => to_unsigned(617, 10), 988 => to_unsigned(467, 10), 989 => to_unsigned(324, 10), 990 => to_unsigned(366, 10), 991 => to_unsigned(79, 10), 992 => to_unsigned(417, 10), 993 => to_unsigned(960, 10), 994 => to_unsigned(879, 10), 995 => to_unsigned(911, 10), 996 => to_unsigned(333, 10), 997 => to_unsigned(905, 10), 998 => to_unsigned(49, 10), 999 => to_unsigned(746, 10), 1000 => to_unsigned(138, 10), 1001 => to_unsigned(369, 10), 1002 => to_unsigned(615, 10), 1003 => to_unsigned(546, 10), 1004 => to_unsigned(935, 10), 1005 => to_unsigned(944, 10), 1006 => to_unsigned(300, 10), 1007 => to_unsigned(748, 10), 1008 => to_unsigned(618, 10), 1009 => to_unsigned(257, 10), 1010 => to_unsigned(968, 10), 1011 => to_unsigned(256, 10), 1012 => to_unsigned(139, 10), 1013 => to_unsigned(922, 10), 1014 => to_unsigned(478, 10), 1015 => to_unsigned(875, 10), 1016 => to_unsigned(938, 10), 1017 => to_unsigned(787, 10), 1018 => to_unsigned(853, 10), 1019 => to_unsigned(879, 10), 1020 => to_unsigned(769, 10), 1021 => to_unsigned(506, 10), 1022 => to_unsigned(956, 10), 1023 => to_unsigned(594, 10), 1024 => to_unsigned(476, 10), 1025 => to_unsigned(574, 10), 1026 => to_unsigned(907, 10), 1027 => to_unsigned(1019, 10), 1028 => to_unsigned(689, 10), 1029 => to_unsigned(191, 10), 1030 => to_unsigned(884, 10), 1031 => to_unsigned(615, 10), 1032 => to_unsigned(649, 10), 1033 => to_unsigned(24, 10), 1034 => to_unsigned(68, 10), 1035 => to_unsigned(794, 10), 1036 => to_unsigned(820, 10), 1037 => to_unsigned(107, 10), 1038 => to_unsigned(566, 10), 1039 => to_unsigned(469, 10), 1040 => to_unsigned(718, 10), 1041 => to_unsigned(157, 10), 1042 => to_unsigned(897, 10), 1043 => to_unsigned(206, 10), 1044 => to_unsigned(256, 10), 1045 => to_unsigned(527, 10), 1046 => to_unsigned(417, 10), 1047 => to_unsigned(672, 10), 1048 => to_unsigned(765, 10), 1049 => to_unsigned(755, 10), 1050 => to_unsigned(741, 10), 1051 => to_unsigned(197, 10), 1052 => to_unsigned(926, 10), 1053 => to_unsigned(502, 10), 1054 => to_unsigned(105, 10), 1055 => to_unsigned(687, 10), 1056 => to_unsigned(498, 10), 1057 => to_unsigned(570, 10), 1058 => to_unsigned(969, 10), 1059 => to_unsigned(373, 10), 1060 => to_unsigned(903, 10), 1061 => to_unsigned(1022, 10), 1062 => to_unsigned(926, 10), 1063 => to_unsigned(341, 10), 1064 => to_unsigned(30, 10), 1065 => to_unsigned(425, 10), 1066 => to_unsigned(8, 10), 1067 => to_unsigned(65, 10), 1068 => to_unsigned(621, 10), 1069 => to_unsigned(469, 10), 1070 => to_unsigned(264, 10), 1071 => to_unsigned(249, 10), 1072 => to_unsigned(749, 10), 1073 => to_unsigned(49, 10), 1074 => to_unsigned(372, 10), 1075 => to_unsigned(64, 10), 1076 => to_unsigned(603, 10), 1077 => to_unsigned(50, 10), 1078 => to_unsigned(176, 10), 1079 => to_unsigned(473, 10), 1080 => to_unsigned(669, 10), 1081 => to_unsigned(583, 10), 1082 => to_unsigned(538, 10), 1083 => to_unsigned(479, 10), 1084 => to_unsigned(398, 10), 1085 => to_unsigned(889, 10), 1086 => to_unsigned(787, 10), 1087 => to_unsigned(126, 10), 1088 => to_unsigned(136, 10), 1089 => to_unsigned(39, 10), 1090 => to_unsigned(925, 10), 1091 => to_unsigned(279, 10), 1092 => to_unsigned(845, 10), 1093 => to_unsigned(40, 10), 1094 => to_unsigned(129, 10), 1095 => to_unsigned(857, 10), 1096 => to_unsigned(472, 10), 1097 => to_unsigned(798, 10), 1098 => to_unsigned(425, 10), 1099 => to_unsigned(848, 10), 1100 => to_unsigned(380, 10), 1101 => to_unsigned(830, 10), 1102 => to_unsigned(843, 10), 1103 => to_unsigned(871, 10), 1104 => to_unsigned(839, 10), 1105 => to_unsigned(614, 10), 1106 => to_unsigned(469, 10), 1107 => to_unsigned(984, 10), 1108 => to_unsigned(293, 10), 1109 => to_unsigned(811, 10), 1110 => to_unsigned(443, 10), 1111 => to_unsigned(676, 10), 1112 => to_unsigned(672, 10), 1113 => to_unsigned(841, 10), 1114 => to_unsigned(753, 10), 1115 => to_unsigned(767, 10), 1116 => to_unsigned(1000, 10), 1117 => to_unsigned(912, 10), 1118 => to_unsigned(419, 10), 1119 => to_unsigned(759, 10), 1120 => to_unsigned(387, 10), 1121 => to_unsigned(551, 10), 1122 => to_unsigned(421, 10), 1123 => to_unsigned(506, 10), 1124 => to_unsigned(259, 10), 1125 => to_unsigned(424, 10), 1126 => to_unsigned(570, 10), 1127 => to_unsigned(483, 10), 1128 => to_unsigned(641, 10), 1129 => to_unsigned(515, 10), 1130 => to_unsigned(523, 10), 1131 => to_unsigned(387, 10), 1132 => to_unsigned(110, 10), 1133 => to_unsigned(510, 10), 1134 => to_unsigned(699, 10), 1135 => to_unsigned(140, 10), 1136 => to_unsigned(864, 10), 1137 => to_unsigned(935, 10), 1138 => to_unsigned(818, 10), 1139 => to_unsigned(768, 10), 1140 => to_unsigned(566, 10), 1141 => to_unsigned(54, 10), 1142 => to_unsigned(623, 10), 1143 => to_unsigned(855, 10), 1144 => to_unsigned(711, 10), 1145 => to_unsigned(699, 10), 1146 => to_unsigned(321, 10), 1147 => to_unsigned(482, 10), 1148 => to_unsigned(781, 10), 1149 => to_unsigned(952, 10), 1150 => to_unsigned(30, 10), 1151 => to_unsigned(341, 10), 1152 => to_unsigned(593, 10), 1153 => to_unsigned(663, 10), 1154 => to_unsigned(931, 10), 1155 => to_unsigned(929, 10), 1156 => to_unsigned(902, 10), 1157 => to_unsigned(24, 10), 1158 => to_unsigned(34, 10), 1159 => to_unsigned(1015, 10), 1160 => to_unsigned(616, 10), 1161 => to_unsigned(441, 10), 1162 => to_unsigned(358, 10), 1163 => to_unsigned(457, 10), 1164 => to_unsigned(664, 10), 1165 => to_unsigned(733, 10), 1166 => to_unsigned(517, 10), 1167 => to_unsigned(240, 10), 1168 => to_unsigned(944, 10), 1169 => to_unsigned(921, 10), 1170 => to_unsigned(452, 10), 1171 => to_unsigned(750, 10), 1172 => to_unsigned(38, 10), 1173 => to_unsigned(384, 10), 1174 => to_unsigned(315, 10), 1175 => to_unsigned(206, 10), 1176 => to_unsigned(73, 10), 1177 => to_unsigned(228, 10), 1178 => to_unsigned(495, 10), 1179 => to_unsigned(946, 10), 1180 => to_unsigned(28, 10), 1181 => to_unsigned(399, 10), 1182 => to_unsigned(706, 10), 1183 => to_unsigned(36, 10), 1184 => to_unsigned(647, 10), 1185 => to_unsigned(977, 10), 1186 => to_unsigned(671, 10), 1187 => to_unsigned(171, 10), 1188 => to_unsigned(41, 10), 1189 => to_unsigned(463, 10), 1190 => to_unsigned(796, 10), 1191 => to_unsigned(382, 10), 1192 => to_unsigned(182, 10), 1193 => to_unsigned(820, 10), 1194 => to_unsigned(118, 10), 1195 => to_unsigned(682, 10), 1196 => to_unsigned(760, 10), 1197 => to_unsigned(415, 10), 1198 => to_unsigned(86, 10), 1199 => to_unsigned(569, 10), 1200 => to_unsigned(498, 10), 1201 => to_unsigned(23, 10), 1202 => to_unsigned(124, 10), 1203 => to_unsigned(836, 10), 1204 => to_unsigned(576, 10), 1205 => to_unsigned(913, 10), 1206 => to_unsigned(198, 10), 1207 => to_unsigned(68, 10), 1208 => to_unsigned(203, 10), 1209 => to_unsigned(992, 10), 1210 => to_unsigned(208, 10), 1211 => to_unsigned(898, 10), 1212 => to_unsigned(506, 10), 1213 => to_unsigned(714, 10), 1214 => to_unsigned(423, 10), 1215 => to_unsigned(510, 10), 1216 => to_unsigned(166, 10), 1217 => to_unsigned(438, 10), 1218 => to_unsigned(764, 10), 1219 => to_unsigned(615, 10), 1220 => to_unsigned(1021, 10), 1221 => to_unsigned(247, 10), 1222 => to_unsigned(128, 10), 1223 => to_unsigned(777, 10), 1224 => to_unsigned(587, 10), 1225 => to_unsigned(428, 10), 1226 => to_unsigned(52, 10), 1227 => to_unsigned(209, 10), 1228 => to_unsigned(356, 10), 1229 => to_unsigned(361, 10), 1230 => to_unsigned(687, 10), 1231 => to_unsigned(709, 10), 1232 => to_unsigned(489, 10), 1233 => to_unsigned(560, 10), 1234 => to_unsigned(422, 10), 1235 => to_unsigned(36, 10), 1236 => to_unsigned(388, 10), 1237 => to_unsigned(763, 10), 1238 => to_unsigned(1009, 10), 1239 => to_unsigned(203, 10), 1240 => to_unsigned(39, 10), 1241 => to_unsigned(221, 10), 1242 => to_unsigned(747, 10), 1243 => to_unsigned(190, 10), 1244 => to_unsigned(685, 10), 1245 => to_unsigned(459, 10), 1246 => to_unsigned(810, 10), 1247 => to_unsigned(160, 10), 1248 => to_unsigned(897, 10), 1249 => to_unsigned(748, 10), 1250 => to_unsigned(175, 10), 1251 => to_unsigned(674, 10), 1252 => to_unsigned(298, 10), 1253 => to_unsigned(298, 10), 1254 => to_unsigned(364, 10), 1255 => to_unsigned(202, 10), 1256 => to_unsigned(426, 10), 1257 => to_unsigned(764, 10), 1258 => to_unsigned(744, 10), 1259 => to_unsigned(558, 10), 1260 => to_unsigned(999, 10), 1261 => to_unsigned(463, 10), 1262 => to_unsigned(621, 10), 1263 => to_unsigned(730, 10), 1264 => to_unsigned(617, 10), 1265 => to_unsigned(552, 10), 1266 => to_unsigned(620, 10), 1267 => to_unsigned(368, 10), 1268 => to_unsigned(848, 10), 1269 => to_unsigned(427, 10), 1270 => to_unsigned(860, 10), 1271 => to_unsigned(448, 10), 1272 => to_unsigned(575, 10), 1273 => to_unsigned(44, 10), 1274 => to_unsigned(893, 10), 1275 => to_unsigned(642, 10), 1276 => to_unsigned(534, 10), 1277 => to_unsigned(380, 10), 1278 => to_unsigned(920, 10), 1279 => to_unsigned(940, 10), 1280 => to_unsigned(851, 10), 1281 => to_unsigned(734, 10), 1282 => to_unsigned(973, 10), 1283 => to_unsigned(391, 10), 1284 => to_unsigned(211, 10), 1285 => to_unsigned(227, 10), 1286 => to_unsigned(309, 10), 1287 => to_unsigned(501, 10), 1288 => to_unsigned(318, 10), 1289 => to_unsigned(413, 10), 1290 => to_unsigned(724, 10), 1291 => to_unsigned(520, 10), 1292 => to_unsigned(970, 10), 1293 => to_unsigned(809, 10), 1294 => to_unsigned(930, 10), 1295 => to_unsigned(174, 10), 1296 => to_unsigned(957, 10), 1297 => to_unsigned(715, 10), 1298 => to_unsigned(253, 10), 1299 => to_unsigned(712, 10), 1300 => to_unsigned(629, 10), 1301 => to_unsigned(311, 10), 1302 => to_unsigned(981, 10), 1303 => to_unsigned(756, 10), 1304 => to_unsigned(580, 10), 1305 => to_unsigned(303, 10), 1306 => to_unsigned(519, 10), 1307 => to_unsigned(248, 10), 1308 => to_unsigned(312, 10), 1309 => to_unsigned(85, 10), 1310 => to_unsigned(86, 10), 1311 => to_unsigned(326, 10), 1312 => to_unsigned(19, 10), 1313 => to_unsigned(683, 10), 1314 => to_unsigned(326, 10), 1315 => to_unsigned(352, 10), 1316 => to_unsigned(507, 10), 1317 => to_unsigned(357, 10), 1318 => to_unsigned(342, 10), 1319 => to_unsigned(361, 10), 1320 => to_unsigned(789, 10), 1321 => to_unsigned(756, 10), 1322 => to_unsigned(139, 10), 1323 => to_unsigned(171, 10), 1324 => to_unsigned(67, 10), 1325 => to_unsigned(736, 10), 1326 => to_unsigned(925, 10), 1327 => to_unsigned(917, 10), 1328 => to_unsigned(209, 10), 1329 => to_unsigned(325, 10), 1330 => to_unsigned(751, 10), 1331 => to_unsigned(475, 10), 1332 => to_unsigned(257, 10), 1333 => to_unsigned(673, 10), 1334 => to_unsigned(424, 10), 1335 => to_unsigned(363, 10), 1336 => to_unsigned(103, 10), 1337 => to_unsigned(761, 10), 1338 => to_unsigned(683, 10), 1339 => to_unsigned(51, 10), 1340 => to_unsigned(997, 10), 1341 => to_unsigned(350, 10), 1342 => to_unsigned(466, 10), 1343 => to_unsigned(438, 10), 1344 => to_unsigned(975, 10), 1345 => to_unsigned(764, 10), 1346 => to_unsigned(307, 10), 1347 => to_unsigned(429, 10), 1348 => to_unsigned(232, 10), 1349 => to_unsigned(349, 10), 1350 => to_unsigned(132, 10), 1351 => to_unsigned(696, 10), 1352 => to_unsigned(432, 10), 1353 => to_unsigned(888, 10), 1354 => to_unsigned(490, 10), 1355 => to_unsigned(404, 10), 1356 => to_unsigned(784, 10), 1357 => to_unsigned(53, 10), 1358 => to_unsigned(981, 10), 1359 => to_unsigned(706, 10), 1360 => to_unsigned(404, 10), 1361 => to_unsigned(1005, 10), 1362 => to_unsigned(952, 10), 1363 => to_unsigned(408, 10), 1364 => to_unsigned(811, 10), 1365 => to_unsigned(340, 10), 1366 => to_unsigned(749, 10), 1367 => to_unsigned(703, 10), 1368 => to_unsigned(15, 10), 1369 => to_unsigned(353, 10), 1370 => to_unsigned(280, 10), 1371 => to_unsigned(344, 10), 1372 => to_unsigned(360, 10), 1373 => to_unsigned(603, 10), 1374 => to_unsigned(317, 10), 1375 => to_unsigned(643, 10), 1376 => to_unsigned(403, 10), 1377 => to_unsigned(652, 10), 1378 => to_unsigned(114, 10), 1379 => to_unsigned(300, 10), 1380 => to_unsigned(842, 10), 1381 => to_unsigned(393, 10), 1382 => to_unsigned(703, 10), 1383 => to_unsigned(988, 10), 1384 => to_unsigned(373, 10), 1385 => to_unsigned(686, 10), 1386 => to_unsigned(735, 10), 1387 => to_unsigned(471, 10), 1388 => to_unsigned(909, 10), 1389 => to_unsigned(581, 10), 1390 => to_unsigned(685, 10), 1391 => to_unsigned(1000, 10), 1392 => to_unsigned(135, 10), 1393 => to_unsigned(297, 10), 1394 => to_unsigned(622, 10), 1395 => to_unsigned(400, 10), 1396 => to_unsigned(178, 10), 1397 => to_unsigned(807, 10), 1398 => to_unsigned(35, 10), 1399 => to_unsigned(874, 10), 1400 => to_unsigned(284, 10), 1401 => to_unsigned(629, 10), 1402 => to_unsigned(81, 10), 1403 => to_unsigned(37, 10), 1404 => to_unsigned(513, 10), 1405 => to_unsigned(465, 10), 1406 => to_unsigned(286, 10), 1407 => to_unsigned(34, 10), 1408 => to_unsigned(884, 10), 1409 => to_unsigned(3, 10), 1410 => to_unsigned(417, 10), 1411 => to_unsigned(171, 10), 1412 => to_unsigned(345, 10), 1413 => to_unsigned(513, 10), 1414 => to_unsigned(354, 10), 1415 => to_unsigned(440, 10), 1416 => to_unsigned(817, 10), 1417 => to_unsigned(103, 10), 1418 => to_unsigned(808, 10), 1419 => to_unsigned(82, 10), 1420 => to_unsigned(553, 10), 1421 => to_unsigned(310, 10), 1422 => to_unsigned(981, 10), 1423 => to_unsigned(687, 10), 1424 => to_unsigned(604, 10), 1425 => to_unsigned(895, 10), 1426 => to_unsigned(961, 10), 1427 => to_unsigned(809, 10), 1428 => to_unsigned(806, 10), 1429 => to_unsigned(396, 10), 1430 => to_unsigned(207, 10), 1431 => to_unsigned(924, 10), 1432 => to_unsigned(281, 10), 1433 => to_unsigned(251, 10), 1434 => to_unsigned(242, 10), 1435 => to_unsigned(53, 10), 1436 => to_unsigned(470, 10), 1437 => to_unsigned(703, 10), 1438 => to_unsigned(347, 10), 1439 => to_unsigned(77, 10), 1440 => to_unsigned(673, 10), 1441 => to_unsigned(462, 10), 1442 => to_unsigned(373, 10), 1443 => to_unsigned(904, 10), 1444 => to_unsigned(196, 10), 1445 => to_unsigned(46, 10), 1446 => to_unsigned(630, 10), 1447 => to_unsigned(853, 10), 1448 => to_unsigned(685, 10), 1449 => to_unsigned(476, 10), 1450 => to_unsigned(790, 10), 1451 => to_unsigned(270, 10), 1452 => to_unsigned(256, 10), 1453 => to_unsigned(434, 10), 1454 => to_unsigned(485, 10), 1455 => to_unsigned(182, 10), 1456 => to_unsigned(178, 10), 1457 => to_unsigned(905, 10), 1458 => to_unsigned(801, 10), 1459 => to_unsigned(244, 10), 1460 => to_unsigned(552, 10), 1461 => to_unsigned(680, 10), 1462 => to_unsigned(755, 10), 1463 => to_unsigned(903, 10), 1464 => to_unsigned(922, 10), 1465 => to_unsigned(669, 10), 1466 => to_unsigned(946, 10), 1467 => to_unsigned(185, 10), 1468 => to_unsigned(529, 10), 1469 => to_unsigned(638, 10), 1470 => to_unsigned(266, 10), 1471 => to_unsigned(299, 10), 1472 => to_unsigned(958, 10), 1473 => to_unsigned(225, 10), 1474 => to_unsigned(961, 10), 1475 => to_unsigned(742, 10), 1476 => to_unsigned(893, 10), 1477 => to_unsigned(787, 10), 1478 => to_unsigned(221, 10), 1479 => to_unsigned(390, 10), 1480 => to_unsigned(5, 10), 1481 => to_unsigned(196, 10), 1482 => to_unsigned(450, 10), 1483 => to_unsigned(759, 10), 1484 => to_unsigned(424, 10), 1485 => to_unsigned(488, 10), 1486 => to_unsigned(976, 10), 1487 => to_unsigned(839, 10), 1488 => to_unsigned(936, 10), 1489 => to_unsigned(792, 10), 1490 => to_unsigned(215, 10), 1491 => to_unsigned(692, 10), 1492 => to_unsigned(378, 10), 1493 => to_unsigned(662, 10), 1494 => to_unsigned(553, 10), 1495 => to_unsigned(774, 10), 1496 => to_unsigned(120, 10), 1497 => to_unsigned(206, 10), 1498 => to_unsigned(563, 10), 1499 => to_unsigned(679, 10), 1500 => to_unsigned(1023, 10), 1501 => to_unsigned(536, 10), 1502 => to_unsigned(31, 10), 1503 => to_unsigned(660, 10), 1504 => to_unsigned(658, 10), 1505 => to_unsigned(803, 10), 1506 => to_unsigned(480, 10), 1507 => to_unsigned(724, 10), 1508 => to_unsigned(88, 10), 1509 => to_unsigned(480, 10), 1510 => to_unsigned(603, 10), 1511 => to_unsigned(812, 10), 1512 => to_unsigned(1018, 10), 1513 => to_unsigned(868, 10), 1514 => to_unsigned(466, 10), 1515 => to_unsigned(150, 10), 1516 => to_unsigned(482, 10), 1517 => to_unsigned(927, 10), 1518 => to_unsigned(690, 10), 1519 => to_unsigned(786, 10), 1520 => to_unsigned(508, 10), 1521 => to_unsigned(78, 10), 1522 => to_unsigned(519, 10), 1523 => to_unsigned(523, 10), 1524 => to_unsigned(703, 10), 1525 => to_unsigned(714, 10), 1526 => to_unsigned(953, 10), 1527 => to_unsigned(314, 10), 1528 => to_unsigned(550, 10), 1529 => to_unsigned(169, 10), 1530 => to_unsigned(982, 10), 1531 => to_unsigned(960, 10), 1532 => to_unsigned(34, 10), 1533 => to_unsigned(209, 10), 1534 => to_unsigned(426, 10), 1535 => to_unsigned(948, 10), 1536 => to_unsigned(70, 10), 1537 => to_unsigned(131, 10), 1538 => to_unsigned(936, 10), 1539 => to_unsigned(891, 10), 1540 => to_unsigned(91, 10), 1541 => to_unsigned(972, 10), 1542 => to_unsigned(679, 10), 1543 => to_unsigned(213, 10), 1544 => to_unsigned(793, 10), 1545 => to_unsigned(768, 10), 1546 => to_unsigned(107, 10), 1547 => to_unsigned(930, 10), 1548 => to_unsigned(381, 10), 1549 => to_unsigned(961, 10), 1550 => to_unsigned(880, 10), 1551 => to_unsigned(555, 10), 1552 => to_unsigned(677, 10), 1553 => to_unsigned(1006, 10), 1554 => to_unsigned(107, 10), 1555 => to_unsigned(473, 10), 1556 => to_unsigned(983, 10), 1557 => to_unsigned(810, 10), 1558 => to_unsigned(499, 10), 1559 => to_unsigned(708, 10), 1560 => to_unsigned(692, 10), 1561 => to_unsigned(455, 10), 1562 => to_unsigned(93, 10), 1563 => to_unsigned(1, 10), 1564 => to_unsigned(23, 10), 1565 => to_unsigned(215, 10), 1566 => to_unsigned(344, 10), 1567 => to_unsigned(345, 10), 1568 => to_unsigned(325, 10), 1569 => to_unsigned(918, 10), 1570 => to_unsigned(1009, 10), 1571 => to_unsigned(80, 10), 1572 => to_unsigned(351, 10), 1573 => to_unsigned(240, 10), 1574 => to_unsigned(704, 10), 1575 => to_unsigned(498, 10), 1576 => to_unsigned(963, 10), 1577 => to_unsigned(353, 10), 1578 => to_unsigned(799, 10), 1579 => to_unsigned(454, 10), 1580 => to_unsigned(52, 10), 1581 => to_unsigned(576, 10), 1582 => to_unsigned(776, 10), 1583 => to_unsigned(792, 10), 1584 => to_unsigned(70, 10), 1585 => to_unsigned(331, 10), 1586 => to_unsigned(964, 10), 1587 => to_unsigned(830, 10), 1588 => to_unsigned(245, 10), 1589 => to_unsigned(101, 10), 1590 => to_unsigned(839, 10), 1591 => to_unsigned(503, 10), 1592 => to_unsigned(537, 10), 1593 => to_unsigned(435, 10), 1594 => to_unsigned(810, 10), 1595 => to_unsigned(645, 10), 1596 => to_unsigned(933, 10), 1597 => to_unsigned(900, 10), 1598 => to_unsigned(764, 10), 1599 => to_unsigned(767, 10), 1600 => to_unsigned(958, 10), 1601 => to_unsigned(810, 10), 1602 => to_unsigned(1017, 10), 1603 => to_unsigned(12, 10), 1604 => to_unsigned(784, 10), 1605 => to_unsigned(185, 10), 1606 => to_unsigned(581, 10), 1607 => to_unsigned(13, 10), 1608 => to_unsigned(779, 10), 1609 => to_unsigned(982, 10), 1610 => to_unsigned(362, 10), 1611 => to_unsigned(295, 10), 1612 => to_unsigned(256, 10), 1613 => to_unsigned(408, 10), 1614 => to_unsigned(880, 10), 1615 => to_unsigned(667, 10), 1616 => to_unsigned(887, 10), 1617 => to_unsigned(670, 10), 1618 => to_unsigned(216, 10), 1619 => to_unsigned(988, 10), 1620 => to_unsigned(408, 10), 1621 => to_unsigned(767, 10), 1622 => to_unsigned(894, 10), 1623 => to_unsigned(94, 10), 1624 => to_unsigned(633, 10), 1625 => to_unsigned(948, 10), 1626 => to_unsigned(366, 10), 1627 => to_unsigned(672, 10), 1628 => to_unsigned(958, 10), 1629 => to_unsigned(829, 10), 1630 => to_unsigned(494, 10), 1631 => to_unsigned(995, 10), 1632 => to_unsigned(86, 10), 1633 => to_unsigned(815, 10), 1634 => to_unsigned(648, 10), 1635 => to_unsigned(515, 10), 1636 => to_unsigned(612, 10), 1637 => to_unsigned(692, 10), 1638 => to_unsigned(206, 10), 1639 => to_unsigned(828, 10), 1640 => to_unsigned(740, 10), 1641 => to_unsigned(827, 10), 1642 => to_unsigned(465, 10), 1643 => to_unsigned(955, 10), 1644 => to_unsigned(979, 10), 1645 => to_unsigned(344, 10), 1646 => to_unsigned(88, 10), 1647 => to_unsigned(99, 10), 1648 => to_unsigned(242, 10), 1649 => to_unsigned(833, 10), 1650 => to_unsigned(204, 10), 1651 => to_unsigned(340, 10), 1652 => to_unsigned(7, 10), 1653 => to_unsigned(86, 10), 1654 => to_unsigned(812, 10), 1655 => to_unsigned(760, 10), 1656 => to_unsigned(207, 10), 1657 => to_unsigned(32, 10), 1658 => to_unsigned(33, 10), 1659 => to_unsigned(333, 10), 1660 => to_unsigned(641, 10), 1661 => to_unsigned(515, 10), 1662 => to_unsigned(423, 10), 1663 => to_unsigned(248, 10), 1664 => to_unsigned(446, 10), 1665 => to_unsigned(62, 10), 1666 => to_unsigned(612, 10), 1667 => to_unsigned(998, 10), 1668 => to_unsigned(283, 10), 1669 => to_unsigned(954, 10), 1670 => to_unsigned(610, 10), 1671 => to_unsigned(365, 10), 1672 => to_unsigned(230, 10), 1673 => to_unsigned(431, 10), 1674 => to_unsigned(921, 10), 1675 => to_unsigned(336, 10), 1676 => to_unsigned(240, 10), 1677 => to_unsigned(114, 10), 1678 => to_unsigned(511, 10), 1679 => to_unsigned(201, 10), 1680 => to_unsigned(665, 10), 1681 => to_unsigned(448, 10), 1682 => to_unsigned(783, 10), 1683 => to_unsigned(501, 10), 1684 => to_unsigned(80, 10), 1685 => to_unsigned(746, 10), 1686 => to_unsigned(509, 10), 1687 => to_unsigned(612, 10), 1688 => to_unsigned(7, 10), 1689 => to_unsigned(407, 10), 1690 => to_unsigned(241, 10), 1691 => to_unsigned(296, 10), 1692 => to_unsigned(550, 10), 1693 => to_unsigned(877, 10), 1694 => to_unsigned(549, 10), 1695 => to_unsigned(625, 10), 1696 => to_unsigned(613, 10), 1697 => to_unsigned(452, 10), 1698 => to_unsigned(226, 10), 1699 => to_unsigned(854, 10), 1700 => to_unsigned(956, 10), 1701 => to_unsigned(250, 10), 1702 => to_unsigned(305, 10), 1703 => to_unsigned(542, 10), 1704 => to_unsigned(763, 10), 1705 => to_unsigned(737, 10), 1706 => to_unsigned(475, 10), 1707 => to_unsigned(327, 10), 1708 => to_unsigned(717, 10), 1709 => to_unsigned(729, 10), 1710 => to_unsigned(421, 10), 1711 => to_unsigned(927, 10), 1712 => to_unsigned(740, 10), 1713 => to_unsigned(250, 10), 1714 => to_unsigned(945, 10), 1715 => to_unsigned(943, 10), 1716 => to_unsigned(309, 10), 1717 => to_unsigned(615, 10), 1718 => to_unsigned(648, 10), 1719 => to_unsigned(786, 10), 1720 => to_unsigned(980, 10), 1721 => to_unsigned(25, 10), 1722 => to_unsigned(423, 10), 1723 => to_unsigned(989, 10), 1724 => to_unsigned(258, 10), 1725 => to_unsigned(488, 10), 1726 => to_unsigned(690, 10), 1727 => to_unsigned(209, 10), 1728 => to_unsigned(616, 10), 1729 => to_unsigned(615, 10), 1730 => to_unsigned(609, 10), 1731 => to_unsigned(3, 10), 1732 => to_unsigned(26, 10), 1733 => to_unsigned(437, 10), 1734 => to_unsigned(111, 10), 1735 => to_unsigned(984, 10), 1736 => to_unsigned(191, 10), 1737 => to_unsigned(255, 10), 1738 => to_unsigned(1023, 10), 1739 => to_unsigned(369, 10), 1740 => to_unsigned(478, 10), 1741 => to_unsigned(627, 10), 1742 => to_unsigned(441, 10), 1743 => to_unsigned(65, 10), 1744 => to_unsigned(618, 10), 1745 => to_unsigned(850, 10), 1746 => to_unsigned(327, 10), 1747 => to_unsigned(683, 10), 1748 => to_unsigned(581, 10), 1749 => to_unsigned(826, 10), 1750 => to_unsigned(424, 10), 1751 => to_unsigned(613, 10), 1752 => to_unsigned(659, 10), 1753 => to_unsigned(34, 10), 1754 => to_unsigned(213, 10), 1755 => to_unsigned(996, 10), 1756 => to_unsigned(88, 10), 1757 => to_unsigned(606, 10), 1758 => to_unsigned(705, 10), 1759 => to_unsigned(640, 10), 1760 => to_unsigned(216, 10), 1761 => to_unsigned(365, 10), 1762 => to_unsigned(815, 10), 1763 => to_unsigned(888, 10), 1764 => to_unsigned(516, 10), 1765 => to_unsigned(64, 10), 1766 => to_unsigned(420, 10), 1767 => to_unsigned(572, 10), 1768 => to_unsigned(690, 10), 1769 => to_unsigned(183, 10), 1770 => to_unsigned(468, 10), 1771 => to_unsigned(836, 10), 1772 => to_unsigned(773, 10), 1773 => to_unsigned(701, 10), 1774 => to_unsigned(462, 10), 1775 => to_unsigned(22, 10), 1776 => to_unsigned(975, 10), 1777 => to_unsigned(83, 10), 1778 => to_unsigned(844, 10), 1779 => to_unsigned(317, 10), 1780 => to_unsigned(167, 10), 1781 => to_unsigned(800, 10), 1782 => to_unsigned(697, 10), 1783 => to_unsigned(30, 10), 1784 => to_unsigned(340, 10), 1785 => to_unsigned(404, 10), 1786 => to_unsigned(442, 10), 1787 => to_unsigned(581, 10), 1788 => to_unsigned(458, 10), 1789 => to_unsigned(344, 10), 1790 => to_unsigned(203, 10), 1791 => to_unsigned(917, 10), 1792 => to_unsigned(252, 10), 1793 => to_unsigned(326, 10), 1794 => to_unsigned(705, 10), 1795 => to_unsigned(436, 10), 1796 => to_unsigned(525, 10), 1797 => to_unsigned(847, 10), 1798 => to_unsigned(623, 10), 1799 => to_unsigned(811, 10), 1800 => to_unsigned(981, 10), 1801 => to_unsigned(835, 10), 1802 => to_unsigned(221, 10), 1803 => to_unsigned(9, 10), 1804 => to_unsigned(566, 10), 1805 => to_unsigned(856, 10), 1806 => to_unsigned(695, 10), 1807 => to_unsigned(484, 10), 1808 => to_unsigned(1020, 10), 1809 => to_unsigned(634, 10), 1810 => to_unsigned(823, 10), 1811 => to_unsigned(184, 10), 1812 => to_unsigned(305, 10), 1813 => to_unsigned(276, 10), 1814 => to_unsigned(421, 10), 1815 => to_unsigned(949, 10), 1816 => to_unsigned(829, 10), 1817 => to_unsigned(1006, 10), 1818 => to_unsigned(467, 10), 1819 => to_unsigned(808, 10), 1820 => to_unsigned(382, 10), 1821 => to_unsigned(579, 10), 1822 => to_unsigned(293, 10), 1823 => to_unsigned(643, 10), 1824 => to_unsigned(468, 10), 1825 => to_unsigned(934, 10), 1826 => to_unsigned(734, 10), 1827 => to_unsigned(801, 10), 1828 => to_unsigned(89, 10), 1829 => to_unsigned(169, 10), 1830 => to_unsigned(748, 10), 1831 => to_unsigned(503, 10), 1832 => to_unsigned(22, 10), 1833 => to_unsigned(485, 10), 1834 => to_unsigned(322, 10), 1835 => to_unsigned(569, 10), 1836 => to_unsigned(667, 10), 1837 => to_unsigned(494, 10), 1838 => to_unsigned(243, 10), 1839 => to_unsigned(229, 10), 1840 => to_unsigned(58, 10), 1841 => to_unsigned(120, 10), 1842 => to_unsigned(156, 10), 1843 => to_unsigned(956, 10), 1844 => to_unsigned(227, 10), 1845 => to_unsigned(815, 10), 1846 => to_unsigned(289, 10), 1847 => to_unsigned(921, 10), 1848 => to_unsigned(630, 10), 1849 => to_unsigned(458, 10), 1850 => to_unsigned(231, 10), 1851 => to_unsigned(456, 10), 1852 => to_unsigned(465, 10), 1853 => to_unsigned(217, 10), 1854 => to_unsigned(775, 10), 1855 => to_unsigned(947, 10), 1856 => to_unsigned(285, 10), 1857 => to_unsigned(167, 10), 1858 => to_unsigned(425, 10), 1859 => to_unsigned(788, 10), 1860 => to_unsigned(289, 10), 1861 => to_unsigned(625, 10), 1862 => to_unsigned(120, 10), 1863 => to_unsigned(252, 10), 1864 => to_unsigned(522, 10), 1865 => to_unsigned(588, 10), 1866 => to_unsigned(559, 10), 1867 => to_unsigned(386, 10), 1868 => to_unsigned(736, 10), 1869 => to_unsigned(984, 10), 1870 => to_unsigned(309, 10), 1871 => to_unsigned(325, 10), 1872 => to_unsigned(403, 10), 1873 => to_unsigned(384, 10), 1874 => to_unsigned(401, 10), 1875 => to_unsigned(471, 10), 1876 => to_unsigned(622, 10), 1877 => to_unsigned(980, 10), 1878 => to_unsigned(58, 10), 1879 => to_unsigned(996, 10), 1880 => to_unsigned(676, 10), 1881 => to_unsigned(396, 10), 1882 => to_unsigned(684, 10), 1883 => to_unsigned(740, 10), 1884 => to_unsigned(847, 10), 1885 => to_unsigned(421, 10), 1886 => to_unsigned(118, 10), 1887 => to_unsigned(408, 10), 1888 => to_unsigned(685, 10), 1889 => to_unsigned(180, 10), 1890 => to_unsigned(852, 10), 1891 => to_unsigned(890, 10), 1892 => to_unsigned(700, 10), 1893 => to_unsigned(391, 10), 1894 => to_unsigned(878, 10), 1895 => to_unsigned(23, 10), 1896 => to_unsigned(788, 10), 1897 => to_unsigned(69, 10), 1898 => to_unsigned(263, 10), 1899 => to_unsigned(804, 10), 1900 => to_unsigned(111, 10), 1901 => to_unsigned(649, 10), 1902 => to_unsigned(197, 10), 1903 => to_unsigned(281, 10), 1904 => to_unsigned(545, 10), 1905 => to_unsigned(468, 10), 1906 => to_unsigned(576, 10), 1907 => to_unsigned(161, 10), 1908 => to_unsigned(83, 10), 1909 => to_unsigned(457, 10), 1910 => to_unsigned(258, 10), 1911 => to_unsigned(528, 10), 1912 => to_unsigned(126, 10), 1913 => to_unsigned(87, 10), 1914 => to_unsigned(829, 10), 1915 => to_unsigned(826, 10), 1916 => to_unsigned(626, 10), 1917 => to_unsigned(25, 10), 1918 => to_unsigned(122, 10), 1919 => to_unsigned(938, 10), 1920 => to_unsigned(720, 10), 1921 => to_unsigned(913, 10), 1922 => to_unsigned(40, 10), 1923 => to_unsigned(316, 10), 1924 => to_unsigned(337, 10), 1925 => to_unsigned(506, 10), 1926 => to_unsigned(253, 10), 1927 => to_unsigned(497, 10), 1928 => to_unsigned(741, 10), 1929 => to_unsigned(425, 10), 1930 => to_unsigned(422, 10), 1931 => to_unsigned(204, 10), 1932 => to_unsigned(198, 10), 1933 => to_unsigned(367, 10), 1934 => to_unsigned(280, 10), 1935 => to_unsigned(289, 10), 1936 => to_unsigned(462, 10), 1937 => to_unsigned(197, 10), 1938 => to_unsigned(9, 10), 1939 => to_unsigned(37, 10), 1940 => to_unsigned(358, 10), 1941 => to_unsigned(907, 10), 1942 => to_unsigned(921, 10), 1943 => to_unsigned(784, 10), 1944 => to_unsigned(83, 10), 1945 => to_unsigned(829, 10), 1946 => to_unsigned(378, 10), 1947 => to_unsigned(919, 10), 1948 => to_unsigned(434, 10), 1949 => to_unsigned(633, 10), 1950 => to_unsigned(880, 10), 1951 => to_unsigned(521, 10), 1952 => to_unsigned(810, 10), 1953 => to_unsigned(425, 10), 1954 => to_unsigned(745, 10), 1955 => to_unsigned(999, 10), 1956 => to_unsigned(26, 10), 1957 => to_unsigned(375, 10), 1958 => to_unsigned(630, 10), 1959 => to_unsigned(810, 10), 1960 => to_unsigned(62, 10), 1961 => to_unsigned(779, 10), 1962 => to_unsigned(967, 10), 1963 => to_unsigned(987, 10), 1964 => to_unsigned(160, 10), 1965 => to_unsigned(637, 10), 1966 => to_unsigned(798, 10), 1967 => to_unsigned(854, 10), 1968 => to_unsigned(285, 10), 1969 => to_unsigned(32, 10), 1970 => to_unsigned(450, 10), 1971 => to_unsigned(406, 10), 1972 => to_unsigned(175, 10), 1973 => to_unsigned(40, 10), 1974 => to_unsigned(239, 10), 1975 => to_unsigned(408, 10), 1976 => to_unsigned(374, 10), 1977 => to_unsigned(1011, 10), 1978 => to_unsigned(654, 10), 1979 => to_unsigned(514, 10), 1980 => to_unsigned(195, 10), 1981 => to_unsigned(545, 10), 1982 => to_unsigned(810, 10), 1983 => to_unsigned(292, 10), 1984 => to_unsigned(128, 10), 1985 => to_unsigned(920, 10), 1986 => to_unsigned(50, 10), 1987 => to_unsigned(294, 10), 1988 => to_unsigned(823, 10), 1989 => to_unsigned(268, 10), 1990 => to_unsigned(637, 10), 1991 => to_unsigned(271, 10), 1992 => to_unsigned(26, 10), 1993 => to_unsigned(919, 10), 1994 => to_unsigned(696, 10), 1995 => to_unsigned(989, 10), 1996 => to_unsigned(784, 10), 1997 => to_unsigned(338, 10), 1998 => to_unsigned(941, 10), 1999 => to_unsigned(673, 10), 2000 => to_unsigned(246, 10), 2001 => to_unsigned(387, 10), 2002 => to_unsigned(570, 10), 2003 => to_unsigned(870, 10), 2004 => to_unsigned(71, 10), 2005 => to_unsigned(57, 10), 2006 => to_unsigned(660, 10), 2007 => to_unsigned(368, 10), 2008 => to_unsigned(472, 10), 2009 => to_unsigned(834, 10), 2010 => to_unsigned(510, 10), 2011 => to_unsigned(60, 10), 2012 => to_unsigned(522, 10), 2013 => to_unsigned(563, 10), 2014 => to_unsigned(866, 10), 2015 => to_unsigned(728, 10), 2016 => to_unsigned(256, 10), 2017 => to_unsigned(70, 10), 2018 => to_unsigned(781, 10), 2019 => to_unsigned(742, 10), 2020 => to_unsigned(25, 10), 2021 => to_unsigned(91, 10), 2022 => to_unsigned(303, 10), 2023 => to_unsigned(325, 10), 2024 => to_unsigned(493, 10), 2025 => to_unsigned(1021, 10), 2026 => to_unsigned(617, 10), 2027 => to_unsigned(23, 10), 2028 => to_unsigned(947, 10), 2029 => to_unsigned(438, 10), 2030 => to_unsigned(280, 10), 2031 => to_unsigned(461, 10), 2032 => to_unsigned(789, 10), 2033 => to_unsigned(525, 10), 2034 => to_unsigned(66, 10), 2035 => to_unsigned(504, 10), 2036 => to_unsigned(681, 10), 2037 => to_unsigned(641, 10), 2038 => to_unsigned(58, 10), 2039 => to_unsigned(1005, 10), 2040 => to_unsigned(564, 10), 2041 => to_unsigned(896, 10), 2042 => to_unsigned(441, 10), 2043 => to_unsigned(894, 10), 2044 => to_unsigned(1020, 10), 2045 => to_unsigned(526, 10), 2046 => to_unsigned(356, 10), 2047 => to_unsigned(135, 10)),
            3 => (0 => to_unsigned(816, 10), 1 => to_unsigned(73, 10), 2 => to_unsigned(108, 10), 3 => to_unsigned(561, 10), 4 => to_unsigned(516, 10), 5 => to_unsigned(16, 10), 6 => to_unsigned(144, 10), 7 => to_unsigned(249, 10), 8 => to_unsigned(831, 10), 9 => to_unsigned(912, 10), 10 => to_unsigned(451, 10), 11 => to_unsigned(872, 10), 12 => to_unsigned(182, 10), 13 => to_unsigned(258, 10), 14 => to_unsigned(544, 10), 15 => to_unsigned(697, 10), 16 => to_unsigned(326, 10), 17 => to_unsigned(981, 10), 18 => to_unsigned(668, 10), 19 => to_unsigned(790, 10), 20 => to_unsigned(667, 10), 21 => to_unsigned(889, 10), 22 => to_unsigned(177, 10), 23 => to_unsigned(894, 10), 24 => to_unsigned(772, 10), 25 => to_unsigned(772, 10), 26 => to_unsigned(991, 10), 27 => to_unsigned(962, 10), 28 => to_unsigned(217, 10), 29 => to_unsigned(734, 10), 30 => to_unsigned(331, 10), 31 => to_unsigned(714, 10), 32 => to_unsigned(194, 10), 33 => to_unsigned(331, 10), 34 => to_unsigned(588, 10), 35 => to_unsigned(468, 10), 36 => to_unsigned(649, 10), 37 => to_unsigned(762, 10), 38 => to_unsigned(35, 10), 39 => to_unsigned(435, 10), 40 => to_unsigned(646, 10), 41 => to_unsigned(510, 10), 42 => to_unsigned(543, 10), 43 => to_unsigned(283, 10), 44 => to_unsigned(10, 10), 45 => to_unsigned(688, 10), 46 => to_unsigned(968, 10), 47 => to_unsigned(217, 10), 48 => to_unsigned(613, 10), 49 => to_unsigned(335, 10), 50 => to_unsigned(538, 10), 51 => to_unsigned(837, 10), 52 => to_unsigned(210, 10), 53 => to_unsigned(960, 10), 54 => to_unsigned(932, 10), 55 => to_unsigned(32, 10), 56 => to_unsigned(37, 10), 57 => to_unsigned(594, 10), 58 => to_unsigned(77, 10), 59 => to_unsigned(723, 10), 60 => to_unsigned(834, 10), 61 => to_unsigned(239, 10), 62 => to_unsigned(761, 10), 63 => to_unsigned(168, 10), 64 => to_unsigned(233, 10), 65 => to_unsigned(128, 10), 66 => to_unsigned(166, 10), 67 => to_unsigned(320, 10), 68 => to_unsigned(905, 10), 69 => to_unsigned(830, 10), 70 => to_unsigned(945, 10), 71 => to_unsigned(515, 10), 72 => to_unsigned(133, 10), 73 => to_unsigned(849, 10), 74 => to_unsigned(764, 10), 75 => to_unsigned(274, 10), 76 => to_unsigned(813, 10), 77 => to_unsigned(715, 10), 78 => to_unsigned(576, 10), 79 => to_unsigned(629, 10), 80 => to_unsigned(294, 10), 81 => to_unsigned(108, 10), 82 => to_unsigned(169, 10), 83 => to_unsigned(529, 10), 84 => to_unsigned(684, 10), 85 => to_unsigned(658, 10), 86 => to_unsigned(447, 10), 87 => to_unsigned(390, 10), 88 => to_unsigned(975, 10), 89 => to_unsigned(822, 10), 90 => to_unsigned(700, 10), 91 => to_unsigned(423, 10), 92 => to_unsigned(384, 10), 93 => to_unsigned(293, 10), 94 => to_unsigned(548, 10), 95 => to_unsigned(135, 10), 96 => to_unsigned(557, 10), 97 => to_unsigned(511, 10), 98 => to_unsigned(907, 10), 99 => to_unsigned(644, 10), 100 => to_unsigned(710, 10), 101 => to_unsigned(550, 10), 102 => to_unsigned(892, 10), 103 => to_unsigned(808, 10), 104 => to_unsigned(830, 10), 105 => to_unsigned(838, 10), 106 => to_unsigned(976, 10), 107 => to_unsigned(674, 10), 108 => to_unsigned(848, 10), 109 => to_unsigned(736, 10), 110 => to_unsigned(1016, 10), 111 => to_unsigned(412, 10), 112 => to_unsigned(996, 10), 113 => to_unsigned(928, 10), 114 => to_unsigned(817, 10), 115 => to_unsigned(1008, 10), 116 => to_unsigned(264, 10), 117 => to_unsigned(789, 10), 118 => to_unsigned(50, 10), 119 => to_unsigned(408, 10), 120 => to_unsigned(400, 10), 121 => to_unsigned(85, 10), 122 => to_unsigned(266, 10), 123 => to_unsigned(160, 10), 124 => to_unsigned(392, 10), 125 => to_unsigned(187, 10), 126 => to_unsigned(485, 10), 127 => to_unsigned(454, 10), 128 => to_unsigned(474, 10), 129 => to_unsigned(106, 10), 130 => to_unsigned(731, 10), 131 => to_unsigned(762, 10), 132 => to_unsigned(45, 10), 133 => to_unsigned(985, 10), 134 => to_unsigned(660, 10), 135 => to_unsigned(468, 10), 136 => to_unsigned(717, 10), 137 => to_unsigned(162, 10), 138 => to_unsigned(260, 10), 139 => to_unsigned(560, 10), 140 => to_unsigned(974, 10), 141 => to_unsigned(536, 10), 142 => to_unsigned(705, 10), 143 => to_unsigned(615, 10), 144 => to_unsigned(811, 10), 145 => to_unsigned(205, 10), 146 => to_unsigned(228, 10), 147 => to_unsigned(481, 10), 148 => to_unsigned(204, 10), 149 => to_unsigned(528, 10), 150 => to_unsigned(57, 10), 151 => to_unsigned(517, 10), 152 => to_unsigned(993, 10), 153 => to_unsigned(379, 10), 154 => to_unsigned(735, 10), 155 => to_unsigned(8, 10), 156 => to_unsigned(33, 10), 157 => to_unsigned(310, 10), 158 => to_unsigned(320, 10), 159 => to_unsigned(416, 10), 160 => to_unsigned(479, 10), 161 => to_unsigned(770, 10), 162 => to_unsigned(490, 10), 163 => to_unsigned(155, 10), 164 => to_unsigned(720, 10), 165 => to_unsigned(87, 10), 166 => to_unsigned(834, 10), 167 => to_unsigned(967, 10), 168 => to_unsigned(741, 10), 169 => to_unsigned(45, 10), 170 => to_unsigned(660, 10), 171 => to_unsigned(704, 10), 172 => to_unsigned(647, 10), 173 => to_unsigned(473, 10), 174 => to_unsigned(792, 10), 175 => to_unsigned(193, 10), 176 => to_unsigned(611, 10), 177 => to_unsigned(318, 10), 178 => to_unsigned(94, 10), 179 => to_unsigned(418, 10), 180 => to_unsigned(220, 10), 181 => to_unsigned(226, 10), 182 => to_unsigned(917, 10), 183 => to_unsigned(343, 10), 184 => to_unsigned(913, 10), 185 => to_unsigned(325, 10), 186 => to_unsigned(895, 10), 187 => to_unsigned(771, 10), 188 => to_unsigned(345, 10), 189 => to_unsigned(149, 10), 190 => to_unsigned(699, 10), 191 => to_unsigned(646, 10), 192 => to_unsigned(701, 10), 193 => to_unsigned(723, 10), 194 => to_unsigned(22, 10), 195 => to_unsigned(535, 10), 196 => to_unsigned(85, 10), 197 => to_unsigned(76, 10), 198 => to_unsigned(662, 10), 199 => to_unsigned(60, 10), 200 => to_unsigned(906, 10), 201 => to_unsigned(718, 10), 202 => to_unsigned(1004, 10), 203 => to_unsigned(185, 10), 204 => to_unsigned(41, 10), 205 => to_unsigned(581, 10), 206 => to_unsigned(679, 10), 207 => to_unsigned(757, 10), 208 => to_unsigned(883, 10), 209 => to_unsigned(458, 10), 210 => to_unsigned(445, 10), 211 => to_unsigned(346, 10), 212 => to_unsigned(410, 10), 213 => to_unsigned(723, 10), 214 => to_unsigned(174, 10), 215 => to_unsigned(628, 10), 216 => to_unsigned(144, 10), 217 => to_unsigned(641, 10), 218 => to_unsigned(211, 10), 219 => to_unsigned(334, 10), 220 => to_unsigned(521, 10), 221 => to_unsigned(831, 10), 222 => to_unsigned(492, 10), 223 => to_unsigned(319, 10), 224 => to_unsigned(444, 10), 225 => to_unsigned(163, 10), 226 => to_unsigned(355, 10), 227 => to_unsigned(136, 10), 228 => to_unsigned(730, 10), 229 => to_unsigned(568, 10), 230 => to_unsigned(371, 10), 231 => to_unsigned(360, 10), 232 => to_unsigned(173, 10), 233 => to_unsigned(845, 10), 234 => to_unsigned(189, 10), 235 => to_unsigned(729, 10), 236 => to_unsigned(300, 10), 237 => to_unsigned(948, 10), 238 => to_unsigned(526, 10), 239 => to_unsigned(496, 10), 240 => to_unsigned(141, 10), 241 => to_unsigned(570, 10), 242 => to_unsigned(902, 10), 243 => to_unsigned(363, 10), 244 => to_unsigned(252, 10), 245 => to_unsigned(584, 10), 246 => to_unsigned(742, 10), 247 => to_unsigned(51, 10), 248 => to_unsigned(782, 10), 249 => to_unsigned(622, 10), 250 => to_unsigned(796, 10), 251 => to_unsigned(157, 10), 252 => to_unsigned(223, 10), 253 => to_unsigned(94, 10), 254 => to_unsigned(264, 10), 255 => to_unsigned(619, 10), 256 => to_unsigned(450, 10), 257 => to_unsigned(56, 10), 258 => to_unsigned(335, 10), 259 => to_unsigned(440, 10), 260 => to_unsigned(952, 10), 261 => to_unsigned(988, 10), 262 => to_unsigned(866, 10), 263 => to_unsigned(805, 10), 264 => to_unsigned(682, 10), 265 => to_unsigned(102, 10), 266 => to_unsigned(357, 10), 267 => to_unsigned(216, 10), 268 => to_unsigned(261, 10), 269 => to_unsigned(910, 10), 270 => to_unsigned(696, 10), 271 => to_unsigned(226, 10), 272 => to_unsigned(395, 10), 273 => to_unsigned(912, 10), 274 => to_unsigned(671, 10), 275 => to_unsigned(242, 10), 276 => to_unsigned(588, 10), 277 => to_unsigned(186, 10), 278 => to_unsigned(955, 10), 279 => to_unsigned(448, 10), 280 => to_unsigned(957, 10), 281 => to_unsigned(866, 10), 282 => to_unsigned(1017, 10), 283 => to_unsigned(576, 10), 284 => to_unsigned(632, 10), 285 => to_unsigned(57, 10), 286 => to_unsigned(656, 10), 287 => to_unsigned(895, 10), 288 => to_unsigned(644, 10), 289 => to_unsigned(356, 10), 290 => to_unsigned(515, 10), 291 => to_unsigned(389, 10), 292 => to_unsigned(734, 10), 293 => to_unsigned(251, 10), 294 => to_unsigned(50, 10), 295 => to_unsigned(383, 10), 296 => to_unsigned(170, 10), 297 => to_unsigned(724, 10), 298 => to_unsigned(432, 10), 299 => to_unsigned(813, 10), 300 => to_unsigned(271, 10), 301 => to_unsigned(229, 10), 302 => to_unsigned(233, 10), 303 => to_unsigned(117, 10), 304 => to_unsigned(732, 10), 305 => to_unsigned(603, 10), 306 => to_unsigned(183, 10), 307 => to_unsigned(187, 10), 308 => to_unsigned(507, 10), 309 => to_unsigned(493, 10), 310 => to_unsigned(183, 10), 311 => to_unsigned(893, 10), 312 => to_unsigned(673, 10), 313 => to_unsigned(267, 10), 314 => to_unsigned(639, 10), 315 => to_unsigned(987, 10), 316 => to_unsigned(802, 10), 317 => to_unsigned(472, 10), 318 => to_unsigned(269, 10), 319 => to_unsigned(391, 10), 320 => to_unsigned(408, 10), 321 => to_unsigned(705, 10), 322 => to_unsigned(99, 10), 323 => to_unsigned(594, 10), 324 => to_unsigned(366, 10), 325 => to_unsigned(296, 10), 326 => to_unsigned(695, 10), 327 => to_unsigned(577, 10), 328 => to_unsigned(234, 10), 329 => to_unsigned(283, 10), 330 => to_unsigned(911, 10), 331 => to_unsigned(143, 10), 332 => to_unsigned(297, 10), 333 => to_unsigned(973, 10), 334 => to_unsigned(518, 10), 335 => to_unsigned(638, 10), 336 => to_unsigned(250, 10), 337 => to_unsigned(224, 10), 338 => to_unsigned(476, 10), 339 => to_unsigned(824, 10), 340 => to_unsigned(180, 10), 341 => to_unsigned(646, 10), 342 => to_unsigned(334, 10), 343 => to_unsigned(415, 10), 344 => to_unsigned(390, 10), 345 => to_unsigned(545, 10), 346 => to_unsigned(383, 10), 347 => to_unsigned(186, 10), 348 => to_unsigned(762, 10), 349 => to_unsigned(894, 10), 350 => to_unsigned(46, 10), 351 => to_unsigned(639, 10), 352 => to_unsigned(538, 10), 353 => to_unsigned(51, 10), 354 => to_unsigned(160, 10), 355 => to_unsigned(700, 10), 356 => to_unsigned(763, 10), 357 => to_unsigned(814, 10), 358 => to_unsigned(95, 10), 359 => to_unsigned(647, 10), 360 => to_unsigned(689, 10), 361 => to_unsigned(807, 10), 362 => to_unsigned(193, 10), 363 => to_unsigned(261, 10), 364 => to_unsigned(613, 10), 365 => to_unsigned(667, 10), 366 => to_unsigned(934, 10), 367 => to_unsigned(557, 10), 368 => to_unsigned(663, 10), 369 => to_unsigned(268, 10), 370 => to_unsigned(649, 10), 371 => to_unsigned(157, 10), 372 => to_unsigned(157, 10), 373 => to_unsigned(13, 10), 374 => to_unsigned(599, 10), 375 => to_unsigned(792, 10), 376 => to_unsigned(649, 10), 377 => to_unsigned(68, 10), 378 => to_unsigned(421, 10), 379 => to_unsigned(440, 10), 380 => to_unsigned(715, 10), 381 => to_unsigned(342, 10), 382 => to_unsigned(188, 10), 383 => to_unsigned(664, 10), 384 => to_unsigned(613, 10), 385 => to_unsigned(104, 10), 386 => to_unsigned(488, 10), 387 => to_unsigned(180, 10), 388 => to_unsigned(565, 10), 389 => to_unsigned(866, 10), 390 => to_unsigned(942, 10), 391 => to_unsigned(673, 10), 392 => to_unsigned(1018, 10), 393 => to_unsigned(653, 10), 394 => to_unsigned(481, 10), 395 => to_unsigned(455, 10), 396 => to_unsigned(524, 10), 397 => to_unsigned(201, 10), 398 => to_unsigned(430, 10), 399 => to_unsigned(285, 10), 400 => to_unsigned(268, 10), 401 => to_unsigned(695, 10), 402 => to_unsigned(48, 10), 403 => to_unsigned(246, 10), 404 => to_unsigned(803, 10), 405 => to_unsigned(34, 10), 406 => to_unsigned(58, 10), 407 => to_unsigned(700, 10), 408 => to_unsigned(641, 10), 409 => to_unsigned(657, 10), 410 => to_unsigned(171, 10), 411 => to_unsigned(752, 10), 412 => to_unsigned(439, 10), 413 => to_unsigned(9, 10), 414 => to_unsigned(439, 10), 415 => to_unsigned(761, 10), 416 => to_unsigned(1021, 10), 417 => to_unsigned(656, 10), 418 => to_unsigned(835, 10), 419 => to_unsigned(681, 10), 420 => to_unsigned(470, 10), 421 => to_unsigned(815, 10), 422 => to_unsigned(724, 10), 423 => to_unsigned(88, 10), 424 => to_unsigned(225, 10), 425 => to_unsigned(507, 10), 426 => to_unsigned(826, 10), 427 => to_unsigned(980, 10), 428 => to_unsigned(213, 10), 429 => to_unsigned(804, 10), 430 => to_unsigned(748, 10), 431 => to_unsigned(268, 10), 432 => to_unsigned(26, 10), 433 => to_unsigned(2, 10), 434 => to_unsigned(1018, 10), 435 => to_unsigned(762, 10), 436 => to_unsigned(790, 10), 437 => to_unsigned(558, 10), 438 => to_unsigned(851, 10), 439 => to_unsigned(249, 10), 440 => to_unsigned(18, 10), 441 => to_unsigned(34, 10), 442 => to_unsigned(95, 10), 443 => to_unsigned(195, 10), 444 => to_unsigned(0, 10), 445 => to_unsigned(667, 10), 446 => to_unsigned(48, 10), 447 => to_unsigned(494, 10), 448 => to_unsigned(726, 10), 449 => to_unsigned(500, 10), 450 => to_unsigned(899, 10), 451 => to_unsigned(764, 10), 452 => to_unsigned(992, 10), 453 => to_unsigned(11, 10), 454 => to_unsigned(624, 10), 455 => to_unsigned(728, 10), 456 => to_unsigned(156, 10), 457 => to_unsigned(296, 10), 458 => to_unsigned(201, 10), 459 => to_unsigned(770, 10), 460 => to_unsigned(462, 10), 461 => to_unsigned(571, 10), 462 => to_unsigned(1012, 10), 463 => to_unsigned(778, 10), 464 => to_unsigned(388, 10), 465 => to_unsigned(713, 10), 466 => to_unsigned(365, 10), 467 => to_unsigned(127, 10), 468 => to_unsigned(90, 10), 469 => to_unsigned(619, 10), 470 => to_unsigned(253, 10), 471 => to_unsigned(264, 10), 472 => to_unsigned(293, 10), 473 => to_unsigned(1000, 10), 474 => to_unsigned(226, 10), 475 => to_unsigned(1004, 10), 476 => to_unsigned(758, 10), 477 => to_unsigned(102, 10), 478 => to_unsigned(859, 10), 479 => to_unsigned(752, 10), 480 => to_unsigned(442, 10), 481 => to_unsigned(954, 10), 482 => to_unsigned(945, 10), 483 => to_unsigned(245, 10), 484 => to_unsigned(275, 10), 485 => to_unsigned(803, 10), 486 => to_unsigned(420, 10), 487 => to_unsigned(636, 10), 488 => to_unsigned(330, 10), 489 => to_unsigned(305, 10), 490 => to_unsigned(658, 10), 491 => to_unsigned(260, 10), 492 => to_unsigned(472, 10), 493 => to_unsigned(975, 10), 494 => to_unsigned(817, 10), 495 => to_unsigned(990, 10), 496 => to_unsigned(269, 10), 497 => to_unsigned(435, 10), 498 => to_unsigned(400, 10), 499 => to_unsigned(439, 10), 500 => to_unsigned(104, 10), 501 => to_unsigned(1005, 10), 502 => to_unsigned(715, 10), 503 => to_unsigned(61, 10), 504 => to_unsigned(354, 10), 505 => to_unsigned(273, 10), 506 => to_unsigned(710, 10), 507 => to_unsigned(536, 10), 508 => to_unsigned(605, 10), 509 => to_unsigned(221, 10), 510 => to_unsigned(578, 10), 511 => to_unsigned(203, 10), 512 => to_unsigned(1018, 10), 513 => to_unsigned(46, 10), 514 => to_unsigned(168, 10), 515 => to_unsigned(721, 10), 516 => to_unsigned(167, 10), 517 => to_unsigned(511, 10), 518 => to_unsigned(777, 10), 519 => to_unsigned(363, 10), 520 => to_unsigned(282, 10), 521 => to_unsigned(788, 10), 522 => to_unsigned(953, 10), 523 => to_unsigned(964, 10), 524 => to_unsigned(618, 10), 525 => to_unsigned(322, 10), 526 => to_unsigned(52, 10), 527 => to_unsigned(807, 10), 528 => to_unsigned(851, 10), 529 => to_unsigned(447, 10), 530 => to_unsigned(372, 10), 531 => to_unsigned(647, 10), 532 => to_unsigned(543, 10), 533 => to_unsigned(96, 10), 534 => to_unsigned(196, 10), 535 => to_unsigned(1012, 10), 536 => to_unsigned(155, 10), 537 => to_unsigned(152, 10), 538 => to_unsigned(1002, 10), 539 => to_unsigned(823, 10), 540 => to_unsigned(648, 10), 541 => to_unsigned(556, 10), 542 => to_unsigned(821, 10), 543 => to_unsigned(730, 10), 544 => to_unsigned(550, 10), 545 => to_unsigned(155, 10), 546 => to_unsigned(226, 10), 547 => to_unsigned(43, 10), 548 => to_unsigned(972, 10), 549 => to_unsigned(751, 10), 550 => to_unsigned(520, 10), 551 => to_unsigned(680, 10), 552 => to_unsigned(632, 10), 553 => to_unsigned(493, 10), 554 => to_unsigned(288, 10), 555 => to_unsigned(448, 10), 556 => to_unsigned(1007, 10), 557 => to_unsigned(721, 10), 558 => to_unsigned(716, 10), 559 => to_unsigned(528, 10), 560 => to_unsigned(117, 10), 561 => to_unsigned(760, 10), 562 => to_unsigned(331, 10), 563 => to_unsigned(591, 10), 564 => to_unsigned(220, 10), 565 => to_unsigned(563, 10), 566 => to_unsigned(448, 10), 567 => to_unsigned(878, 10), 568 => to_unsigned(732, 10), 569 => to_unsigned(932, 10), 570 => to_unsigned(60, 10), 571 => to_unsigned(530, 10), 572 => to_unsigned(721, 10), 573 => to_unsigned(153, 10), 574 => to_unsigned(552, 10), 575 => to_unsigned(921, 10), 576 => to_unsigned(772, 10), 577 => to_unsigned(906, 10), 578 => to_unsigned(97, 10), 579 => to_unsigned(86, 10), 580 => to_unsigned(225, 10), 581 => to_unsigned(366, 10), 582 => to_unsigned(210, 10), 583 => to_unsigned(675, 10), 584 => to_unsigned(752, 10), 585 => to_unsigned(596, 10), 586 => to_unsigned(901, 10), 587 => to_unsigned(314, 10), 588 => to_unsigned(611, 10), 589 => to_unsigned(431, 10), 590 => to_unsigned(461, 10), 591 => to_unsigned(488, 10), 592 => to_unsigned(103, 10), 593 => to_unsigned(414, 10), 594 => to_unsigned(395, 10), 595 => to_unsigned(8, 10), 596 => to_unsigned(121, 10), 597 => to_unsigned(26, 10), 598 => to_unsigned(104, 10), 599 => to_unsigned(95, 10), 600 => to_unsigned(986, 10), 601 => to_unsigned(562, 10), 602 => to_unsigned(229, 10), 603 => to_unsigned(19, 10), 604 => to_unsigned(439, 10), 605 => to_unsigned(252, 10), 606 => to_unsigned(799, 10), 607 => to_unsigned(966, 10), 608 => to_unsigned(947, 10), 609 => to_unsigned(293, 10), 610 => to_unsigned(651, 10), 611 => to_unsigned(335, 10), 612 => to_unsigned(940, 10), 613 => to_unsigned(309, 10), 614 => to_unsigned(132, 10), 615 => to_unsigned(483, 10), 616 => to_unsigned(242, 10), 617 => to_unsigned(913, 10), 618 => to_unsigned(492, 10), 619 => to_unsigned(537, 10), 620 => to_unsigned(950, 10), 621 => to_unsigned(378, 10), 622 => to_unsigned(588, 10), 623 => to_unsigned(768, 10), 624 => to_unsigned(864, 10), 625 => to_unsigned(966, 10), 626 => to_unsigned(739, 10), 627 => to_unsigned(425, 10), 628 => to_unsigned(360, 10), 629 => to_unsigned(83, 10), 630 => to_unsigned(635, 10), 631 => to_unsigned(99, 10), 632 => to_unsigned(349, 10), 633 => to_unsigned(490, 10), 634 => to_unsigned(727, 10), 635 => to_unsigned(793, 10), 636 => to_unsigned(212, 10), 637 => to_unsigned(891, 10), 638 => to_unsigned(428, 10), 639 => to_unsigned(328, 10), 640 => to_unsigned(38, 10), 641 => to_unsigned(470, 10), 642 => to_unsigned(231, 10), 643 => to_unsigned(306, 10), 644 => to_unsigned(1013, 10), 645 => to_unsigned(655, 10), 646 => to_unsigned(511, 10), 647 => to_unsigned(900, 10), 648 => to_unsigned(715, 10), 649 => to_unsigned(282, 10), 650 => to_unsigned(75, 10), 651 => to_unsigned(794, 10), 652 => to_unsigned(972, 10), 653 => to_unsigned(796, 10), 654 => to_unsigned(896, 10), 655 => to_unsigned(325, 10), 656 => to_unsigned(57, 10), 657 => to_unsigned(486, 10), 658 => to_unsigned(525, 10), 659 => to_unsigned(790, 10), 660 => to_unsigned(763, 10), 661 => to_unsigned(251, 10), 662 => to_unsigned(984, 10), 663 => to_unsigned(317, 10), 664 => to_unsigned(602, 10), 665 => to_unsigned(574, 10), 666 => to_unsigned(645, 10), 667 => to_unsigned(850, 10), 668 => to_unsigned(812, 10), 669 => to_unsigned(366, 10), 670 => to_unsigned(220, 10), 671 => to_unsigned(579, 10), 672 => to_unsigned(23, 10), 673 => to_unsigned(905, 10), 674 => to_unsigned(435, 10), 675 => to_unsigned(517, 10), 676 => to_unsigned(218, 10), 677 => to_unsigned(545, 10), 678 => to_unsigned(129, 10), 679 => to_unsigned(63, 10), 680 => to_unsigned(480, 10), 681 => to_unsigned(84, 10), 682 => to_unsigned(505, 10), 683 => to_unsigned(701, 10), 684 => to_unsigned(495, 10), 685 => to_unsigned(347, 10), 686 => to_unsigned(746, 10), 687 => to_unsigned(204, 10), 688 => to_unsigned(287, 10), 689 => to_unsigned(237, 10), 690 => to_unsigned(475, 10), 691 => to_unsigned(954, 10), 692 => to_unsigned(387, 10), 693 => to_unsigned(243, 10), 694 => to_unsigned(596, 10), 695 => to_unsigned(394, 10), 696 => to_unsigned(179, 10), 697 => to_unsigned(73, 10), 698 => to_unsigned(965, 10), 699 => to_unsigned(141, 10), 700 => to_unsigned(316, 10), 701 => to_unsigned(616, 10), 702 => to_unsigned(849, 10), 703 => to_unsigned(442, 10), 704 => to_unsigned(301, 10), 705 => to_unsigned(153, 10), 706 => to_unsigned(899, 10), 707 => to_unsigned(448, 10), 708 => to_unsigned(758, 10), 709 => to_unsigned(718, 10), 710 => to_unsigned(244, 10), 711 => to_unsigned(782, 10), 712 => to_unsigned(215, 10), 713 => to_unsigned(966, 10), 714 => to_unsigned(271, 10), 715 => to_unsigned(517, 10), 716 => to_unsigned(822, 10), 717 => to_unsigned(512, 10), 718 => to_unsigned(743, 10), 719 => to_unsigned(711, 10), 720 => to_unsigned(957, 10), 721 => to_unsigned(337, 10), 722 => to_unsigned(800, 10), 723 => to_unsigned(58, 10), 724 => to_unsigned(541, 10), 725 => to_unsigned(927, 10), 726 => to_unsigned(463, 10), 727 => to_unsigned(715, 10), 728 => to_unsigned(1003, 10), 729 => to_unsigned(415, 10), 730 => to_unsigned(274, 10), 731 => to_unsigned(107, 10), 732 => to_unsigned(102, 10), 733 => to_unsigned(470, 10), 734 => to_unsigned(327, 10), 735 => to_unsigned(756, 10), 736 => to_unsigned(483, 10), 737 => to_unsigned(702, 10), 738 => to_unsigned(531, 10), 739 => to_unsigned(325, 10), 740 => to_unsigned(689, 10), 741 => to_unsigned(192, 10), 742 => to_unsigned(491, 10), 743 => to_unsigned(385, 10), 744 => to_unsigned(818, 10), 745 => to_unsigned(693, 10), 746 => to_unsigned(572, 10), 747 => to_unsigned(570, 10), 748 => to_unsigned(974, 10), 749 => to_unsigned(884, 10), 750 => to_unsigned(697, 10), 751 => to_unsigned(658, 10), 752 => to_unsigned(169, 10), 753 => to_unsigned(774, 10), 754 => to_unsigned(228, 10), 755 => to_unsigned(171, 10), 756 => to_unsigned(753, 10), 757 => to_unsigned(928, 10), 758 => to_unsigned(843, 10), 759 => to_unsigned(215, 10), 760 => to_unsigned(635, 10), 761 => to_unsigned(792, 10), 762 => to_unsigned(50, 10), 763 => to_unsigned(392, 10), 764 => to_unsigned(117, 10), 765 => to_unsigned(595, 10), 766 => to_unsigned(258, 10), 767 => to_unsigned(498, 10), 768 => to_unsigned(28, 10), 769 => to_unsigned(38, 10), 770 => to_unsigned(248, 10), 771 => to_unsigned(430, 10), 772 => to_unsigned(811, 10), 773 => to_unsigned(865, 10), 774 => to_unsigned(884, 10), 775 => to_unsigned(13, 10), 776 => to_unsigned(301, 10), 777 => to_unsigned(545, 10), 778 => to_unsigned(778, 10), 779 => to_unsigned(883, 10), 780 => to_unsigned(855, 10), 781 => to_unsigned(893, 10), 782 => to_unsigned(845, 10), 783 => to_unsigned(371, 10), 784 => to_unsigned(494, 10), 785 => to_unsigned(798, 10), 786 => to_unsigned(64, 10), 787 => to_unsigned(363, 10), 788 => to_unsigned(199, 10), 789 => to_unsigned(323, 10), 790 => to_unsigned(638, 10), 791 => to_unsigned(366, 10), 792 => to_unsigned(128, 10), 793 => to_unsigned(863, 10), 794 => to_unsigned(392, 10), 795 => to_unsigned(323, 10), 796 => to_unsigned(523, 10), 797 => to_unsigned(407, 10), 798 => to_unsigned(532, 10), 799 => to_unsigned(769, 10), 800 => to_unsigned(710, 10), 801 => to_unsigned(238, 10), 802 => to_unsigned(1020, 10), 803 => to_unsigned(324, 10), 804 => to_unsigned(170, 10), 805 => to_unsigned(355, 10), 806 => to_unsigned(124, 10), 807 => to_unsigned(239, 10), 808 => to_unsigned(278, 10), 809 => to_unsigned(158, 10), 810 => to_unsigned(38, 10), 811 => to_unsigned(331, 10), 812 => to_unsigned(820, 10), 813 => to_unsigned(866, 10), 814 => to_unsigned(503, 10), 815 => to_unsigned(707, 10), 816 => to_unsigned(369, 10), 817 => to_unsigned(490, 10), 818 => to_unsigned(192, 10), 819 => to_unsigned(6, 10), 820 => to_unsigned(545, 10), 821 => to_unsigned(1022, 10), 822 => to_unsigned(285, 10), 823 => to_unsigned(341, 10), 824 => to_unsigned(14, 10), 825 => to_unsigned(820, 10), 826 => to_unsigned(598, 10), 827 => to_unsigned(91, 10), 828 => to_unsigned(195, 10), 829 => to_unsigned(881, 10), 830 => to_unsigned(1023, 10), 831 => to_unsigned(862, 10), 832 => to_unsigned(103, 10), 833 => to_unsigned(430, 10), 834 => to_unsigned(343, 10), 835 => to_unsigned(24, 10), 836 => to_unsigned(235, 10), 837 => to_unsigned(397, 10), 838 => to_unsigned(416, 10), 839 => to_unsigned(32, 10), 840 => to_unsigned(242, 10), 841 => to_unsigned(374, 10), 842 => to_unsigned(497, 10), 843 => to_unsigned(793, 10), 844 => to_unsigned(841, 10), 845 => to_unsigned(357, 10), 846 => to_unsigned(364, 10), 847 => to_unsigned(657, 10), 848 => to_unsigned(663, 10), 849 => to_unsigned(291, 10), 850 => to_unsigned(1019, 10), 851 => to_unsigned(377, 10), 852 => to_unsigned(803, 10), 853 => to_unsigned(674, 10), 854 => to_unsigned(84, 10), 855 => to_unsigned(453, 10), 856 => to_unsigned(788, 10), 857 => to_unsigned(774, 10), 858 => to_unsigned(904, 10), 859 => to_unsigned(768, 10), 860 => to_unsigned(829, 10), 861 => to_unsigned(748, 10), 862 => to_unsigned(601, 10), 863 => to_unsigned(358, 10), 864 => to_unsigned(71, 10), 865 => to_unsigned(457, 10), 866 => to_unsigned(378, 10), 867 => to_unsigned(774, 10), 868 => to_unsigned(221, 10), 869 => to_unsigned(453, 10), 870 => to_unsigned(932, 10), 871 => to_unsigned(669, 10), 872 => to_unsigned(103, 10), 873 => to_unsigned(531, 10), 874 => to_unsigned(559, 10), 875 => to_unsigned(406, 10), 876 => to_unsigned(67, 10), 877 => to_unsigned(135, 10), 878 => to_unsigned(568, 10), 879 => to_unsigned(93, 10), 880 => to_unsigned(212, 10), 881 => to_unsigned(840, 10), 882 => to_unsigned(658, 10), 883 => to_unsigned(406, 10), 884 => to_unsigned(150, 10), 885 => to_unsigned(469, 10), 886 => to_unsigned(558, 10), 887 => to_unsigned(295, 10), 888 => to_unsigned(568, 10), 889 => to_unsigned(162, 10), 890 => to_unsigned(572, 10), 891 => to_unsigned(610, 10), 892 => to_unsigned(1023, 10), 893 => to_unsigned(464, 10), 894 => to_unsigned(909, 10), 895 => to_unsigned(540, 10), 896 => to_unsigned(248, 10), 897 => to_unsigned(571, 10), 898 => to_unsigned(13, 10), 899 => to_unsigned(417, 10), 900 => to_unsigned(634, 10), 901 => to_unsigned(666, 10), 902 => to_unsigned(77, 10), 903 => to_unsigned(953, 10), 904 => to_unsigned(125, 10), 905 => to_unsigned(586, 10), 906 => to_unsigned(506, 10), 907 => to_unsigned(599, 10), 908 => to_unsigned(213, 10), 909 => to_unsigned(603, 10), 910 => to_unsigned(493, 10), 911 => to_unsigned(567, 10), 912 => to_unsigned(508, 10), 913 => to_unsigned(85, 10), 914 => to_unsigned(735, 10), 915 => to_unsigned(486, 10), 916 => to_unsigned(466, 10), 917 => to_unsigned(603, 10), 918 => to_unsigned(765, 10), 919 => to_unsigned(474, 10), 920 => to_unsigned(279, 10), 921 => to_unsigned(199, 10), 922 => to_unsigned(909, 10), 923 => to_unsigned(788, 10), 924 => to_unsigned(478, 10), 925 => to_unsigned(291, 10), 926 => to_unsigned(970, 10), 927 => to_unsigned(419, 10), 928 => to_unsigned(709, 10), 929 => to_unsigned(805, 10), 930 => to_unsigned(406, 10), 931 => to_unsigned(673, 10), 932 => to_unsigned(18, 10), 933 => to_unsigned(896, 10), 934 => to_unsigned(287, 10), 935 => to_unsigned(492, 10), 936 => to_unsigned(798, 10), 937 => to_unsigned(173, 10), 938 => to_unsigned(130, 10), 939 => to_unsigned(149, 10), 940 => to_unsigned(786, 10), 941 => to_unsigned(336, 10), 942 => to_unsigned(611, 10), 943 => to_unsigned(1023, 10), 944 => to_unsigned(780, 10), 945 => to_unsigned(840, 10), 946 => to_unsigned(380, 10), 947 => to_unsigned(986, 10), 948 => to_unsigned(700, 10), 949 => to_unsigned(99, 10), 950 => to_unsigned(905, 10), 951 => to_unsigned(31, 10), 952 => to_unsigned(236, 10), 953 => to_unsigned(49, 10), 954 => to_unsigned(319, 10), 955 => to_unsigned(107, 10), 956 => to_unsigned(815, 10), 957 => to_unsigned(896, 10), 958 => to_unsigned(941, 10), 959 => to_unsigned(892, 10), 960 => to_unsigned(822, 10), 961 => to_unsigned(980, 10), 962 => to_unsigned(732, 10), 963 => to_unsigned(806, 10), 964 => to_unsigned(36, 10), 965 => to_unsigned(414, 10), 966 => to_unsigned(33, 10), 967 => to_unsigned(99, 10), 968 => to_unsigned(105, 10), 969 => to_unsigned(630, 10), 970 => to_unsigned(382, 10), 971 => to_unsigned(538, 10), 972 => to_unsigned(814, 10), 973 => to_unsigned(18, 10), 974 => to_unsigned(728, 10), 975 => to_unsigned(344, 10), 976 => to_unsigned(462, 10), 977 => to_unsigned(220, 10), 978 => to_unsigned(498, 10), 979 => to_unsigned(553, 10), 980 => to_unsigned(275, 10), 981 => to_unsigned(770, 10), 982 => to_unsigned(298, 10), 983 => to_unsigned(561, 10), 984 => to_unsigned(250, 10), 985 => to_unsigned(669, 10), 986 => to_unsigned(449, 10), 987 => to_unsigned(789, 10), 988 => to_unsigned(886, 10), 989 => to_unsigned(721, 10), 990 => to_unsigned(503, 10), 991 => to_unsigned(857, 10), 992 => to_unsigned(78, 10), 993 => to_unsigned(889, 10), 994 => to_unsigned(86, 10), 995 => to_unsigned(207, 10), 996 => to_unsigned(754, 10), 997 => to_unsigned(466, 10), 998 => to_unsigned(1023, 10), 999 => to_unsigned(395, 10), 1000 => to_unsigned(310, 10), 1001 => to_unsigned(280, 10), 1002 => to_unsigned(837, 10), 1003 => to_unsigned(235, 10), 1004 => to_unsigned(518, 10), 1005 => to_unsigned(573, 10), 1006 => to_unsigned(41, 10), 1007 => to_unsigned(188, 10), 1008 => to_unsigned(107, 10), 1009 => to_unsigned(687, 10), 1010 => to_unsigned(396, 10), 1011 => to_unsigned(652, 10), 1012 => to_unsigned(301, 10), 1013 => to_unsigned(549, 10), 1014 => to_unsigned(338, 10), 1015 => to_unsigned(457, 10), 1016 => to_unsigned(200, 10), 1017 => to_unsigned(309, 10), 1018 => to_unsigned(552, 10), 1019 => to_unsigned(904, 10), 1020 => to_unsigned(256, 10), 1021 => to_unsigned(288, 10), 1022 => to_unsigned(396, 10), 1023 => to_unsigned(244, 10), 1024 => to_unsigned(20, 10), 1025 => to_unsigned(249, 10), 1026 => to_unsigned(1019, 10), 1027 => to_unsigned(501, 10), 1028 => to_unsigned(370, 10), 1029 => to_unsigned(783, 10), 1030 => to_unsigned(791, 10), 1031 => to_unsigned(446, 10), 1032 => to_unsigned(54, 10), 1033 => to_unsigned(364, 10), 1034 => to_unsigned(977, 10), 1035 => to_unsigned(343, 10), 1036 => to_unsigned(9, 10), 1037 => to_unsigned(621, 10), 1038 => to_unsigned(482, 10), 1039 => to_unsigned(480, 10), 1040 => to_unsigned(873, 10), 1041 => to_unsigned(582, 10), 1042 => to_unsigned(1015, 10), 1043 => to_unsigned(475, 10), 1044 => to_unsigned(675, 10), 1045 => to_unsigned(723, 10), 1046 => to_unsigned(934, 10), 1047 => to_unsigned(321, 10), 1048 => to_unsigned(289, 10), 1049 => to_unsigned(613, 10), 1050 => to_unsigned(353, 10), 1051 => to_unsigned(929, 10), 1052 => to_unsigned(131, 10), 1053 => to_unsigned(854, 10), 1054 => to_unsigned(357, 10), 1055 => to_unsigned(122, 10), 1056 => to_unsigned(690, 10), 1057 => to_unsigned(929, 10), 1058 => to_unsigned(515, 10), 1059 => to_unsigned(333, 10), 1060 => to_unsigned(418, 10), 1061 => to_unsigned(847, 10), 1062 => to_unsigned(939, 10), 1063 => to_unsigned(481, 10), 1064 => to_unsigned(30, 10), 1065 => to_unsigned(937, 10), 1066 => to_unsigned(924, 10), 1067 => to_unsigned(649, 10), 1068 => to_unsigned(779, 10), 1069 => to_unsigned(153, 10), 1070 => to_unsigned(752, 10), 1071 => to_unsigned(252, 10), 1072 => to_unsigned(313, 10), 1073 => to_unsigned(585, 10), 1074 => to_unsigned(508, 10), 1075 => to_unsigned(318, 10), 1076 => to_unsigned(96, 10), 1077 => to_unsigned(917, 10), 1078 => to_unsigned(996, 10), 1079 => to_unsigned(203, 10), 1080 => to_unsigned(675, 10), 1081 => to_unsigned(184, 10), 1082 => to_unsigned(889, 10), 1083 => to_unsigned(428, 10), 1084 => to_unsigned(706, 10), 1085 => to_unsigned(96, 10), 1086 => to_unsigned(92, 10), 1087 => to_unsigned(612, 10), 1088 => to_unsigned(760, 10), 1089 => to_unsigned(586, 10), 1090 => to_unsigned(355, 10), 1091 => to_unsigned(285, 10), 1092 => to_unsigned(189, 10), 1093 => to_unsigned(491, 10), 1094 => to_unsigned(41, 10), 1095 => to_unsigned(983, 10), 1096 => to_unsigned(933, 10), 1097 => to_unsigned(703, 10), 1098 => to_unsigned(157, 10), 1099 => to_unsigned(353, 10), 1100 => to_unsigned(253, 10), 1101 => to_unsigned(35, 10), 1102 => to_unsigned(746, 10), 1103 => to_unsigned(208, 10), 1104 => to_unsigned(84, 10), 1105 => to_unsigned(33, 10), 1106 => to_unsigned(643, 10), 1107 => to_unsigned(351, 10), 1108 => to_unsigned(237, 10), 1109 => to_unsigned(100, 10), 1110 => to_unsigned(968, 10), 1111 => to_unsigned(344, 10), 1112 => to_unsigned(702, 10), 1113 => to_unsigned(537, 10), 1114 => to_unsigned(857, 10), 1115 => to_unsigned(293, 10), 1116 => to_unsigned(714, 10), 1117 => to_unsigned(224, 10), 1118 => to_unsigned(707, 10), 1119 => to_unsigned(639, 10), 1120 => to_unsigned(703, 10), 1121 => to_unsigned(725, 10), 1122 => to_unsigned(1000, 10), 1123 => to_unsigned(589, 10), 1124 => to_unsigned(96, 10), 1125 => to_unsigned(618, 10), 1126 => to_unsigned(5, 10), 1127 => to_unsigned(277, 10), 1128 => to_unsigned(168, 10), 1129 => to_unsigned(141, 10), 1130 => to_unsigned(27, 10), 1131 => to_unsigned(546, 10), 1132 => to_unsigned(384, 10), 1133 => to_unsigned(567, 10), 1134 => to_unsigned(761, 10), 1135 => to_unsigned(44, 10), 1136 => to_unsigned(743, 10), 1137 => to_unsigned(176, 10), 1138 => to_unsigned(367, 10), 1139 => to_unsigned(307, 10), 1140 => to_unsigned(827, 10), 1141 => to_unsigned(529, 10), 1142 => to_unsigned(352, 10), 1143 => to_unsigned(504, 10), 1144 => to_unsigned(736, 10), 1145 => to_unsigned(779, 10), 1146 => to_unsigned(426, 10), 1147 => to_unsigned(710, 10), 1148 => to_unsigned(210, 10), 1149 => to_unsigned(801, 10), 1150 => to_unsigned(51, 10), 1151 => to_unsigned(436, 10), 1152 => to_unsigned(837, 10), 1153 => to_unsigned(81, 10), 1154 => to_unsigned(950, 10), 1155 => to_unsigned(266, 10), 1156 => to_unsigned(204, 10), 1157 => to_unsigned(41, 10), 1158 => to_unsigned(465, 10), 1159 => to_unsigned(927, 10), 1160 => to_unsigned(259, 10), 1161 => to_unsigned(744, 10), 1162 => to_unsigned(226, 10), 1163 => to_unsigned(426, 10), 1164 => to_unsigned(862, 10), 1165 => to_unsigned(646, 10), 1166 => to_unsigned(832, 10), 1167 => to_unsigned(4, 10), 1168 => to_unsigned(644, 10), 1169 => to_unsigned(575, 10), 1170 => to_unsigned(748, 10), 1171 => to_unsigned(448, 10), 1172 => to_unsigned(1011, 10), 1173 => to_unsigned(483, 10), 1174 => to_unsigned(342, 10), 1175 => to_unsigned(990, 10), 1176 => to_unsigned(487, 10), 1177 => to_unsigned(925, 10), 1178 => to_unsigned(790, 10), 1179 => to_unsigned(87, 10), 1180 => to_unsigned(305, 10), 1181 => to_unsigned(794, 10), 1182 => to_unsigned(118, 10), 1183 => to_unsigned(824, 10), 1184 => to_unsigned(139, 10), 1185 => to_unsigned(898, 10), 1186 => to_unsigned(981, 10), 1187 => to_unsigned(12, 10), 1188 => to_unsigned(976, 10), 1189 => to_unsigned(2, 10), 1190 => to_unsigned(91, 10), 1191 => to_unsigned(716, 10), 1192 => to_unsigned(117, 10), 1193 => to_unsigned(121, 10), 1194 => to_unsigned(633, 10), 1195 => to_unsigned(745, 10), 1196 => to_unsigned(35, 10), 1197 => to_unsigned(640, 10), 1198 => to_unsigned(317, 10), 1199 => to_unsigned(77, 10), 1200 => to_unsigned(511, 10), 1201 => to_unsigned(613, 10), 1202 => to_unsigned(402, 10), 1203 => to_unsigned(931, 10), 1204 => to_unsigned(522, 10), 1205 => to_unsigned(275, 10), 1206 => to_unsigned(748, 10), 1207 => to_unsigned(667, 10), 1208 => to_unsigned(265, 10), 1209 => to_unsigned(624, 10), 1210 => to_unsigned(422, 10), 1211 => to_unsigned(890, 10), 1212 => to_unsigned(780, 10), 1213 => to_unsigned(751, 10), 1214 => to_unsigned(230, 10), 1215 => to_unsigned(497, 10), 1216 => to_unsigned(102, 10), 1217 => to_unsigned(69, 10), 1218 => to_unsigned(342, 10), 1219 => to_unsigned(62, 10), 1220 => to_unsigned(12, 10), 1221 => to_unsigned(578, 10), 1222 => to_unsigned(59, 10), 1223 => to_unsigned(896, 10), 1224 => to_unsigned(497, 10), 1225 => to_unsigned(24, 10), 1226 => to_unsigned(362, 10), 1227 => to_unsigned(733, 10), 1228 => to_unsigned(476, 10), 1229 => to_unsigned(992, 10), 1230 => to_unsigned(132, 10), 1231 => to_unsigned(968, 10), 1232 => to_unsigned(402, 10), 1233 => to_unsigned(813, 10), 1234 => to_unsigned(476, 10), 1235 => to_unsigned(199, 10), 1236 => to_unsigned(584, 10), 1237 => to_unsigned(912, 10), 1238 => to_unsigned(598, 10), 1239 => to_unsigned(874, 10), 1240 => to_unsigned(79, 10), 1241 => to_unsigned(895, 10), 1242 => to_unsigned(276, 10), 1243 => to_unsigned(560, 10), 1244 => to_unsigned(469, 10), 1245 => to_unsigned(599, 10), 1246 => to_unsigned(481, 10), 1247 => to_unsigned(322, 10), 1248 => to_unsigned(560, 10), 1249 => to_unsigned(730, 10), 1250 => to_unsigned(139, 10), 1251 => to_unsigned(152, 10), 1252 => to_unsigned(399, 10), 1253 => to_unsigned(879, 10), 1254 => to_unsigned(665, 10), 1255 => to_unsigned(895, 10), 1256 => to_unsigned(901, 10), 1257 => to_unsigned(534, 10), 1258 => to_unsigned(310, 10), 1259 => to_unsigned(819, 10), 1260 => to_unsigned(162, 10), 1261 => to_unsigned(157, 10), 1262 => to_unsigned(140, 10), 1263 => to_unsigned(300, 10), 1264 => to_unsigned(826, 10), 1265 => to_unsigned(892, 10), 1266 => to_unsigned(276, 10), 1267 => to_unsigned(319, 10), 1268 => to_unsigned(942, 10), 1269 => to_unsigned(353, 10), 1270 => to_unsigned(587, 10), 1271 => to_unsigned(814, 10), 1272 => to_unsigned(350, 10), 1273 => to_unsigned(110, 10), 1274 => to_unsigned(760, 10), 1275 => to_unsigned(267, 10), 1276 => to_unsigned(966, 10), 1277 => to_unsigned(863, 10), 1278 => to_unsigned(802, 10), 1279 => to_unsigned(297, 10), 1280 => to_unsigned(149, 10), 1281 => to_unsigned(714, 10), 1282 => to_unsigned(91, 10), 1283 => to_unsigned(81, 10), 1284 => to_unsigned(486, 10), 1285 => to_unsigned(825, 10), 1286 => to_unsigned(390, 10), 1287 => to_unsigned(907, 10), 1288 => to_unsigned(189, 10), 1289 => to_unsigned(368, 10), 1290 => to_unsigned(989, 10), 1291 => to_unsigned(461, 10), 1292 => to_unsigned(878, 10), 1293 => to_unsigned(659, 10), 1294 => to_unsigned(249, 10), 1295 => to_unsigned(7, 10), 1296 => to_unsigned(313, 10), 1297 => to_unsigned(656, 10), 1298 => to_unsigned(838, 10), 1299 => to_unsigned(168, 10), 1300 => to_unsigned(975, 10), 1301 => to_unsigned(190, 10), 1302 => to_unsigned(194, 10), 1303 => to_unsigned(522, 10), 1304 => to_unsigned(297, 10), 1305 => to_unsigned(938, 10), 1306 => to_unsigned(424, 10), 1307 => to_unsigned(925, 10), 1308 => to_unsigned(74, 10), 1309 => to_unsigned(330, 10), 1310 => to_unsigned(671, 10), 1311 => to_unsigned(593, 10), 1312 => to_unsigned(1019, 10), 1313 => to_unsigned(867, 10), 1314 => to_unsigned(932, 10), 1315 => to_unsigned(484, 10), 1316 => to_unsigned(61, 10), 1317 => to_unsigned(849, 10), 1318 => to_unsigned(881, 10), 1319 => to_unsigned(469, 10), 1320 => to_unsigned(923, 10), 1321 => to_unsigned(281, 10), 1322 => to_unsigned(943, 10), 1323 => to_unsigned(182, 10), 1324 => to_unsigned(456, 10), 1325 => to_unsigned(993, 10), 1326 => to_unsigned(762, 10), 1327 => to_unsigned(367, 10), 1328 => to_unsigned(457, 10), 1329 => to_unsigned(907, 10), 1330 => to_unsigned(176, 10), 1331 => to_unsigned(1007, 10), 1332 => to_unsigned(604, 10), 1333 => to_unsigned(784, 10), 1334 => to_unsigned(240, 10), 1335 => to_unsigned(962, 10), 1336 => to_unsigned(200, 10), 1337 => to_unsigned(417, 10), 1338 => to_unsigned(635, 10), 1339 => to_unsigned(688, 10), 1340 => to_unsigned(398, 10), 1341 => to_unsigned(680, 10), 1342 => to_unsigned(321, 10), 1343 => to_unsigned(686, 10), 1344 => to_unsigned(223, 10), 1345 => to_unsigned(790, 10), 1346 => to_unsigned(1005, 10), 1347 => to_unsigned(192, 10), 1348 => to_unsigned(716, 10), 1349 => to_unsigned(168, 10), 1350 => to_unsigned(760, 10), 1351 => to_unsigned(511, 10), 1352 => to_unsigned(448, 10), 1353 => to_unsigned(988, 10), 1354 => to_unsigned(159, 10), 1355 => to_unsigned(60, 10), 1356 => to_unsigned(382, 10), 1357 => to_unsigned(284, 10), 1358 => to_unsigned(124, 10), 1359 => to_unsigned(504, 10), 1360 => to_unsigned(697, 10), 1361 => to_unsigned(83, 10), 1362 => to_unsigned(1011, 10), 1363 => to_unsigned(96, 10), 1364 => to_unsigned(106, 10), 1365 => to_unsigned(299, 10), 1366 => to_unsigned(503, 10), 1367 => to_unsigned(580, 10), 1368 => to_unsigned(498, 10), 1369 => to_unsigned(721, 10), 1370 => to_unsigned(93, 10), 1371 => to_unsigned(486, 10), 1372 => to_unsigned(538, 10), 1373 => to_unsigned(729, 10), 1374 => to_unsigned(978, 10), 1375 => to_unsigned(435, 10), 1376 => to_unsigned(852, 10), 1377 => to_unsigned(303, 10), 1378 => to_unsigned(825, 10), 1379 => to_unsigned(41, 10), 1380 => to_unsigned(455, 10), 1381 => to_unsigned(226, 10), 1382 => to_unsigned(412, 10), 1383 => to_unsigned(672, 10), 1384 => to_unsigned(497, 10), 1385 => to_unsigned(486, 10), 1386 => to_unsigned(652, 10), 1387 => to_unsigned(600, 10), 1388 => to_unsigned(110, 10), 1389 => to_unsigned(494, 10), 1390 => to_unsigned(199, 10), 1391 => to_unsigned(457, 10), 1392 => to_unsigned(956, 10), 1393 => to_unsigned(295, 10), 1394 => to_unsigned(301, 10), 1395 => to_unsigned(161, 10), 1396 => to_unsigned(94, 10), 1397 => to_unsigned(995, 10), 1398 => to_unsigned(60, 10), 1399 => to_unsigned(930, 10), 1400 => to_unsigned(999, 10), 1401 => to_unsigned(450, 10), 1402 => to_unsigned(157, 10), 1403 => to_unsigned(888, 10), 1404 => to_unsigned(167, 10), 1405 => to_unsigned(831, 10), 1406 => to_unsigned(662, 10), 1407 => to_unsigned(739, 10), 1408 => to_unsigned(53, 10), 1409 => to_unsigned(704, 10), 1410 => to_unsigned(26, 10), 1411 => to_unsigned(68, 10), 1412 => to_unsigned(501, 10), 1413 => to_unsigned(43, 10), 1414 => to_unsigned(431, 10), 1415 => to_unsigned(137, 10), 1416 => to_unsigned(582, 10), 1417 => to_unsigned(925, 10), 1418 => to_unsigned(5, 10), 1419 => to_unsigned(513, 10), 1420 => to_unsigned(892, 10), 1421 => to_unsigned(598, 10), 1422 => to_unsigned(26, 10), 1423 => to_unsigned(861, 10), 1424 => to_unsigned(645, 10), 1425 => to_unsigned(400, 10), 1426 => to_unsigned(922, 10), 1427 => to_unsigned(300, 10), 1428 => to_unsigned(282, 10), 1429 => to_unsigned(78, 10), 1430 => to_unsigned(856, 10), 1431 => to_unsigned(648, 10), 1432 => to_unsigned(787, 10), 1433 => to_unsigned(989, 10), 1434 => to_unsigned(887, 10), 1435 => to_unsigned(315, 10), 1436 => to_unsigned(75, 10), 1437 => to_unsigned(174, 10), 1438 => to_unsigned(789, 10), 1439 => to_unsigned(450, 10), 1440 => to_unsigned(189, 10), 1441 => to_unsigned(57, 10), 1442 => to_unsigned(410, 10), 1443 => to_unsigned(53, 10), 1444 => to_unsigned(368, 10), 1445 => to_unsigned(1003, 10), 1446 => to_unsigned(452, 10), 1447 => to_unsigned(121, 10), 1448 => to_unsigned(918, 10), 1449 => to_unsigned(338, 10), 1450 => to_unsigned(678, 10), 1451 => to_unsigned(449, 10), 1452 => to_unsigned(644, 10), 1453 => to_unsigned(125, 10), 1454 => to_unsigned(231, 10), 1455 => to_unsigned(403, 10), 1456 => to_unsigned(859, 10), 1457 => to_unsigned(391, 10), 1458 => to_unsigned(368, 10), 1459 => to_unsigned(373, 10), 1460 => to_unsigned(477, 10), 1461 => to_unsigned(866, 10), 1462 => to_unsigned(856, 10), 1463 => to_unsigned(825, 10), 1464 => to_unsigned(460, 10), 1465 => to_unsigned(325, 10), 1466 => to_unsigned(556, 10), 1467 => to_unsigned(13, 10), 1468 => to_unsigned(496, 10), 1469 => to_unsigned(422, 10), 1470 => to_unsigned(207, 10), 1471 => to_unsigned(0, 10), 1472 => to_unsigned(113, 10), 1473 => to_unsigned(435, 10), 1474 => to_unsigned(708, 10), 1475 => to_unsigned(45, 10), 1476 => to_unsigned(662, 10), 1477 => to_unsigned(798, 10), 1478 => to_unsigned(509, 10), 1479 => to_unsigned(544, 10), 1480 => to_unsigned(631, 10), 1481 => to_unsigned(607, 10), 1482 => to_unsigned(45, 10), 1483 => to_unsigned(100, 10), 1484 => to_unsigned(899, 10), 1485 => to_unsigned(700, 10), 1486 => to_unsigned(931, 10), 1487 => to_unsigned(19, 10), 1488 => to_unsigned(610, 10), 1489 => to_unsigned(657, 10), 1490 => to_unsigned(236, 10), 1491 => to_unsigned(259, 10), 1492 => to_unsigned(700, 10), 1493 => to_unsigned(456, 10), 1494 => to_unsigned(65, 10), 1495 => to_unsigned(655, 10), 1496 => to_unsigned(873, 10), 1497 => to_unsigned(264, 10), 1498 => to_unsigned(376, 10), 1499 => to_unsigned(308, 10), 1500 => to_unsigned(918, 10), 1501 => to_unsigned(10, 10), 1502 => to_unsigned(44, 10), 1503 => to_unsigned(140, 10), 1504 => to_unsigned(3, 10), 1505 => to_unsigned(278, 10), 1506 => to_unsigned(652, 10), 1507 => to_unsigned(665, 10), 1508 => to_unsigned(693, 10), 1509 => to_unsigned(90, 10), 1510 => to_unsigned(552, 10), 1511 => to_unsigned(169, 10), 1512 => to_unsigned(640, 10), 1513 => to_unsigned(695, 10), 1514 => to_unsigned(59, 10), 1515 => to_unsigned(742, 10), 1516 => to_unsigned(180, 10), 1517 => to_unsigned(155, 10), 1518 => to_unsigned(552, 10), 1519 => to_unsigned(484, 10), 1520 => to_unsigned(725, 10), 1521 => to_unsigned(21, 10), 1522 => to_unsigned(454, 10), 1523 => to_unsigned(76, 10), 1524 => to_unsigned(647, 10), 1525 => to_unsigned(131, 10), 1526 => to_unsigned(504, 10), 1527 => to_unsigned(970, 10), 1528 => to_unsigned(27, 10), 1529 => to_unsigned(697, 10), 1530 => to_unsigned(241, 10), 1531 => to_unsigned(497, 10), 1532 => to_unsigned(344, 10), 1533 => to_unsigned(177, 10), 1534 => to_unsigned(174, 10), 1535 => to_unsigned(713, 10), 1536 => to_unsigned(492, 10), 1537 => to_unsigned(1004, 10), 1538 => to_unsigned(36, 10), 1539 => to_unsigned(520, 10), 1540 => to_unsigned(393, 10), 1541 => to_unsigned(483, 10), 1542 => to_unsigned(385, 10), 1543 => to_unsigned(678, 10), 1544 => to_unsigned(404, 10), 1545 => to_unsigned(45, 10), 1546 => to_unsigned(857, 10), 1547 => to_unsigned(172, 10), 1548 => to_unsigned(601, 10), 1549 => to_unsigned(965, 10), 1550 => to_unsigned(320, 10), 1551 => to_unsigned(1022, 10), 1552 => to_unsigned(103, 10), 1553 => to_unsigned(314, 10), 1554 => to_unsigned(966, 10), 1555 => to_unsigned(326, 10), 1556 => to_unsigned(615, 10), 1557 => to_unsigned(754, 10), 1558 => to_unsigned(529, 10), 1559 => to_unsigned(779, 10), 1560 => to_unsigned(17, 10), 1561 => to_unsigned(805, 10), 1562 => to_unsigned(606, 10), 1563 => to_unsigned(185, 10), 1564 => to_unsigned(1010, 10), 1565 => to_unsigned(881, 10), 1566 => to_unsigned(713, 10), 1567 => to_unsigned(780, 10), 1568 => to_unsigned(913, 10), 1569 => to_unsigned(638, 10), 1570 => to_unsigned(804, 10), 1571 => to_unsigned(672, 10), 1572 => to_unsigned(383, 10), 1573 => to_unsigned(899, 10), 1574 => to_unsigned(505, 10), 1575 => to_unsigned(886, 10), 1576 => to_unsigned(972, 10), 1577 => to_unsigned(117, 10), 1578 => to_unsigned(239, 10), 1579 => to_unsigned(677, 10), 1580 => to_unsigned(500, 10), 1581 => to_unsigned(711, 10), 1582 => to_unsigned(238, 10), 1583 => to_unsigned(701, 10), 1584 => to_unsigned(517, 10), 1585 => to_unsigned(145, 10), 1586 => to_unsigned(274, 10), 1587 => to_unsigned(530, 10), 1588 => to_unsigned(849, 10), 1589 => to_unsigned(545, 10), 1590 => to_unsigned(650, 10), 1591 => to_unsigned(305, 10), 1592 => to_unsigned(521, 10), 1593 => to_unsigned(666, 10), 1594 => to_unsigned(132, 10), 1595 => to_unsigned(872, 10), 1596 => to_unsigned(601, 10), 1597 => to_unsigned(114, 10), 1598 => to_unsigned(229, 10), 1599 => to_unsigned(327, 10), 1600 => to_unsigned(353, 10), 1601 => to_unsigned(785, 10), 1602 => to_unsigned(764, 10), 1603 => to_unsigned(495, 10), 1604 => to_unsigned(487, 10), 1605 => to_unsigned(624, 10), 1606 => to_unsigned(17, 10), 1607 => to_unsigned(870, 10), 1608 => to_unsigned(712, 10), 1609 => to_unsigned(614, 10), 1610 => to_unsigned(570, 10), 1611 => to_unsigned(87, 10), 1612 => to_unsigned(951, 10), 1613 => to_unsigned(162, 10), 1614 => to_unsigned(741, 10), 1615 => to_unsigned(987, 10), 1616 => to_unsigned(708, 10), 1617 => to_unsigned(642, 10), 1618 => to_unsigned(493, 10), 1619 => to_unsigned(881, 10), 1620 => to_unsigned(793, 10), 1621 => to_unsigned(326, 10), 1622 => to_unsigned(138, 10), 1623 => to_unsigned(531, 10), 1624 => to_unsigned(941, 10), 1625 => to_unsigned(847, 10), 1626 => to_unsigned(84, 10), 1627 => to_unsigned(437, 10), 1628 => to_unsigned(975, 10), 1629 => to_unsigned(182, 10), 1630 => to_unsigned(803, 10), 1631 => to_unsigned(943, 10), 1632 => to_unsigned(711, 10), 1633 => to_unsigned(872, 10), 1634 => to_unsigned(828, 10), 1635 => to_unsigned(548, 10), 1636 => to_unsigned(625, 10), 1637 => to_unsigned(924, 10), 1638 => to_unsigned(428, 10), 1639 => to_unsigned(558, 10), 1640 => to_unsigned(393, 10), 1641 => to_unsigned(356, 10), 1642 => to_unsigned(87, 10), 1643 => to_unsigned(163, 10), 1644 => to_unsigned(92, 10), 1645 => to_unsigned(18, 10), 1646 => to_unsigned(590, 10), 1647 => to_unsigned(743, 10), 1648 => to_unsigned(148, 10), 1649 => to_unsigned(36, 10), 1650 => to_unsigned(840, 10), 1651 => to_unsigned(368, 10), 1652 => to_unsigned(871, 10), 1653 => to_unsigned(525, 10), 1654 => to_unsigned(1015, 10), 1655 => to_unsigned(619, 10), 1656 => to_unsigned(488, 10), 1657 => to_unsigned(277, 10), 1658 => to_unsigned(315, 10), 1659 => to_unsigned(239, 10), 1660 => to_unsigned(189, 10), 1661 => to_unsigned(480, 10), 1662 => to_unsigned(288, 10), 1663 => to_unsigned(30, 10), 1664 => to_unsigned(585, 10), 1665 => to_unsigned(91, 10), 1666 => to_unsigned(445, 10), 1667 => to_unsigned(924, 10), 1668 => to_unsigned(824, 10), 1669 => to_unsigned(1003, 10), 1670 => to_unsigned(791, 10), 1671 => to_unsigned(348, 10), 1672 => to_unsigned(952, 10), 1673 => to_unsigned(322, 10), 1674 => to_unsigned(788, 10), 1675 => to_unsigned(342, 10), 1676 => to_unsigned(608, 10), 1677 => to_unsigned(903, 10), 1678 => to_unsigned(440, 10), 1679 => to_unsigned(277, 10), 1680 => to_unsigned(596, 10), 1681 => to_unsigned(915, 10), 1682 => to_unsigned(857, 10), 1683 => to_unsigned(175, 10), 1684 => to_unsigned(421, 10), 1685 => to_unsigned(88, 10), 1686 => to_unsigned(851, 10), 1687 => to_unsigned(439, 10), 1688 => to_unsigned(682, 10), 1689 => to_unsigned(525, 10), 1690 => to_unsigned(428, 10), 1691 => to_unsigned(603, 10), 1692 => to_unsigned(342, 10), 1693 => to_unsigned(347, 10), 1694 => to_unsigned(643, 10), 1695 => to_unsigned(441, 10), 1696 => to_unsigned(161, 10), 1697 => to_unsigned(797, 10), 1698 => to_unsigned(341, 10), 1699 => to_unsigned(66, 10), 1700 => to_unsigned(38, 10), 1701 => to_unsigned(408, 10), 1702 => to_unsigned(209, 10), 1703 => to_unsigned(589, 10), 1704 => to_unsigned(457, 10), 1705 => to_unsigned(745, 10), 1706 => to_unsigned(537, 10), 1707 => to_unsigned(37, 10), 1708 => to_unsigned(782, 10), 1709 => to_unsigned(925, 10), 1710 => to_unsigned(367, 10), 1711 => to_unsigned(903, 10), 1712 => to_unsigned(314, 10), 1713 => to_unsigned(923, 10), 1714 => to_unsigned(924, 10), 1715 => to_unsigned(854, 10), 1716 => to_unsigned(68, 10), 1717 => to_unsigned(963, 10), 1718 => to_unsigned(280, 10), 1719 => to_unsigned(231, 10), 1720 => to_unsigned(154, 10), 1721 => to_unsigned(250, 10), 1722 => to_unsigned(649, 10), 1723 => to_unsigned(955, 10), 1724 => to_unsigned(873, 10), 1725 => to_unsigned(244, 10), 1726 => to_unsigned(183, 10), 1727 => to_unsigned(839, 10), 1728 => to_unsigned(596, 10), 1729 => to_unsigned(395, 10), 1730 => to_unsigned(198, 10), 1731 => to_unsigned(348, 10), 1732 => to_unsigned(877, 10), 1733 => to_unsigned(258, 10), 1734 => to_unsigned(167, 10), 1735 => to_unsigned(569, 10), 1736 => to_unsigned(250, 10), 1737 => to_unsigned(923, 10), 1738 => to_unsigned(415, 10), 1739 => to_unsigned(931, 10), 1740 => to_unsigned(140, 10), 1741 => to_unsigned(832, 10), 1742 => to_unsigned(767, 10), 1743 => to_unsigned(663, 10), 1744 => to_unsigned(645, 10), 1745 => to_unsigned(695, 10), 1746 => to_unsigned(192, 10), 1747 => to_unsigned(803, 10), 1748 => to_unsigned(383, 10), 1749 => to_unsigned(10, 10), 1750 => to_unsigned(669, 10), 1751 => to_unsigned(319, 10), 1752 => to_unsigned(977, 10), 1753 => to_unsigned(816, 10), 1754 => to_unsigned(1000, 10), 1755 => to_unsigned(210, 10), 1756 => to_unsigned(571, 10), 1757 => to_unsigned(116, 10), 1758 => to_unsigned(175, 10), 1759 => to_unsigned(957, 10), 1760 => to_unsigned(138, 10), 1761 => to_unsigned(147, 10), 1762 => to_unsigned(741, 10), 1763 => to_unsigned(77, 10), 1764 => to_unsigned(185, 10), 1765 => to_unsigned(963, 10), 1766 => to_unsigned(548, 10), 1767 => to_unsigned(515, 10), 1768 => to_unsigned(419, 10), 1769 => to_unsigned(967, 10), 1770 => to_unsigned(758, 10), 1771 => to_unsigned(842, 10), 1772 => to_unsigned(84, 10), 1773 => to_unsigned(860, 10), 1774 => to_unsigned(584, 10), 1775 => to_unsigned(8, 10), 1776 => to_unsigned(465, 10), 1777 => to_unsigned(977, 10), 1778 => to_unsigned(380, 10), 1779 => to_unsigned(709, 10), 1780 => to_unsigned(991, 10), 1781 => to_unsigned(221, 10), 1782 => to_unsigned(955, 10), 1783 => to_unsigned(720, 10), 1784 => to_unsigned(441, 10), 1785 => to_unsigned(372, 10), 1786 => to_unsigned(854, 10), 1787 => to_unsigned(739, 10), 1788 => to_unsigned(562, 10), 1789 => to_unsigned(867, 10), 1790 => to_unsigned(592, 10), 1791 => to_unsigned(117, 10), 1792 => to_unsigned(411, 10), 1793 => to_unsigned(608, 10), 1794 => to_unsigned(303, 10), 1795 => to_unsigned(450, 10), 1796 => to_unsigned(11, 10), 1797 => to_unsigned(82, 10), 1798 => to_unsigned(216, 10), 1799 => to_unsigned(536, 10), 1800 => to_unsigned(128, 10), 1801 => to_unsigned(621, 10), 1802 => to_unsigned(444, 10), 1803 => to_unsigned(200, 10), 1804 => to_unsigned(87, 10), 1805 => to_unsigned(513, 10), 1806 => to_unsigned(251, 10), 1807 => to_unsigned(349, 10), 1808 => to_unsigned(47, 10), 1809 => to_unsigned(614, 10), 1810 => to_unsigned(230, 10), 1811 => to_unsigned(236, 10), 1812 => to_unsigned(1010, 10), 1813 => to_unsigned(434, 10), 1814 => to_unsigned(977, 10), 1815 => to_unsigned(211, 10), 1816 => to_unsigned(125, 10), 1817 => to_unsigned(729, 10), 1818 => to_unsigned(638, 10), 1819 => to_unsigned(965, 10), 1820 => to_unsigned(507, 10), 1821 => to_unsigned(750, 10), 1822 => to_unsigned(853, 10), 1823 => to_unsigned(546, 10), 1824 => to_unsigned(481, 10), 1825 => to_unsigned(806, 10), 1826 => to_unsigned(754, 10), 1827 => to_unsigned(895, 10), 1828 => to_unsigned(475, 10), 1829 => to_unsigned(361, 10), 1830 => to_unsigned(997, 10), 1831 => to_unsigned(817, 10), 1832 => to_unsigned(508, 10), 1833 => to_unsigned(900, 10), 1834 => to_unsigned(211, 10), 1835 => to_unsigned(819, 10), 1836 => to_unsigned(801, 10), 1837 => to_unsigned(853, 10), 1838 => to_unsigned(132, 10), 1839 => to_unsigned(435, 10), 1840 => to_unsigned(729, 10), 1841 => to_unsigned(893, 10), 1842 => to_unsigned(243, 10), 1843 => to_unsigned(71, 10), 1844 => to_unsigned(440, 10), 1845 => to_unsigned(638, 10), 1846 => to_unsigned(804, 10), 1847 => to_unsigned(563, 10), 1848 => to_unsigned(223, 10), 1849 => to_unsigned(61, 10), 1850 => to_unsigned(701, 10), 1851 => to_unsigned(367, 10), 1852 => to_unsigned(706, 10), 1853 => to_unsigned(953, 10), 1854 => to_unsigned(153, 10), 1855 => to_unsigned(908, 10), 1856 => to_unsigned(756, 10), 1857 => to_unsigned(957, 10), 1858 => to_unsigned(889, 10), 1859 => to_unsigned(381, 10), 1860 => to_unsigned(901, 10), 1861 => to_unsigned(675, 10), 1862 => to_unsigned(222, 10), 1863 => to_unsigned(244, 10), 1864 => to_unsigned(692, 10), 1865 => to_unsigned(649, 10), 1866 => to_unsigned(49, 10), 1867 => to_unsigned(1011, 10), 1868 => to_unsigned(465, 10), 1869 => to_unsigned(184, 10), 1870 => to_unsigned(157, 10), 1871 => to_unsigned(203, 10), 1872 => to_unsigned(189, 10), 1873 => to_unsigned(418, 10), 1874 => to_unsigned(1003, 10), 1875 => to_unsigned(248, 10), 1876 => to_unsigned(890, 10), 1877 => to_unsigned(939, 10), 1878 => to_unsigned(801, 10), 1879 => to_unsigned(890, 10), 1880 => to_unsigned(510, 10), 1881 => to_unsigned(156, 10), 1882 => to_unsigned(534, 10), 1883 => to_unsigned(89, 10), 1884 => to_unsigned(987, 10), 1885 => to_unsigned(17, 10), 1886 => to_unsigned(767, 10), 1887 => to_unsigned(33, 10), 1888 => to_unsigned(609, 10), 1889 => to_unsigned(1012, 10), 1890 => to_unsigned(601, 10), 1891 => to_unsigned(468, 10), 1892 => to_unsigned(379, 10), 1893 => to_unsigned(7, 10), 1894 => to_unsigned(192, 10), 1895 => to_unsigned(268, 10), 1896 => to_unsigned(241, 10), 1897 => to_unsigned(327, 10), 1898 => to_unsigned(940, 10), 1899 => to_unsigned(599, 10), 1900 => to_unsigned(550, 10), 1901 => to_unsigned(2, 10), 1902 => to_unsigned(955, 10), 1903 => to_unsigned(585, 10), 1904 => to_unsigned(926, 10), 1905 => to_unsigned(190, 10), 1906 => to_unsigned(306, 10), 1907 => to_unsigned(666, 10), 1908 => to_unsigned(524, 10), 1909 => to_unsigned(914, 10), 1910 => to_unsigned(487, 10), 1911 => to_unsigned(753, 10), 1912 => to_unsigned(413, 10), 1913 => to_unsigned(186, 10), 1914 => to_unsigned(1006, 10), 1915 => to_unsigned(934, 10), 1916 => to_unsigned(759, 10), 1917 => to_unsigned(326, 10), 1918 => to_unsigned(66, 10), 1919 => to_unsigned(636, 10), 1920 => to_unsigned(305, 10), 1921 => to_unsigned(461, 10), 1922 => to_unsigned(248, 10), 1923 => to_unsigned(691, 10), 1924 => to_unsigned(1023, 10), 1925 => to_unsigned(848, 10), 1926 => to_unsigned(799, 10), 1927 => to_unsigned(648, 10), 1928 => to_unsigned(873, 10), 1929 => to_unsigned(871, 10), 1930 => to_unsigned(671, 10), 1931 => to_unsigned(921, 10), 1932 => to_unsigned(18, 10), 1933 => to_unsigned(979, 10), 1934 => to_unsigned(860, 10), 1935 => to_unsigned(833, 10), 1936 => to_unsigned(441, 10), 1937 => to_unsigned(346, 10), 1938 => to_unsigned(115, 10), 1939 => to_unsigned(414, 10), 1940 => to_unsigned(405, 10), 1941 => to_unsigned(884, 10), 1942 => to_unsigned(843, 10), 1943 => to_unsigned(291, 10), 1944 => to_unsigned(994, 10), 1945 => to_unsigned(637, 10), 1946 => to_unsigned(182, 10), 1947 => to_unsigned(832, 10), 1948 => to_unsigned(761, 10), 1949 => to_unsigned(575, 10), 1950 => to_unsigned(728, 10), 1951 => to_unsigned(174, 10), 1952 => to_unsigned(608, 10), 1953 => to_unsigned(168, 10), 1954 => to_unsigned(570, 10), 1955 => to_unsigned(324, 10), 1956 => to_unsigned(413, 10), 1957 => to_unsigned(51, 10), 1958 => to_unsigned(54, 10), 1959 => to_unsigned(56, 10), 1960 => to_unsigned(1012, 10), 1961 => to_unsigned(850, 10), 1962 => to_unsigned(564, 10), 1963 => to_unsigned(101, 10), 1964 => to_unsigned(487, 10), 1965 => to_unsigned(66, 10), 1966 => to_unsigned(883, 10), 1967 => to_unsigned(545, 10), 1968 => to_unsigned(985, 10), 1969 => to_unsigned(923, 10), 1970 => to_unsigned(877, 10), 1971 => to_unsigned(470, 10), 1972 => to_unsigned(810, 10), 1973 => to_unsigned(881, 10), 1974 => to_unsigned(6, 10), 1975 => to_unsigned(949, 10), 1976 => to_unsigned(605, 10), 1977 => to_unsigned(32, 10), 1978 => to_unsigned(871, 10), 1979 => to_unsigned(407, 10), 1980 => to_unsigned(165, 10), 1981 => to_unsigned(650, 10), 1982 => to_unsigned(905, 10), 1983 => to_unsigned(321, 10), 1984 => to_unsigned(832, 10), 1985 => to_unsigned(515, 10), 1986 => to_unsigned(665, 10), 1987 => to_unsigned(189, 10), 1988 => to_unsigned(616, 10), 1989 => to_unsigned(716, 10), 1990 => to_unsigned(195, 10), 1991 => to_unsigned(738, 10), 1992 => to_unsigned(219, 10), 1993 => to_unsigned(49, 10), 1994 => to_unsigned(513, 10), 1995 => to_unsigned(776, 10), 1996 => to_unsigned(102, 10), 1997 => to_unsigned(97, 10), 1998 => to_unsigned(363, 10), 1999 => to_unsigned(95, 10), 2000 => to_unsigned(669, 10), 2001 => to_unsigned(560, 10), 2002 => to_unsigned(188, 10), 2003 => to_unsigned(764, 10), 2004 => to_unsigned(365, 10), 2005 => to_unsigned(205, 10), 2006 => to_unsigned(974, 10), 2007 => to_unsigned(668, 10), 2008 => to_unsigned(80, 10), 2009 => to_unsigned(739, 10), 2010 => to_unsigned(88, 10), 2011 => to_unsigned(301, 10), 2012 => to_unsigned(390, 10), 2013 => to_unsigned(274, 10), 2014 => to_unsigned(312, 10), 2015 => to_unsigned(673, 10), 2016 => to_unsigned(1020, 10), 2017 => to_unsigned(520, 10), 2018 => to_unsigned(846, 10), 2019 => to_unsigned(146, 10), 2020 => to_unsigned(489, 10), 2021 => to_unsigned(699, 10), 2022 => to_unsigned(551, 10), 2023 => to_unsigned(664, 10), 2024 => to_unsigned(908, 10), 2025 => to_unsigned(521, 10), 2026 => to_unsigned(496, 10), 2027 => to_unsigned(353, 10), 2028 => to_unsigned(255, 10), 2029 => to_unsigned(433, 10), 2030 => to_unsigned(353, 10), 2031 => to_unsigned(562, 10), 2032 => to_unsigned(728, 10), 2033 => to_unsigned(399, 10), 2034 => to_unsigned(238, 10), 2035 => to_unsigned(167, 10), 2036 => to_unsigned(326, 10), 2037 => to_unsigned(829, 10), 2038 => to_unsigned(401, 10), 2039 => to_unsigned(904, 10), 2040 => to_unsigned(111, 10), 2041 => to_unsigned(449, 10), 2042 => to_unsigned(647, 10), 2043 => to_unsigned(276, 10), 2044 => to_unsigned(680, 10), 2045 => to_unsigned(72, 10), 2046 => to_unsigned(372, 10), 2047 => to_unsigned(128, 10)),
            4 => (0 => to_unsigned(887, 10), 1 => to_unsigned(553, 10), 2 => to_unsigned(898, 10), 3 => to_unsigned(32, 10), 4 => to_unsigned(470, 10), 5 => to_unsigned(380, 10), 6 => to_unsigned(522, 10), 7 => to_unsigned(990, 10), 8 => to_unsigned(904, 10), 9 => to_unsigned(21, 10), 10 => to_unsigned(631, 10), 11 => to_unsigned(569, 10), 12 => to_unsigned(557, 10), 13 => to_unsigned(323, 10), 14 => to_unsigned(197, 10), 15 => to_unsigned(283, 10), 16 => to_unsigned(218, 10), 17 => to_unsigned(396, 10), 18 => to_unsigned(320, 10), 19 => to_unsigned(3, 10), 20 => to_unsigned(957, 10), 21 => to_unsigned(427, 10), 22 => to_unsigned(608, 10), 23 => to_unsigned(552, 10), 24 => to_unsigned(20, 10), 25 => to_unsigned(782, 10), 26 => to_unsigned(536, 10), 27 => to_unsigned(835, 10), 28 => to_unsigned(288, 10), 29 => to_unsigned(329, 10), 30 => to_unsigned(326, 10), 31 => to_unsigned(67, 10), 32 => to_unsigned(826, 10), 33 => to_unsigned(412, 10), 34 => to_unsigned(515, 10), 35 => to_unsigned(463, 10), 36 => to_unsigned(224, 10), 37 => to_unsigned(422, 10), 38 => to_unsigned(620, 10), 39 => to_unsigned(860, 10), 40 => to_unsigned(1013, 10), 41 => to_unsigned(754, 10), 42 => to_unsigned(709, 10), 43 => to_unsigned(1, 10), 44 => to_unsigned(145, 10), 45 => to_unsigned(190, 10), 46 => to_unsigned(431, 10), 47 => to_unsigned(264, 10), 48 => to_unsigned(329, 10), 49 => to_unsigned(436, 10), 50 => to_unsigned(909, 10), 51 => to_unsigned(880, 10), 52 => to_unsigned(553, 10), 53 => to_unsigned(24, 10), 54 => to_unsigned(575, 10), 55 => to_unsigned(964, 10), 56 => to_unsigned(71, 10), 57 => to_unsigned(69, 10), 58 => to_unsigned(615, 10), 59 => to_unsigned(660, 10), 60 => to_unsigned(835, 10), 61 => to_unsigned(449, 10), 62 => to_unsigned(201, 10), 63 => to_unsigned(346, 10), 64 => to_unsigned(833, 10), 65 => to_unsigned(168, 10), 66 => to_unsigned(368, 10), 67 => to_unsigned(358, 10), 68 => to_unsigned(942, 10), 69 => to_unsigned(405, 10), 70 => to_unsigned(332, 10), 71 => to_unsigned(70, 10), 72 => to_unsigned(416, 10), 73 => to_unsigned(426, 10), 74 => to_unsigned(852, 10), 75 => to_unsigned(716, 10), 76 => to_unsigned(342, 10), 77 => to_unsigned(20, 10), 78 => to_unsigned(109, 10), 79 => to_unsigned(929, 10), 80 => to_unsigned(928, 10), 81 => to_unsigned(777, 10), 82 => to_unsigned(187, 10), 83 => to_unsigned(612, 10), 84 => to_unsigned(1023, 10), 85 => to_unsigned(131, 10), 86 => to_unsigned(745, 10), 87 => to_unsigned(575, 10), 88 => to_unsigned(62, 10), 89 => to_unsigned(392, 10), 90 => to_unsigned(284, 10), 91 => to_unsigned(243, 10), 92 => to_unsigned(13, 10), 93 => to_unsigned(471, 10), 94 => to_unsigned(839, 10), 95 => to_unsigned(382, 10), 96 => to_unsigned(511, 10), 97 => to_unsigned(627, 10), 98 => to_unsigned(396, 10), 99 => to_unsigned(898, 10), 100 => to_unsigned(740, 10), 101 => to_unsigned(109, 10), 102 => to_unsigned(589, 10), 103 => to_unsigned(279, 10), 104 => to_unsigned(894, 10), 105 => to_unsigned(231, 10), 106 => to_unsigned(187, 10), 107 => to_unsigned(249, 10), 108 => to_unsigned(118, 10), 109 => to_unsigned(201, 10), 110 => to_unsigned(231, 10), 111 => to_unsigned(894, 10), 112 => to_unsigned(847, 10), 113 => to_unsigned(11, 10), 114 => to_unsigned(9, 10), 115 => to_unsigned(830, 10), 116 => to_unsigned(577, 10), 117 => to_unsigned(218, 10), 118 => to_unsigned(395, 10), 119 => to_unsigned(863, 10), 120 => to_unsigned(816, 10), 121 => to_unsigned(314, 10), 122 => to_unsigned(75, 10), 123 => to_unsigned(129, 10), 124 => to_unsigned(121, 10), 125 => to_unsigned(968, 10), 126 => to_unsigned(921, 10), 127 => to_unsigned(1016, 10), 128 => to_unsigned(286, 10), 129 => to_unsigned(417, 10), 130 => to_unsigned(236, 10), 131 => to_unsigned(87, 10), 132 => to_unsigned(788, 10), 133 => to_unsigned(817, 10), 134 => to_unsigned(904, 10), 135 => to_unsigned(320, 10), 136 => to_unsigned(930, 10), 137 => to_unsigned(670, 10), 138 => to_unsigned(870, 10), 139 => to_unsigned(468, 10), 140 => to_unsigned(165, 10), 141 => to_unsigned(790, 10), 142 => to_unsigned(573, 10), 143 => to_unsigned(298, 10), 144 => to_unsigned(304, 10), 145 => to_unsigned(982, 10), 146 => to_unsigned(105, 10), 147 => to_unsigned(20, 10), 148 => to_unsigned(939, 10), 149 => to_unsigned(391, 10), 150 => to_unsigned(705, 10), 151 => to_unsigned(120, 10), 152 => to_unsigned(429, 10), 153 => to_unsigned(542, 10), 154 => to_unsigned(652, 10), 155 => to_unsigned(453, 10), 156 => to_unsigned(824, 10), 157 => to_unsigned(149, 10), 158 => to_unsigned(197, 10), 159 => to_unsigned(16, 10), 160 => to_unsigned(555, 10), 161 => to_unsigned(382, 10), 162 => to_unsigned(535, 10), 163 => to_unsigned(168, 10), 164 => to_unsigned(1022, 10), 165 => to_unsigned(421, 10), 166 => to_unsigned(367, 10), 167 => to_unsigned(944, 10), 168 => to_unsigned(807, 10), 169 => to_unsigned(616, 10), 170 => to_unsigned(806, 10), 171 => to_unsigned(427, 10), 172 => to_unsigned(1018, 10), 173 => to_unsigned(688, 10), 174 => to_unsigned(896, 10), 175 => to_unsigned(137, 10), 176 => to_unsigned(764, 10), 177 => to_unsigned(911, 10), 178 => to_unsigned(436, 10), 179 => to_unsigned(748, 10), 180 => to_unsigned(53, 10), 181 => to_unsigned(766, 10), 182 => to_unsigned(388, 10), 183 => to_unsigned(668, 10), 184 => to_unsigned(497, 10), 185 => to_unsigned(35, 10), 186 => to_unsigned(532, 10), 187 => to_unsigned(262, 10), 188 => to_unsigned(553, 10), 189 => to_unsigned(927, 10), 190 => to_unsigned(217, 10), 191 => to_unsigned(848, 10), 192 => to_unsigned(964, 10), 193 => to_unsigned(238, 10), 194 => to_unsigned(397, 10), 195 => to_unsigned(929, 10), 196 => to_unsigned(145, 10), 197 => to_unsigned(111, 10), 198 => to_unsigned(577, 10), 199 => to_unsigned(601, 10), 200 => to_unsigned(559, 10), 201 => to_unsigned(342, 10), 202 => to_unsigned(554, 10), 203 => to_unsigned(150, 10), 204 => to_unsigned(977, 10), 205 => to_unsigned(835, 10), 206 => to_unsigned(147, 10), 207 => to_unsigned(814, 10), 208 => to_unsigned(285, 10), 209 => to_unsigned(758, 10), 210 => to_unsigned(324, 10), 211 => to_unsigned(468, 10), 212 => to_unsigned(365, 10), 213 => to_unsigned(926, 10), 214 => to_unsigned(684, 10), 215 => to_unsigned(463, 10), 216 => to_unsigned(929, 10), 217 => to_unsigned(1020, 10), 218 => to_unsigned(772, 10), 219 => to_unsigned(979, 10), 220 => to_unsigned(933, 10), 221 => to_unsigned(52, 10), 222 => to_unsigned(320, 10), 223 => to_unsigned(529, 10), 224 => to_unsigned(657, 10), 225 => to_unsigned(1009, 10), 226 => to_unsigned(423, 10), 227 => to_unsigned(616, 10), 228 => to_unsigned(274, 10), 229 => to_unsigned(389, 10), 230 => to_unsigned(866, 10), 231 => to_unsigned(899, 10), 232 => to_unsigned(314, 10), 233 => to_unsigned(512, 10), 234 => to_unsigned(631, 10), 235 => to_unsigned(547, 10), 236 => to_unsigned(281, 10), 237 => to_unsigned(340, 10), 238 => to_unsigned(605, 10), 239 => to_unsigned(449, 10), 240 => to_unsigned(910, 10), 241 => to_unsigned(556, 10), 242 => to_unsigned(742, 10), 243 => to_unsigned(260, 10), 244 => to_unsigned(710, 10), 245 => to_unsigned(657, 10), 246 => to_unsigned(221, 10), 247 => to_unsigned(445, 10), 248 => to_unsigned(824, 10), 249 => to_unsigned(897, 10), 250 => to_unsigned(272, 10), 251 => to_unsigned(194, 10), 252 => to_unsigned(590, 10), 253 => to_unsigned(362, 10), 254 => to_unsigned(689, 10), 255 => to_unsigned(24, 10), 256 => to_unsigned(837, 10), 257 => to_unsigned(889, 10), 258 => to_unsigned(405, 10), 259 => to_unsigned(520, 10), 260 => to_unsigned(712, 10), 261 => to_unsigned(289, 10), 262 => to_unsigned(69, 10), 263 => to_unsigned(608, 10), 264 => to_unsigned(1013, 10), 265 => to_unsigned(256, 10), 266 => to_unsigned(811, 10), 267 => to_unsigned(371, 10), 268 => to_unsigned(262, 10), 269 => to_unsigned(398, 10), 270 => to_unsigned(165, 10), 271 => to_unsigned(348, 10), 272 => to_unsigned(464, 10), 273 => to_unsigned(309, 10), 274 => to_unsigned(29, 10), 275 => to_unsigned(1012, 10), 276 => to_unsigned(978, 10), 277 => to_unsigned(861, 10), 278 => to_unsigned(632, 10), 279 => to_unsigned(122, 10), 280 => to_unsigned(741, 10), 281 => to_unsigned(131, 10), 282 => to_unsigned(1002, 10), 283 => to_unsigned(74, 10), 284 => to_unsigned(297, 10), 285 => to_unsigned(423, 10), 286 => to_unsigned(96, 10), 287 => to_unsigned(416, 10), 288 => to_unsigned(156, 10), 289 => to_unsigned(270, 10), 290 => to_unsigned(479, 10), 291 => to_unsigned(866, 10), 292 => to_unsigned(830, 10), 293 => to_unsigned(829, 10), 294 => to_unsigned(357, 10), 295 => to_unsigned(227, 10), 296 => to_unsigned(835, 10), 297 => to_unsigned(909, 10), 298 => to_unsigned(914, 10), 299 => to_unsigned(337, 10), 300 => to_unsigned(317, 10), 301 => to_unsigned(290, 10), 302 => to_unsigned(610, 10), 303 => to_unsigned(339, 10), 304 => to_unsigned(498, 10), 305 => to_unsigned(452, 10), 306 => to_unsigned(587, 10), 307 => to_unsigned(917, 10), 308 => to_unsigned(131, 10), 309 => to_unsigned(113, 10), 310 => to_unsigned(34, 10), 311 => to_unsigned(211, 10), 312 => to_unsigned(858, 10), 313 => to_unsigned(712, 10), 314 => to_unsigned(489, 10), 315 => to_unsigned(462, 10), 316 => to_unsigned(931, 10), 317 => to_unsigned(716, 10), 318 => to_unsigned(465, 10), 319 => to_unsigned(106, 10), 320 => to_unsigned(983, 10), 321 => to_unsigned(465, 10), 322 => to_unsigned(224, 10), 323 => to_unsigned(177, 10), 324 => to_unsigned(523, 10), 325 => to_unsigned(616, 10), 326 => to_unsigned(322, 10), 327 => to_unsigned(752, 10), 328 => to_unsigned(790, 10), 329 => to_unsigned(196, 10), 330 => to_unsigned(297, 10), 331 => to_unsigned(810, 10), 332 => to_unsigned(911, 10), 333 => to_unsigned(187, 10), 334 => to_unsigned(316, 10), 335 => to_unsigned(337, 10), 336 => to_unsigned(871, 10), 337 => to_unsigned(205, 10), 338 => to_unsigned(607, 10), 339 => to_unsigned(867, 10), 340 => to_unsigned(892, 10), 341 => to_unsigned(881, 10), 342 => to_unsigned(515, 10), 343 => to_unsigned(506, 10), 344 => to_unsigned(941, 10), 345 => to_unsigned(665, 10), 346 => to_unsigned(307, 10), 347 => to_unsigned(924, 10), 348 => to_unsigned(338, 10), 349 => to_unsigned(108, 10), 350 => to_unsigned(735, 10), 351 => to_unsigned(919, 10), 352 => to_unsigned(622, 10), 353 => to_unsigned(266, 10), 354 => to_unsigned(909, 10), 355 => to_unsigned(845, 10), 356 => to_unsigned(525, 10), 357 => to_unsigned(979, 10), 358 => to_unsigned(833, 10), 359 => to_unsigned(3, 10), 360 => to_unsigned(140, 10), 361 => to_unsigned(8, 10), 362 => to_unsigned(1011, 10), 363 => to_unsigned(778, 10), 364 => to_unsigned(893, 10), 365 => to_unsigned(774, 10), 366 => to_unsigned(820, 10), 367 => to_unsigned(415, 10), 368 => to_unsigned(887, 10), 369 => to_unsigned(299, 10), 370 => to_unsigned(991, 10), 371 => to_unsigned(661, 10), 372 => to_unsigned(269, 10), 373 => to_unsigned(327, 10), 374 => to_unsigned(301, 10), 375 => to_unsigned(540, 10), 376 => to_unsigned(338, 10), 377 => to_unsigned(925, 10), 378 => to_unsigned(317, 10), 379 => to_unsigned(410, 10), 380 => to_unsigned(306, 10), 381 => to_unsigned(527, 10), 382 => to_unsigned(942, 10), 383 => to_unsigned(833, 10), 384 => to_unsigned(109, 10), 385 => to_unsigned(691, 10), 386 => to_unsigned(793, 10), 387 => to_unsigned(530, 10), 388 => to_unsigned(1013, 10), 389 => to_unsigned(551, 10), 390 => to_unsigned(688, 10), 391 => to_unsigned(813, 10), 392 => to_unsigned(918, 10), 393 => to_unsigned(539, 10), 394 => to_unsigned(459, 10), 395 => to_unsigned(44, 10), 396 => to_unsigned(678, 10), 397 => to_unsigned(241, 10), 398 => to_unsigned(0, 10), 399 => to_unsigned(649, 10), 400 => to_unsigned(534, 10), 401 => to_unsigned(837, 10), 402 => to_unsigned(637, 10), 403 => to_unsigned(919, 10), 404 => to_unsigned(838, 10), 405 => to_unsigned(854, 10), 406 => to_unsigned(983, 10), 407 => to_unsigned(833, 10), 408 => to_unsigned(951, 10), 409 => to_unsigned(183, 10), 410 => to_unsigned(922, 10), 411 => to_unsigned(671, 10), 412 => to_unsigned(915, 10), 413 => to_unsigned(957, 10), 414 => to_unsigned(281, 10), 415 => to_unsigned(1000, 10), 416 => to_unsigned(839, 10), 417 => to_unsigned(523, 10), 418 => to_unsigned(379, 10), 419 => to_unsigned(185, 10), 420 => to_unsigned(567, 10), 421 => to_unsigned(785, 10), 422 => to_unsigned(950, 10), 423 => to_unsigned(104, 10), 424 => to_unsigned(256, 10), 425 => to_unsigned(779, 10), 426 => to_unsigned(548, 10), 427 => to_unsigned(739, 10), 428 => to_unsigned(205, 10), 429 => to_unsigned(764, 10), 430 => to_unsigned(264, 10), 431 => to_unsigned(319, 10), 432 => to_unsigned(998, 10), 433 => to_unsigned(394, 10), 434 => to_unsigned(729, 10), 435 => to_unsigned(745, 10), 436 => to_unsigned(9, 10), 437 => to_unsigned(630, 10), 438 => to_unsigned(84, 10), 439 => to_unsigned(260, 10), 440 => to_unsigned(443, 10), 441 => to_unsigned(39, 10), 442 => to_unsigned(720, 10), 443 => to_unsigned(466, 10), 444 => to_unsigned(750, 10), 445 => to_unsigned(718, 10), 446 => to_unsigned(215, 10), 447 => to_unsigned(750, 10), 448 => to_unsigned(308, 10), 449 => to_unsigned(355, 10), 450 => to_unsigned(123, 10), 451 => to_unsigned(560, 10), 452 => to_unsigned(286, 10), 453 => to_unsigned(3, 10), 454 => to_unsigned(10, 10), 455 => to_unsigned(288, 10), 456 => to_unsigned(149, 10), 457 => to_unsigned(937, 10), 458 => to_unsigned(890, 10), 459 => to_unsigned(110, 10), 460 => to_unsigned(353, 10), 461 => to_unsigned(658, 10), 462 => to_unsigned(225, 10), 463 => to_unsigned(179, 10), 464 => to_unsigned(204, 10), 465 => to_unsigned(191, 10), 466 => to_unsigned(564, 10), 467 => to_unsigned(450, 10), 468 => to_unsigned(857, 10), 469 => to_unsigned(490, 10), 470 => to_unsigned(478, 10), 471 => to_unsigned(691, 10), 472 => to_unsigned(348, 10), 473 => to_unsigned(169, 10), 474 => to_unsigned(785, 10), 475 => to_unsigned(910, 10), 476 => to_unsigned(827, 10), 477 => to_unsigned(828, 10), 478 => to_unsigned(13, 10), 479 => to_unsigned(609, 10), 480 => to_unsigned(790, 10), 481 => to_unsigned(244, 10), 482 => to_unsigned(957, 10), 483 => to_unsigned(344, 10), 484 => to_unsigned(414, 10), 485 => to_unsigned(906, 10), 486 => to_unsigned(643, 10), 487 => to_unsigned(159, 10), 488 => to_unsigned(1009, 10), 489 => to_unsigned(32, 10), 490 => to_unsigned(909, 10), 491 => to_unsigned(177, 10), 492 => to_unsigned(551, 10), 493 => to_unsigned(384, 10), 494 => to_unsigned(750, 10), 495 => to_unsigned(536, 10), 496 => to_unsigned(340, 10), 497 => to_unsigned(555, 10), 498 => to_unsigned(361, 10), 499 => to_unsigned(730, 10), 500 => to_unsigned(219, 10), 501 => to_unsigned(983, 10), 502 => to_unsigned(90, 10), 503 => to_unsigned(457, 10), 504 => to_unsigned(865, 10), 505 => to_unsigned(346, 10), 506 => to_unsigned(425, 10), 507 => to_unsigned(1007, 10), 508 => to_unsigned(159, 10), 509 => to_unsigned(552, 10), 510 => to_unsigned(223, 10), 511 => to_unsigned(264, 10), 512 => to_unsigned(433, 10), 513 => to_unsigned(676, 10), 514 => to_unsigned(337, 10), 515 => to_unsigned(862, 10), 516 => to_unsigned(385, 10), 517 => to_unsigned(186, 10), 518 => to_unsigned(285, 10), 519 => to_unsigned(245, 10), 520 => to_unsigned(208, 10), 521 => to_unsigned(84, 10), 522 => to_unsigned(648, 10), 523 => to_unsigned(631, 10), 524 => to_unsigned(292, 10), 525 => to_unsigned(861, 10), 526 => to_unsigned(699, 10), 527 => to_unsigned(235, 10), 528 => to_unsigned(108, 10), 529 => to_unsigned(271, 10), 530 => to_unsigned(13, 10), 531 => to_unsigned(665, 10), 532 => to_unsigned(766, 10), 533 => to_unsigned(229, 10), 534 => to_unsigned(720, 10), 535 => to_unsigned(818, 10), 536 => to_unsigned(907, 10), 537 => to_unsigned(302, 10), 538 => to_unsigned(130, 10), 539 => to_unsigned(161, 10), 540 => to_unsigned(476, 10), 541 => to_unsigned(602, 10), 542 => to_unsigned(681, 10), 543 => to_unsigned(257, 10), 544 => to_unsigned(410, 10), 545 => to_unsigned(456, 10), 546 => to_unsigned(339, 10), 547 => to_unsigned(411, 10), 548 => to_unsigned(761, 10), 549 => to_unsigned(611, 10), 550 => to_unsigned(150, 10), 551 => to_unsigned(729, 10), 552 => to_unsigned(216, 10), 553 => to_unsigned(364, 10), 554 => to_unsigned(852, 10), 555 => to_unsigned(932, 10), 556 => to_unsigned(245, 10), 557 => to_unsigned(920, 10), 558 => to_unsigned(542, 10), 559 => to_unsigned(652, 10), 560 => to_unsigned(820, 10), 561 => to_unsigned(247, 10), 562 => to_unsigned(746, 10), 563 => to_unsigned(568, 10), 564 => to_unsigned(220, 10), 565 => to_unsigned(754, 10), 566 => to_unsigned(68, 10), 567 => to_unsigned(961, 10), 568 => to_unsigned(69, 10), 569 => to_unsigned(172, 10), 570 => to_unsigned(341, 10), 571 => to_unsigned(762, 10), 572 => to_unsigned(625, 10), 573 => to_unsigned(920, 10), 574 => to_unsigned(136, 10), 575 => to_unsigned(760, 10), 576 => to_unsigned(492, 10), 577 => to_unsigned(122, 10), 578 => to_unsigned(368, 10), 579 => to_unsigned(378, 10), 580 => to_unsigned(414, 10), 581 => to_unsigned(288, 10), 582 => to_unsigned(341, 10), 583 => to_unsigned(963, 10), 584 => to_unsigned(185, 10), 585 => to_unsigned(885, 10), 586 => to_unsigned(852, 10), 587 => to_unsigned(337, 10), 588 => to_unsigned(126, 10), 589 => to_unsigned(145, 10), 590 => to_unsigned(331, 10), 591 => to_unsigned(402, 10), 592 => to_unsigned(889, 10), 593 => to_unsigned(675, 10), 594 => to_unsigned(826, 10), 595 => to_unsigned(597, 10), 596 => to_unsigned(493, 10), 597 => to_unsigned(299, 10), 598 => to_unsigned(447, 10), 599 => to_unsigned(354, 10), 600 => to_unsigned(371, 10), 601 => to_unsigned(97, 10), 602 => to_unsigned(969, 10), 603 => to_unsigned(155, 10), 604 => to_unsigned(983, 10), 605 => to_unsigned(959, 10), 606 => to_unsigned(1001, 10), 607 => to_unsigned(563, 10), 608 => to_unsigned(571, 10), 609 => to_unsigned(676, 10), 610 => to_unsigned(688, 10), 611 => to_unsigned(225, 10), 612 => to_unsigned(395, 10), 613 => to_unsigned(237, 10), 614 => to_unsigned(584, 10), 615 => to_unsigned(747, 10), 616 => to_unsigned(494, 10), 617 => to_unsigned(861, 10), 618 => to_unsigned(417, 10), 619 => to_unsigned(687, 10), 620 => to_unsigned(142, 10), 621 => to_unsigned(990, 10), 622 => to_unsigned(366, 10), 623 => to_unsigned(671, 10), 624 => to_unsigned(215, 10), 625 => to_unsigned(831, 10), 626 => to_unsigned(683, 10), 627 => to_unsigned(533, 10), 628 => to_unsigned(386, 10), 629 => to_unsigned(666, 10), 630 => to_unsigned(228, 10), 631 => to_unsigned(494, 10), 632 => to_unsigned(9, 10), 633 => to_unsigned(385, 10), 634 => to_unsigned(952, 10), 635 => to_unsigned(835, 10), 636 => to_unsigned(849, 10), 637 => to_unsigned(257, 10), 638 => to_unsigned(112, 10), 639 => to_unsigned(286, 10), 640 => to_unsigned(546, 10), 641 => to_unsigned(993, 10), 642 => to_unsigned(943, 10), 643 => to_unsigned(944, 10), 644 => to_unsigned(10, 10), 645 => to_unsigned(249, 10), 646 => to_unsigned(646, 10), 647 => to_unsigned(517, 10), 648 => to_unsigned(298, 10), 649 => to_unsigned(198, 10), 650 => to_unsigned(105, 10), 651 => to_unsigned(678, 10), 652 => to_unsigned(517, 10), 653 => to_unsigned(316, 10), 654 => to_unsigned(670, 10), 655 => to_unsigned(571, 10), 656 => to_unsigned(8, 10), 657 => to_unsigned(191, 10), 658 => to_unsigned(209, 10), 659 => to_unsigned(375, 10), 660 => to_unsigned(598, 10), 661 => to_unsigned(131, 10), 662 => to_unsigned(783, 10), 663 => to_unsigned(614, 10), 664 => to_unsigned(366, 10), 665 => to_unsigned(500, 10), 666 => to_unsigned(862, 10), 667 => to_unsigned(6, 10), 668 => to_unsigned(605, 10), 669 => to_unsigned(22, 10), 670 => to_unsigned(10, 10), 671 => to_unsigned(668, 10), 672 => to_unsigned(903, 10), 673 => to_unsigned(347, 10), 674 => to_unsigned(496, 10), 675 => to_unsigned(83, 10), 676 => to_unsigned(514, 10), 677 => to_unsigned(371, 10), 678 => to_unsigned(327, 10), 679 => to_unsigned(460, 10), 680 => to_unsigned(179, 10), 681 => to_unsigned(275, 10), 682 => to_unsigned(243, 10), 683 => to_unsigned(606, 10), 684 => to_unsigned(798, 10), 685 => to_unsigned(126, 10), 686 => to_unsigned(283, 10), 687 => to_unsigned(783, 10), 688 => to_unsigned(47, 10), 689 => to_unsigned(535, 10), 690 => to_unsigned(954, 10), 691 => to_unsigned(862, 10), 692 => to_unsigned(979, 10), 693 => to_unsigned(136, 10), 694 => to_unsigned(653, 10), 695 => to_unsigned(294, 10), 696 => to_unsigned(678, 10), 697 => to_unsigned(258, 10), 698 => to_unsigned(810, 10), 699 => to_unsigned(51, 10), 700 => to_unsigned(68, 10), 701 => to_unsigned(806, 10), 702 => to_unsigned(709, 10), 703 => to_unsigned(571, 10), 704 => to_unsigned(959, 10), 705 => to_unsigned(437, 10), 706 => to_unsigned(62, 10), 707 => to_unsigned(366, 10), 708 => to_unsigned(626, 10), 709 => to_unsigned(417, 10), 710 => to_unsigned(88, 10), 711 => to_unsigned(620, 10), 712 => to_unsigned(220, 10), 713 => to_unsigned(725, 10), 714 => to_unsigned(253, 10), 715 => to_unsigned(172, 10), 716 => to_unsigned(654, 10), 717 => to_unsigned(242, 10), 718 => to_unsigned(372, 10), 719 => to_unsigned(708, 10), 720 => to_unsigned(361, 10), 721 => to_unsigned(81, 10), 722 => to_unsigned(719, 10), 723 => to_unsigned(665, 10), 724 => to_unsigned(959, 10), 725 => to_unsigned(164, 10), 726 => to_unsigned(396, 10), 727 => to_unsigned(550, 10), 728 => to_unsigned(187, 10), 729 => to_unsigned(477, 10), 730 => to_unsigned(542, 10), 731 => to_unsigned(354, 10), 732 => to_unsigned(467, 10), 733 => to_unsigned(1002, 10), 734 => to_unsigned(851, 10), 735 => to_unsigned(543, 10), 736 => to_unsigned(1001, 10), 737 => to_unsigned(868, 10), 738 => to_unsigned(233, 10), 739 => to_unsigned(843, 10), 740 => to_unsigned(7, 10), 741 => to_unsigned(69, 10), 742 => to_unsigned(333, 10), 743 => to_unsigned(958, 10), 744 => to_unsigned(482, 10), 745 => to_unsigned(430, 10), 746 => to_unsigned(544, 10), 747 => to_unsigned(32, 10), 748 => to_unsigned(540, 10), 749 => to_unsigned(12, 10), 750 => to_unsigned(93, 10), 751 => to_unsigned(1011, 10), 752 => to_unsigned(74, 10), 753 => to_unsigned(1002, 10), 754 => to_unsigned(55, 10), 755 => to_unsigned(841, 10), 756 => to_unsigned(1011, 10), 757 => to_unsigned(305, 10), 758 => to_unsigned(507, 10), 759 => to_unsigned(19, 10), 760 => to_unsigned(214, 10), 761 => to_unsigned(407, 10), 762 => to_unsigned(542, 10), 763 => to_unsigned(956, 10), 764 => to_unsigned(436, 10), 765 => to_unsigned(781, 10), 766 => to_unsigned(498, 10), 767 => to_unsigned(799, 10), 768 => to_unsigned(186, 10), 769 => to_unsigned(252, 10), 770 => to_unsigned(656, 10), 771 => to_unsigned(786, 10), 772 => to_unsigned(897, 10), 773 => to_unsigned(15, 10), 774 => to_unsigned(672, 10), 775 => to_unsigned(78, 10), 776 => to_unsigned(841, 10), 777 => to_unsigned(774, 10), 778 => to_unsigned(755, 10), 779 => to_unsigned(879, 10), 780 => to_unsigned(195, 10), 781 => to_unsigned(70, 10), 782 => to_unsigned(886, 10), 783 => to_unsigned(207, 10), 784 => to_unsigned(733, 10), 785 => to_unsigned(853, 10), 786 => to_unsigned(179, 10), 787 => to_unsigned(842, 10), 788 => to_unsigned(186, 10), 789 => to_unsigned(973, 10), 790 => to_unsigned(859, 10), 791 => to_unsigned(922, 10), 792 => to_unsigned(538, 10), 793 => to_unsigned(745, 10), 794 => to_unsigned(580, 10), 795 => to_unsigned(827, 10), 796 => to_unsigned(925, 10), 797 => to_unsigned(688, 10), 798 => to_unsigned(348, 10), 799 => to_unsigned(317, 10), 800 => to_unsigned(700, 10), 801 => to_unsigned(911, 10), 802 => to_unsigned(878, 10), 803 => to_unsigned(505, 10), 804 => to_unsigned(91, 10), 805 => to_unsigned(424, 10), 806 => to_unsigned(160, 10), 807 => to_unsigned(685, 10), 808 => to_unsigned(113, 10), 809 => to_unsigned(398, 10), 810 => to_unsigned(836, 10), 811 => to_unsigned(345, 10), 812 => to_unsigned(480, 10), 813 => to_unsigned(268, 10), 814 => to_unsigned(684, 10), 815 => to_unsigned(873, 10), 816 => to_unsigned(315, 10), 817 => to_unsigned(426, 10), 818 => to_unsigned(959, 10), 819 => to_unsigned(820, 10), 820 => to_unsigned(397, 10), 821 => to_unsigned(436, 10), 822 => to_unsigned(178, 10), 823 => to_unsigned(120, 10), 824 => to_unsigned(946, 10), 825 => to_unsigned(881, 10), 826 => to_unsigned(965, 10), 827 => to_unsigned(471, 10), 828 => to_unsigned(741, 10), 829 => to_unsigned(628, 10), 830 => to_unsigned(990, 10), 831 => to_unsigned(476, 10), 832 => to_unsigned(182, 10), 833 => to_unsigned(981, 10), 834 => to_unsigned(851, 10), 835 => to_unsigned(856, 10), 836 => to_unsigned(377, 10), 837 => to_unsigned(687, 10), 838 => to_unsigned(599, 10), 839 => to_unsigned(941, 10), 840 => to_unsigned(62, 10), 841 => to_unsigned(266, 10), 842 => to_unsigned(606, 10), 843 => to_unsigned(96, 10), 844 => to_unsigned(981, 10), 845 => to_unsigned(872, 10), 846 => to_unsigned(54, 10), 847 => to_unsigned(862, 10), 848 => to_unsigned(646, 10), 849 => to_unsigned(921, 10), 850 => to_unsigned(517, 10), 851 => to_unsigned(695, 10), 852 => to_unsigned(735, 10), 853 => to_unsigned(47, 10), 854 => to_unsigned(494, 10), 855 => to_unsigned(411, 10), 856 => to_unsigned(345, 10), 857 => to_unsigned(417, 10), 858 => to_unsigned(731, 10), 859 => to_unsigned(912, 10), 860 => to_unsigned(656, 10), 861 => to_unsigned(335, 10), 862 => to_unsigned(734, 10), 863 => to_unsigned(418, 10), 864 => to_unsigned(443, 10), 865 => to_unsigned(69, 10), 866 => to_unsigned(72, 10), 867 => to_unsigned(656, 10), 868 => to_unsigned(230, 10), 869 => to_unsigned(819, 10), 870 => to_unsigned(487, 10), 871 => to_unsigned(604, 10), 872 => to_unsigned(645, 10), 873 => to_unsigned(0, 10), 874 => to_unsigned(723, 10), 875 => to_unsigned(535, 10), 876 => to_unsigned(508, 10), 877 => to_unsigned(158, 10), 878 => to_unsigned(756, 10), 879 => to_unsigned(622, 10), 880 => to_unsigned(806, 10), 881 => to_unsigned(680, 10), 882 => to_unsigned(738, 10), 883 => to_unsigned(593, 10), 884 => to_unsigned(639, 10), 885 => to_unsigned(911, 10), 886 => to_unsigned(74, 10), 887 => to_unsigned(274, 10), 888 => to_unsigned(488, 10), 889 => to_unsigned(283, 10), 890 => to_unsigned(307, 10), 891 => to_unsigned(892, 10), 892 => to_unsigned(426, 10), 893 => to_unsigned(486, 10), 894 => to_unsigned(718, 10), 895 => to_unsigned(815, 10), 896 => to_unsigned(337, 10), 897 => to_unsigned(252, 10), 898 => to_unsigned(375, 10), 899 => to_unsigned(169, 10), 900 => to_unsigned(236, 10), 901 => to_unsigned(899, 10), 902 => to_unsigned(496, 10), 903 => to_unsigned(117, 10), 904 => to_unsigned(921, 10), 905 => to_unsigned(216, 10), 906 => to_unsigned(876, 10), 907 => to_unsigned(991, 10), 908 => to_unsigned(215, 10), 909 => to_unsigned(1021, 10), 910 => to_unsigned(335, 10), 911 => to_unsigned(21, 10), 912 => to_unsigned(60, 10), 913 => to_unsigned(29, 10), 914 => to_unsigned(534, 10), 915 => to_unsigned(24, 10), 916 => to_unsigned(67, 10), 917 => to_unsigned(649, 10), 918 => to_unsigned(550, 10), 919 => to_unsigned(832, 10), 920 => to_unsigned(335, 10), 921 => to_unsigned(492, 10), 922 => to_unsigned(1001, 10), 923 => to_unsigned(142, 10), 924 => to_unsigned(581, 10), 925 => to_unsigned(81, 10), 926 => to_unsigned(698, 10), 927 => to_unsigned(361, 10), 928 => to_unsigned(579, 10), 929 => to_unsigned(240, 10), 930 => to_unsigned(211, 10), 931 => to_unsigned(82, 10), 932 => to_unsigned(363, 10), 933 => to_unsigned(689, 10), 934 => to_unsigned(625, 10), 935 => to_unsigned(385, 10), 936 => to_unsigned(647, 10), 937 => to_unsigned(520, 10), 938 => to_unsigned(543, 10), 939 => to_unsigned(636, 10), 940 => to_unsigned(270, 10), 941 => to_unsigned(206, 10), 942 => to_unsigned(404, 10), 943 => to_unsigned(146, 10), 944 => to_unsigned(751, 10), 945 => to_unsigned(163, 10), 946 => to_unsigned(812, 10), 947 => to_unsigned(1000, 10), 948 => to_unsigned(359, 10), 949 => to_unsigned(671, 10), 950 => to_unsigned(193, 10), 951 => to_unsigned(730, 10), 952 => to_unsigned(249, 10), 953 => to_unsigned(408, 10), 954 => to_unsigned(294, 10), 955 => to_unsigned(41, 10), 956 => to_unsigned(735, 10), 957 => to_unsigned(184, 10), 958 => to_unsigned(587, 10), 959 => to_unsigned(496, 10), 960 => to_unsigned(571, 10), 961 => to_unsigned(803, 10), 962 => to_unsigned(331, 10), 963 => to_unsigned(753, 10), 964 => to_unsigned(559, 10), 965 => to_unsigned(433, 10), 966 => to_unsigned(753, 10), 967 => to_unsigned(370, 10), 968 => to_unsigned(239, 10), 969 => to_unsigned(882, 10), 970 => to_unsigned(365, 10), 971 => to_unsigned(285, 10), 972 => to_unsigned(996, 10), 973 => to_unsigned(818, 10), 974 => to_unsigned(121, 10), 975 => to_unsigned(906, 10), 976 => to_unsigned(554, 10), 977 => to_unsigned(538, 10), 978 => to_unsigned(1020, 10), 979 => to_unsigned(203, 10), 980 => to_unsigned(697, 10), 981 => to_unsigned(105, 10), 982 => to_unsigned(455, 10), 983 => to_unsigned(893, 10), 984 => to_unsigned(372, 10), 985 => to_unsigned(736, 10), 986 => to_unsigned(219, 10), 987 => to_unsigned(263, 10), 988 => to_unsigned(439, 10), 989 => to_unsigned(212, 10), 990 => to_unsigned(401, 10), 991 => to_unsigned(74, 10), 992 => to_unsigned(988, 10), 993 => to_unsigned(710, 10), 994 => to_unsigned(568, 10), 995 => to_unsigned(412, 10), 996 => to_unsigned(255, 10), 997 => to_unsigned(656, 10), 998 => to_unsigned(61, 10), 999 => to_unsigned(836, 10), 1000 => to_unsigned(197, 10), 1001 => to_unsigned(472, 10), 1002 => to_unsigned(684, 10), 1003 => to_unsigned(310, 10), 1004 => to_unsigned(1008, 10), 1005 => to_unsigned(928, 10), 1006 => to_unsigned(622, 10), 1007 => to_unsigned(716, 10), 1008 => to_unsigned(439, 10), 1009 => to_unsigned(449, 10), 1010 => to_unsigned(751, 10), 1011 => to_unsigned(268, 10), 1012 => to_unsigned(409, 10), 1013 => to_unsigned(576, 10), 1014 => to_unsigned(325, 10), 1015 => to_unsigned(76, 10), 1016 => to_unsigned(926, 10), 1017 => to_unsigned(680, 10), 1018 => to_unsigned(913, 10), 1019 => to_unsigned(412, 10), 1020 => to_unsigned(500, 10), 1021 => to_unsigned(284, 10), 1022 => to_unsigned(11, 10), 1023 => to_unsigned(605, 10), 1024 => to_unsigned(577, 10), 1025 => to_unsigned(104, 10), 1026 => to_unsigned(384, 10), 1027 => to_unsigned(108, 10), 1028 => to_unsigned(690, 10), 1029 => to_unsigned(762, 10), 1030 => to_unsigned(411, 10), 1031 => to_unsigned(184, 10), 1032 => to_unsigned(1020, 10), 1033 => to_unsigned(79, 10), 1034 => to_unsigned(875, 10), 1035 => to_unsigned(692, 10), 1036 => to_unsigned(272, 10), 1037 => to_unsigned(346, 10), 1038 => to_unsigned(589, 10), 1039 => to_unsigned(537, 10), 1040 => to_unsigned(1001, 10), 1041 => to_unsigned(919, 10), 1042 => to_unsigned(316, 10), 1043 => to_unsigned(967, 10), 1044 => to_unsigned(403, 10), 1045 => to_unsigned(486, 10), 1046 => to_unsigned(577, 10), 1047 => to_unsigned(107, 10), 1048 => to_unsigned(446, 10), 1049 => to_unsigned(168, 10), 1050 => to_unsigned(324, 10), 1051 => to_unsigned(143, 10), 1052 => to_unsigned(21, 10), 1053 => to_unsigned(275, 10), 1054 => to_unsigned(668, 10), 1055 => to_unsigned(737, 10), 1056 => to_unsigned(650, 10), 1057 => to_unsigned(24, 10), 1058 => to_unsigned(153, 10), 1059 => to_unsigned(181, 10), 1060 => to_unsigned(519, 10), 1061 => to_unsigned(404, 10), 1062 => to_unsigned(867, 10), 1063 => to_unsigned(215, 10), 1064 => to_unsigned(702, 10), 1065 => to_unsigned(446, 10), 1066 => to_unsigned(974, 10), 1067 => to_unsigned(143, 10), 1068 => to_unsigned(644, 10), 1069 => to_unsigned(363, 10), 1070 => to_unsigned(612, 10), 1071 => to_unsigned(222, 10), 1072 => to_unsigned(96, 10), 1073 => to_unsigned(871, 10), 1074 => to_unsigned(490, 10), 1075 => to_unsigned(597, 10), 1076 => to_unsigned(627, 10), 1077 => to_unsigned(897, 10), 1078 => to_unsigned(690, 10), 1079 => to_unsigned(23, 10), 1080 => to_unsigned(64, 10), 1081 => to_unsigned(270, 10), 1082 => to_unsigned(475, 10), 1083 => to_unsigned(500, 10), 1084 => to_unsigned(205, 10), 1085 => to_unsigned(293, 10), 1086 => to_unsigned(564, 10), 1087 => to_unsigned(354, 10), 1088 => to_unsigned(716, 10), 1089 => to_unsigned(386, 10), 1090 => to_unsigned(114, 10), 1091 => to_unsigned(353, 10), 1092 => to_unsigned(503, 10), 1093 => to_unsigned(206, 10), 1094 => to_unsigned(913, 10), 1095 => to_unsigned(1001, 10), 1096 => to_unsigned(300, 10), 1097 => to_unsigned(711, 10), 1098 => to_unsigned(27, 10), 1099 => to_unsigned(407, 10), 1100 => to_unsigned(99, 10), 1101 => to_unsigned(751, 10), 1102 => to_unsigned(577, 10), 1103 => to_unsigned(71, 10), 1104 => to_unsigned(57, 10), 1105 => to_unsigned(503, 10), 1106 => to_unsigned(843, 10), 1107 => to_unsigned(185, 10), 1108 => to_unsigned(231, 10), 1109 => to_unsigned(266, 10), 1110 => to_unsigned(8, 10), 1111 => to_unsigned(782, 10), 1112 => to_unsigned(989, 10), 1113 => to_unsigned(607, 10), 1114 => to_unsigned(794, 10), 1115 => to_unsigned(819, 10), 1116 => to_unsigned(425, 10), 1117 => to_unsigned(976, 10), 1118 => to_unsigned(41, 10), 1119 => to_unsigned(759, 10), 1120 => to_unsigned(253, 10), 1121 => to_unsigned(813, 10), 1122 => to_unsigned(351, 10), 1123 => to_unsigned(666, 10), 1124 => to_unsigned(757, 10), 1125 => to_unsigned(101, 10), 1126 => to_unsigned(767, 10), 1127 => to_unsigned(965, 10), 1128 => to_unsigned(589, 10), 1129 => to_unsigned(777, 10), 1130 => to_unsigned(277, 10), 1131 => to_unsigned(2, 10), 1132 => to_unsigned(239, 10), 1133 => to_unsigned(416, 10), 1134 => to_unsigned(580, 10), 1135 => to_unsigned(124, 10), 1136 => to_unsigned(936, 10), 1137 => to_unsigned(774, 10), 1138 => to_unsigned(193, 10), 1139 => to_unsigned(309, 10), 1140 => to_unsigned(374, 10), 1141 => to_unsigned(359, 10), 1142 => to_unsigned(52, 10), 1143 => to_unsigned(574, 10), 1144 => to_unsigned(234, 10), 1145 => to_unsigned(831, 10), 1146 => to_unsigned(375, 10), 1147 => to_unsigned(204, 10), 1148 => to_unsigned(826, 10), 1149 => to_unsigned(429, 10), 1150 => to_unsigned(854, 10), 1151 => to_unsigned(1000, 10), 1152 => to_unsigned(588, 10), 1153 => to_unsigned(272, 10), 1154 => to_unsigned(323, 10), 1155 => to_unsigned(214, 10), 1156 => to_unsigned(767, 10), 1157 => to_unsigned(792, 10), 1158 => to_unsigned(133, 10), 1159 => to_unsigned(724, 10), 1160 => to_unsigned(765, 10), 1161 => to_unsigned(778, 10), 1162 => to_unsigned(104, 10), 1163 => to_unsigned(188, 10), 1164 => to_unsigned(345, 10), 1165 => to_unsigned(26, 10), 1166 => to_unsigned(665, 10), 1167 => to_unsigned(222, 10), 1168 => to_unsigned(281, 10), 1169 => to_unsigned(581, 10), 1170 => to_unsigned(283, 10), 1171 => to_unsigned(192, 10), 1172 => to_unsigned(801, 10), 1173 => to_unsigned(770, 10), 1174 => to_unsigned(457, 10), 1175 => to_unsigned(206, 10), 1176 => to_unsigned(445, 10), 1177 => to_unsigned(807, 10), 1178 => to_unsigned(407, 10), 1179 => to_unsigned(1003, 10), 1180 => to_unsigned(436, 10), 1181 => to_unsigned(197, 10), 1182 => to_unsigned(34, 10), 1183 => to_unsigned(479, 10), 1184 => to_unsigned(898, 10), 1185 => to_unsigned(356, 10), 1186 => to_unsigned(718, 10), 1187 => to_unsigned(795, 10), 1188 => to_unsigned(667, 10), 1189 => to_unsigned(192, 10), 1190 => to_unsigned(341, 10), 1191 => to_unsigned(1002, 10), 1192 => to_unsigned(248, 10), 1193 => to_unsigned(741, 10), 1194 => to_unsigned(785, 10), 1195 => to_unsigned(840, 10), 1196 => to_unsigned(136, 10), 1197 => to_unsigned(813, 10), 1198 => to_unsigned(781, 10), 1199 => to_unsigned(532, 10), 1200 => to_unsigned(624, 10), 1201 => to_unsigned(405, 10), 1202 => to_unsigned(343, 10), 1203 => to_unsigned(129, 10), 1204 => to_unsigned(934, 10), 1205 => to_unsigned(750, 10), 1206 => to_unsigned(824, 10), 1207 => to_unsigned(587, 10), 1208 => to_unsigned(664, 10), 1209 => to_unsigned(1015, 10), 1210 => to_unsigned(861, 10), 1211 => to_unsigned(415, 10), 1212 => to_unsigned(661, 10), 1213 => to_unsigned(732, 10), 1214 => to_unsigned(716, 10), 1215 => to_unsigned(732, 10), 1216 => to_unsigned(488, 10), 1217 => to_unsigned(321, 10), 1218 => to_unsigned(607, 10), 1219 => to_unsigned(950, 10), 1220 => to_unsigned(650, 10), 1221 => to_unsigned(732, 10), 1222 => to_unsigned(48, 10), 1223 => to_unsigned(874, 10), 1224 => to_unsigned(997, 10), 1225 => to_unsigned(789, 10), 1226 => to_unsigned(715, 10), 1227 => to_unsigned(499, 10), 1228 => to_unsigned(132, 10), 1229 => to_unsigned(1020, 10), 1230 => to_unsigned(486, 10), 1231 => to_unsigned(123, 10), 1232 => to_unsigned(108, 10), 1233 => to_unsigned(206, 10), 1234 => to_unsigned(437, 10), 1235 => to_unsigned(483, 10), 1236 => to_unsigned(504, 10), 1237 => to_unsigned(695, 10), 1238 => to_unsigned(999, 10), 1239 => to_unsigned(426, 10), 1240 => to_unsigned(760, 10), 1241 => to_unsigned(607, 10), 1242 => to_unsigned(555, 10), 1243 => to_unsigned(328, 10), 1244 => to_unsigned(763, 10), 1245 => to_unsigned(918, 10), 1246 => to_unsigned(551, 10), 1247 => to_unsigned(936, 10), 1248 => to_unsigned(34, 10), 1249 => to_unsigned(291, 10), 1250 => to_unsigned(500, 10), 1251 => to_unsigned(996, 10), 1252 => to_unsigned(436, 10), 1253 => to_unsigned(223, 10), 1254 => to_unsigned(766, 10), 1255 => to_unsigned(699, 10), 1256 => to_unsigned(420, 10), 1257 => to_unsigned(561, 10), 1258 => to_unsigned(530, 10), 1259 => to_unsigned(437, 10), 1260 => to_unsigned(397, 10), 1261 => to_unsigned(310, 10), 1262 => to_unsigned(246, 10), 1263 => to_unsigned(191, 10), 1264 => to_unsigned(697, 10), 1265 => to_unsigned(47, 10), 1266 => to_unsigned(907, 10), 1267 => to_unsigned(747, 10), 1268 => to_unsigned(242, 10), 1269 => to_unsigned(981, 10), 1270 => to_unsigned(704, 10), 1271 => to_unsigned(894, 10), 1272 => to_unsigned(634, 10), 1273 => to_unsigned(681, 10), 1274 => to_unsigned(657, 10), 1275 => to_unsigned(145, 10), 1276 => to_unsigned(765, 10), 1277 => to_unsigned(417, 10), 1278 => to_unsigned(40, 10), 1279 => to_unsigned(227, 10), 1280 => to_unsigned(419, 10), 1281 => to_unsigned(290, 10), 1282 => to_unsigned(859, 10), 1283 => to_unsigned(483, 10), 1284 => to_unsigned(115, 10), 1285 => to_unsigned(544, 10), 1286 => to_unsigned(664, 10), 1287 => to_unsigned(635, 10), 1288 => to_unsigned(9, 10), 1289 => to_unsigned(603, 10), 1290 => to_unsigned(941, 10), 1291 => to_unsigned(922, 10), 1292 => to_unsigned(525, 10), 1293 => to_unsigned(164, 10), 1294 => to_unsigned(298, 10), 1295 => to_unsigned(764, 10), 1296 => to_unsigned(280, 10), 1297 => to_unsigned(816, 10), 1298 => to_unsigned(307, 10), 1299 => to_unsigned(988, 10), 1300 => to_unsigned(496, 10), 1301 => to_unsigned(504, 10), 1302 => to_unsigned(483, 10), 1303 => to_unsigned(159, 10), 1304 => to_unsigned(672, 10), 1305 => to_unsigned(172, 10), 1306 => to_unsigned(602, 10), 1307 => to_unsigned(136, 10), 1308 => to_unsigned(17, 10), 1309 => to_unsigned(623, 10), 1310 => to_unsigned(662, 10), 1311 => to_unsigned(413, 10), 1312 => to_unsigned(768, 10), 1313 => to_unsigned(494, 10), 1314 => to_unsigned(518, 10), 1315 => to_unsigned(207, 10), 1316 => to_unsigned(149, 10), 1317 => to_unsigned(594, 10), 1318 => to_unsigned(963, 10), 1319 => to_unsigned(117, 10), 1320 => to_unsigned(115, 10), 1321 => to_unsigned(535, 10), 1322 => to_unsigned(314, 10), 1323 => to_unsigned(139, 10), 1324 => to_unsigned(54, 10), 1325 => to_unsigned(320, 10), 1326 => to_unsigned(228, 10), 1327 => to_unsigned(24, 10), 1328 => to_unsigned(964, 10), 1329 => to_unsigned(41, 10), 1330 => to_unsigned(290, 10), 1331 => to_unsigned(194, 10), 1332 => to_unsigned(136, 10), 1333 => to_unsigned(931, 10), 1334 => to_unsigned(1002, 10), 1335 => to_unsigned(644, 10), 1336 => to_unsigned(195, 10), 1337 => to_unsigned(420, 10), 1338 => to_unsigned(578, 10), 1339 => to_unsigned(908, 10), 1340 => to_unsigned(831, 10), 1341 => to_unsigned(345, 10), 1342 => to_unsigned(636, 10), 1343 => to_unsigned(792, 10), 1344 => to_unsigned(545, 10), 1345 => to_unsigned(943, 10), 1346 => to_unsigned(432, 10), 1347 => to_unsigned(300, 10), 1348 => to_unsigned(995, 10), 1349 => to_unsigned(824, 10), 1350 => to_unsigned(739, 10), 1351 => to_unsigned(393, 10), 1352 => to_unsigned(175, 10), 1353 => to_unsigned(900, 10), 1354 => to_unsigned(331, 10), 1355 => to_unsigned(360, 10), 1356 => to_unsigned(26, 10), 1357 => to_unsigned(777, 10), 1358 => to_unsigned(857, 10), 1359 => to_unsigned(123, 10), 1360 => to_unsigned(841, 10), 1361 => to_unsigned(412, 10), 1362 => to_unsigned(89, 10), 1363 => to_unsigned(749, 10), 1364 => to_unsigned(324, 10), 1365 => to_unsigned(542, 10), 1366 => to_unsigned(559, 10), 1367 => to_unsigned(417, 10), 1368 => to_unsigned(117, 10), 1369 => to_unsigned(605, 10), 1370 => to_unsigned(733, 10), 1371 => to_unsigned(468, 10), 1372 => to_unsigned(309, 10), 1373 => to_unsigned(760, 10), 1374 => to_unsigned(759, 10), 1375 => to_unsigned(336, 10), 1376 => to_unsigned(863, 10), 1377 => to_unsigned(422, 10), 1378 => to_unsigned(193, 10), 1379 => to_unsigned(321, 10), 1380 => to_unsigned(493, 10), 1381 => to_unsigned(670, 10), 1382 => to_unsigned(809, 10), 1383 => to_unsigned(1023, 10), 1384 => to_unsigned(1012, 10), 1385 => to_unsigned(165, 10), 1386 => to_unsigned(298, 10), 1387 => to_unsigned(513, 10), 1388 => to_unsigned(702, 10), 1389 => to_unsigned(5, 10), 1390 => to_unsigned(654, 10), 1391 => to_unsigned(137, 10), 1392 => to_unsigned(981, 10), 1393 => to_unsigned(579, 10), 1394 => to_unsigned(30, 10), 1395 => to_unsigned(663, 10), 1396 => to_unsigned(337, 10), 1397 => to_unsigned(138, 10), 1398 => to_unsigned(559, 10), 1399 => to_unsigned(1021, 10), 1400 => to_unsigned(439, 10), 1401 => to_unsigned(688, 10), 1402 => to_unsigned(390, 10), 1403 => to_unsigned(326, 10), 1404 => to_unsigned(21, 10), 1405 => to_unsigned(419, 10), 1406 => to_unsigned(235, 10), 1407 => to_unsigned(283, 10), 1408 => to_unsigned(912, 10), 1409 => to_unsigned(806, 10), 1410 => to_unsigned(164, 10), 1411 => to_unsigned(263, 10), 1412 => to_unsigned(14, 10), 1413 => to_unsigned(549, 10), 1414 => to_unsigned(964, 10), 1415 => to_unsigned(287, 10), 1416 => to_unsigned(584, 10), 1417 => to_unsigned(419, 10), 1418 => to_unsigned(327, 10), 1419 => to_unsigned(87, 10), 1420 => to_unsigned(314, 10), 1421 => to_unsigned(952, 10), 1422 => to_unsigned(579, 10), 1423 => to_unsigned(875, 10), 1424 => to_unsigned(465, 10), 1425 => to_unsigned(872, 10), 1426 => to_unsigned(892, 10), 1427 => to_unsigned(309, 10), 1428 => to_unsigned(923, 10), 1429 => to_unsigned(292, 10), 1430 => to_unsigned(996, 10), 1431 => to_unsigned(209, 10), 1432 => to_unsigned(673, 10), 1433 => to_unsigned(936, 10), 1434 => to_unsigned(365, 10), 1435 => to_unsigned(424, 10), 1436 => to_unsigned(723, 10), 1437 => to_unsigned(287, 10), 1438 => to_unsigned(882, 10), 1439 => to_unsigned(598, 10), 1440 => to_unsigned(515, 10), 1441 => to_unsigned(364, 10), 1442 => to_unsigned(512, 10), 1443 => to_unsigned(800, 10), 1444 => to_unsigned(901, 10), 1445 => to_unsigned(232, 10), 1446 => to_unsigned(775, 10), 1447 => to_unsigned(197, 10), 1448 => to_unsigned(143, 10), 1449 => to_unsigned(621, 10), 1450 => to_unsigned(984, 10), 1451 => to_unsigned(746, 10), 1452 => to_unsigned(587, 10), 1453 => to_unsigned(960, 10), 1454 => to_unsigned(250, 10), 1455 => to_unsigned(289, 10), 1456 => to_unsigned(418, 10), 1457 => to_unsigned(544, 10), 1458 => to_unsigned(318, 10), 1459 => to_unsigned(814, 10), 1460 => to_unsigned(184, 10), 1461 => to_unsigned(322, 10), 1462 => to_unsigned(312, 10), 1463 => to_unsigned(31, 10), 1464 => to_unsigned(592, 10), 1465 => to_unsigned(198, 10), 1466 => to_unsigned(522, 10), 1467 => to_unsigned(790, 10), 1468 => to_unsigned(182, 10), 1469 => to_unsigned(142, 10), 1470 => to_unsigned(163, 10), 1471 => to_unsigned(180, 10), 1472 => to_unsigned(579, 10), 1473 => to_unsigned(618, 10), 1474 => to_unsigned(816, 10), 1475 => to_unsigned(435, 10), 1476 => to_unsigned(230, 10), 1477 => to_unsigned(874, 10), 1478 => to_unsigned(570, 10), 1479 => to_unsigned(470, 10), 1480 => to_unsigned(173, 10), 1481 => to_unsigned(557, 10), 1482 => to_unsigned(758, 10), 1483 => to_unsigned(741, 10), 1484 => to_unsigned(889, 10), 1485 => to_unsigned(464, 10), 1486 => to_unsigned(865, 10), 1487 => to_unsigned(660, 10), 1488 => to_unsigned(510, 10), 1489 => to_unsigned(935, 10), 1490 => to_unsigned(610, 10), 1491 => to_unsigned(170, 10), 1492 => to_unsigned(445, 10), 1493 => to_unsigned(822, 10), 1494 => to_unsigned(864, 10), 1495 => to_unsigned(609, 10), 1496 => to_unsigned(497, 10), 1497 => to_unsigned(816, 10), 1498 => to_unsigned(689, 10), 1499 => to_unsigned(991, 10), 1500 => to_unsigned(341, 10), 1501 => to_unsigned(128, 10), 1502 => to_unsigned(534, 10), 1503 => to_unsigned(575, 10), 1504 => to_unsigned(849, 10), 1505 => to_unsigned(960, 10), 1506 => to_unsigned(293, 10), 1507 => to_unsigned(636, 10), 1508 => to_unsigned(557, 10), 1509 => to_unsigned(502, 10), 1510 => to_unsigned(47, 10), 1511 => to_unsigned(8, 10), 1512 => to_unsigned(1014, 10), 1513 => to_unsigned(432, 10), 1514 => to_unsigned(41, 10), 1515 => to_unsigned(929, 10), 1516 => to_unsigned(247, 10), 1517 => to_unsigned(85, 10), 1518 => to_unsigned(101, 10), 1519 => to_unsigned(608, 10), 1520 => to_unsigned(464, 10), 1521 => to_unsigned(17, 10), 1522 => to_unsigned(538, 10), 1523 => to_unsigned(773, 10), 1524 => to_unsigned(939, 10), 1525 => to_unsigned(918, 10), 1526 => to_unsigned(708, 10), 1527 => to_unsigned(312, 10), 1528 => to_unsigned(585, 10), 1529 => to_unsigned(213, 10), 1530 => to_unsigned(811, 10), 1531 => to_unsigned(917, 10), 1532 => to_unsigned(319, 10), 1533 => to_unsigned(952, 10), 1534 => to_unsigned(665, 10), 1535 => to_unsigned(911, 10), 1536 => to_unsigned(929, 10), 1537 => to_unsigned(114, 10), 1538 => to_unsigned(472, 10), 1539 => to_unsigned(197, 10), 1540 => to_unsigned(318, 10), 1541 => to_unsigned(710, 10), 1542 => to_unsigned(695, 10), 1543 => to_unsigned(141, 10), 1544 => to_unsigned(987, 10), 1545 => to_unsigned(268, 10), 1546 => to_unsigned(130, 10), 1547 => to_unsigned(596, 10), 1548 => to_unsigned(62, 10), 1549 => to_unsigned(758, 10), 1550 => to_unsigned(768, 10), 1551 => to_unsigned(19, 10), 1552 => to_unsigned(675, 10), 1553 => to_unsigned(854, 10), 1554 => to_unsigned(531, 10), 1555 => to_unsigned(761, 10), 1556 => to_unsigned(635, 10), 1557 => to_unsigned(385, 10), 1558 => to_unsigned(542, 10), 1559 => to_unsigned(503, 10), 1560 => to_unsigned(749, 10), 1561 => to_unsigned(995, 10), 1562 => to_unsigned(956, 10), 1563 => to_unsigned(204, 10), 1564 => to_unsigned(883, 10), 1565 => to_unsigned(243, 10), 1566 => to_unsigned(703, 10), 1567 => to_unsigned(25, 10), 1568 => to_unsigned(817, 10), 1569 => to_unsigned(529, 10), 1570 => to_unsigned(336, 10), 1571 => to_unsigned(271, 10), 1572 => to_unsigned(1014, 10), 1573 => to_unsigned(793, 10), 1574 => to_unsigned(79, 10), 1575 => to_unsigned(825, 10), 1576 => to_unsigned(1023, 10), 1577 => to_unsigned(936, 10), 1578 => to_unsigned(283, 10), 1579 => to_unsigned(266, 10), 1580 => to_unsigned(264, 10), 1581 => to_unsigned(753, 10), 1582 => to_unsigned(728, 10), 1583 => to_unsigned(510, 10), 1584 => to_unsigned(660, 10), 1585 => to_unsigned(236, 10), 1586 => to_unsigned(719, 10), 1587 => to_unsigned(222, 10), 1588 => to_unsigned(179, 10), 1589 => to_unsigned(857, 10), 1590 => to_unsigned(484, 10), 1591 => to_unsigned(568, 10), 1592 => to_unsigned(766, 10), 1593 => to_unsigned(649, 10), 1594 => to_unsigned(878, 10), 1595 => to_unsigned(863, 10), 1596 => to_unsigned(163, 10), 1597 => to_unsigned(457, 10), 1598 => to_unsigned(393, 10), 1599 => to_unsigned(784, 10), 1600 => to_unsigned(103, 10), 1601 => to_unsigned(781, 10), 1602 => to_unsigned(993, 10), 1603 => to_unsigned(880, 10), 1604 => to_unsigned(552, 10), 1605 => to_unsigned(353, 10), 1606 => to_unsigned(623, 10), 1607 => to_unsigned(437, 10), 1608 => to_unsigned(107, 10), 1609 => to_unsigned(941, 10), 1610 => to_unsigned(915, 10), 1611 => to_unsigned(890, 10), 1612 => to_unsigned(652, 10), 1613 => to_unsigned(9, 10), 1614 => to_unsigned(41, 10), 1615 => to_unsigned(272, 10), 1616 => to_unsigned(35, 10), 1617 => to_unsigned(325, 10), 1618 => to_unsigned(997, 10), 1619 => to_unsigned(929, 10), 1620 => to_unsigned(547, 10), 1621 => to_unsigned(453, 10), 1622 => to_unsigned(474, 10), 1623 => to_unsigned(93, 10), 1624 => to_unsigned(305, 10), 1625 => to_unsigned(288, 10), 1626 => to_unsigned(763, 10), 1627 => to_unsigned(430, 10), 1628 => to_unsigned(332, 10), 1629 => to_unsigned(419, 10), 1630 => to_unsigned(619, 10), 1631 => to_unsigned(813, 10), 1632 => to_unsigned(772, 10), 1633 => to_unsigned(891, 10), 1634 => to_unsigned(490, 10), 1635 => to_unsigned(773, 10), 1636 => to_unsigned(937, 10), 1637 => to_unsigned(345, 10), 1638 => to_unsigned(857, 10), 1639 => to_unsigned(182, 10), 1640 => to_unsigned(53, 10), 1641 => to_unsigned(3, 10), 1642 => to_unsigned(556, 10), 1643 => to_unsigned(539, 10), 1644 => to_unsigned(345, 10), 1645 => to_unsigned(300, 10), 1646 => to_unsigned(433, 10), 1647 => to_unsigned(681, 10), 1648 => to_unsigned(978, 10), 1649 => to_unsigned(970, 10), 1650 => to_unsigned(955, 10), 1651 => to_unsigned(602, 10), 1652 => to_unsigned(84, 10), 1653 => to_unsigned(736, 10), 1654 => to_unsigned(12, 10), 1655 => to_unsigned(337, 10), 1656 => to_unsigned(605, 10), 1657 => to_unsigned(329, 10), 1658 => to_unsigned(965, 10), 1659 => to_unsigned(194, 10), 1660 => to_unsigned(705, 10), 1661 => to_unsigned(696, 10), 1662 => to_unsigned(99, 10), 1663 => to_unsigned(787, 10), 1664 => to_unsigned(231, 10), 1665 => to_unsigned(148, 10), 1666 => to_unsigned(639, 10), 1667 => to_unsigned(293, 10), 1668 => to_unsigned(1014, 10), 1669 => to_unsigned(267, 10), 1670 => to_unsigned(658, 10), 1671 => to_unsigned(631, 10), 1672 => to_unsigned(802, 10), 1673 => to_unsigned(54, 10), 1674 => to_unsigned(665, 10), 1675 => to_unsigned(594, 10), 1676 => to_unsigned(362, 10), 1677 => to_unsigned(683, 10), 1678 => to_unsigned(941, 10), 1679 => to_unsigned(944, 10), 1680 => to_unsigned(649, 10), 1681 => to_unsigned(756, 10), 1682 => to_unsigned(539, 10), 1683 => to_unsigned(279, 10), 1684 => to_unsigned(769, 10), 1685 => to_unsigned(950, 10), 1686 => to_unsigned(915, 10), 1687 => to_unsigned(378, 10), 1688 => to_unsigned(774, 10), 1689 => to_unsigned(28, 10), 1690 => to_unsigned(92, 10), 1691 => to_unsigned(477, 10), 1692 => to_unsigned(95, 10), 1693 => to_unsigned(848, 10), 1694 => to_unsigned(305, 10), 1695 => to_unsigned(357, 10), 1696 => to_unsigned(623, 10), 1697 => to_unsigned(615, 10), 1698 => to_unsigned(100, 10), 1699 => to_unsigned(171, 10), 1700 => to_unsigned(31, 10), 1701 => to_unsigned(65, 10), 1702 => to_unsigned(250, 10), 1703 => to_unsigned(920, 10), 1704 => to_unsigned(34, 10), 1705 => to_unsigned(381, 10), 1706 => to_unsigned(100, 10), 1707 => to_unsigned(298, 10), 1708 => to_unsigned(203, 10), 1709 => to_unsigned(219, 10), 1710 => to_unsigned(241, 10), 1711 => to_unsigned(479, 10), 1712 => to_unsigned(680, 10), 1713 => to_unsigned(256, 10), 1714 => to_unsigned(707, 10), 1715 => to_unsigned(322, 10), 1716 => to_unsigned(66, 10), 1717 => to_unsigned(301, 10), 1718 => to_unsigned(209, 10), 1719 => to_unsigned(780, 10), 1720 => to_unsigned(1012, 10), 1721 => to_unsigned(359, 10), 1722 => to_unsigned(489, 10), 1723 => to_unsigned(343, 10), 1724 => to_unsigned(262, 10), 1725 => to_unsigned(86, 10), 1726 => to_unsigned(828, 10), 1727 => to_unsigned(639, 10), 1728 => to_unsigned(51, 10), 1729 => to_unsigned(568, 10), 1730 => to_unsigned(206, 10), 1731 => to_unsigned(941, 10), 1732 => to_unsigned(320, 10), 1733 => to_unsigned(124, 10), 1734 => to_unsigned(916, 10), 1735 => to_unsigned(292, 10), 1736 => to_unsigned(96, 10), 1737 => to_unsigned(740, 10), 1738 => to_unsigned(530, 10), 1739 => to_unsigned(946, 10), 1740 => to_unsigned(931, 10), 1741 => to_unsigned(793, 10), 1742 => to_unsigned(862, 10), 1743 => to_unsigned(479, 10), 1744 => to_unsigned(510, 10), 1745 => to_unsigned(699, 10), 1746 => to_unsigned(1021, 10), 1747 => to_unsigned(527, 10), 1748 => to_unsigned(728, 10), 1749 => to_unsigned(790, 10), 1750 => to_unsigned(834, 10), 1751 => to_unsigned(23, 10), 1752 => to_unsigned(161, 10), 1753 => to_unsigned(373, 10), 1754 => to_unsigned(874, 10), 1755 => to_unsigned(372, 10), 1756 => to_unsigned(456, 10), 1757 => to_unsigned(617, 10), 1758 => to_unsigned(431, 10), 1759 => to_unsigned(315, 10), 1760 => to_unsigned(365, 10), 1761 => to_unsigned(440, 10), 1762 => to_unsigned(463, 10), 1763 => to_unsigned(19, 10), 1764 => to_unsigned(78, 10), 1765 => to_unsigned(294, 10), 1766 => to_unsigned(37, 10), 1767 => to_unsigned(803, 10), 1768 => to_unsigned(267, 10), 1769 => to_unsigned(870, 10), 1770 => to_unsigned(668, 10), 1771 => to_unsigned(227, 10), 1772 => to_unsigned(810, 10), 1773 => to_unsigned(223, 10), 1774 => to_unsigned(685, 10), 1775 => to_unsigned(209, 10), 1776 => to_unsigned(553, 10), 1777 => to_unsigned(334, 10), 1778 => to_unsigned(552, 10), 1779 => to_unsigned(114, 10), 1780 => to_unsigned(931, 10), 1781 => to_unsigned(190, 10), 1782 => to_unsigned(421, 10), 1783 => to_unsigned(735, 10), 1784 => to_unsigned(567, 10), 1785 => to_unsigned(802, 10), 1786 => to_unsigned(750, 10), 1787 => to_unsigned(287, 10), 1788 => to_unsigned(467, 10), 1789 => to_unsigned(403, 10), 1790 => to_unsigned(313, 10), 1791 => to_unsigned(613, 10), 1792 => to_unsigned(23, 10), 1793 => to_unsigned(588, 10), 1794 => to_unsigned(238, 10), 1795 => to_unsigned(80, 10), 1796 => to_unsigned(865, 10), 1797 => to_unsigned(951, 10), 1798 => to_unsigned(542, 10), 1799 => to_unsigned(91, 10), 1800 => to_unsigned(504, 10), 1801 => to_unsigned(230, 10), 1802 => to_unsigned(387, 10), 1803 => to_unsigned(854, 10), 1804 => to_unsigned(385, 10), 1805 => to_unsigned(526, 10), 1806 => to_unsigned(923, 10), 1807 => to_unsigned(640, 10), 1808 => to_unsigned(747, 10), 1809 => to_unsigned(9, 10), 1810 => to_unsigned(291, 10), 1811 => to_unsigned(846, 10), 1812 => to_unsigned(544, 10), 1813 => to_unsigned(698, 10), 1814 => to_unsigned(666, 10), 1815 => to_unsigned(268, 10), 1816 => to_unsigned(820, 10), 1817 => to_unsigned(953, 10), 1818 => to_unsigned(173, 10), 1819 => to_unsigned(846, 10), 1820 => to_unsigned(19, 10), 1821 => to_unsigned(605, 10), 1822 => to_unsigned(1011, 10), 1823 => to_unsigned(374, 10), 1824 => to_unsigned(891, 10), 1825 => to_unsigned(849, 10), 1826 => to_unsigned(70, 10), 1827 => to_unsigned(239, 10), 1828 => to_unsigned(161, 10), 1829 => to_unsigned(205, 10), 1830 => to_unsigned(214, 10), 1831 => to_unsigned(299, 10), 1832 => to_unsigned(768, 10), 1833 => to_unsigned(57, 10), 1834 => to_unsigned(662, 10), 1835 => to_unsigned(238, 10), 1836 => to_unsigned(782, 10), 1837 => to_unsigned(868, 10), 1838 => to_unsigned(504, 10), 1839 => to_unsigned(581, 10), 1840 => to_unsigned(266, 10), 1841 => to_unsigned(67, 10), 1842 => to_unsigned(4, 10), 1843 => to_unsigned(180, 10), 1844 => to_unsigned(60, 10), 1845 => to_unsigned(308, 10), 1846 => to_unsigned(959, 10), 1847 => to_unsigned(734, 10), 1848 => to_unsigned(389, 10), 1849 => to_unsigned(523, 10), 1850 => to_unsigned(60, 10), 1851 => to_unsigned(141, 10), 1852 => to_unsigned(652, 10), 1853 => to_unsigned(903, 10), 1854 => to_unsigned(312, 10), 1855 => to_unsigned(389, 10), 1856 => to_unsigned(825, 10), 1857 => to_unsigned(906, 10), 1858 => to_unsigned(414, 10), 1859 => to_unsigned(387, 10), 1860 => to_unsigned(738, 10), 1861 => to_unsigned(378, 10), 1862 => to_unsigned(317, 10), 1863 => to_unsigned(641, 10), 1864 => to_unsigned(811, 10), 1865 => to_unsigned(400, 10), 1866 => to_unsigned(935, 10), 1867 => to_unsigned(913, 10), 1868 => to_unsigned(564, 10), 1869 => to_unsigned(1006, 10), 1870 => to_unsigned(436, 10), 1871 => to_unsigned(634, 10), 1872 => to_unsigned(880, 10), 1873 => to_unsigned(519, 10), 1874 => to_unsigned(146, 10), 1875 => to_unsigned(405, 10), 1876 => to_unsigned(662, 10), 1877 => to_unsigned(798, 10), 1878 => to_unsigned(324, 10), 1879 => to_unsigned(863, 10), 1880 => to_unsigned(387, 10), 1881 => to_unsigned(689, 10), 1882 => to_unsigned(752, 10), 1883 => to_unsigned(137, 10), 1884 => to_unsigned(137, 10), 1885 => to_unsigned(674, 10), 1886 => to_unsigned(742, 10), 1887 => to_unsigned(247, 10), 1888 => to_unsigned(862, 10), 1889 => to_unsigned(76, 10), 1890 => to_unsigned(432, 10), 1891 => to_unsigned(945, 10), 1892 => to_unsigned(136, 10), 1893 => to_unsigned(895, 10), 1894 => to_unsigned(1015, 10), 1895 => to_unsigned(238, 10), 1896 => to_unsigned(24, 10), 1897 => to_unsigned(164, 10), 1898 => to_unsigned(119, 10), 1899 => to_unsigned(265, 10), 1900 => to_unsigned(6, 10), 1901 => to_unsigned(776, 10), 1902 => to_unsigned(760, 10), 1903 => to_unsigned(81, 10), 1904 => to_unsigned(329, 10), 1905 => to_unsigned(953, 10), 1906 => to_unsigned(890, 10), 1907 => to_unsigned(129, 10), 1908 => to_unsigned(676, 10), 1909 => to_unsigned(0, 10), 1910 => to_unsigned(570, 10), 1911 => to_unsigned(297, 10), 1912 => to_unsigned(718, 10), 1913 => to_unsigned(566, 10), 1914 => to_unsigned(475, 10), 1915 => to_unsigned(538, 10), 1916 => to_unsigned(674, 10), 1917 => to_unsigned(197, 10), 1918 => to_unsigned(126, 10), 1919 => to_unsigned(7, 10), 1920 => to_unsigned(754, 10), 1921 => to_unsigned(210, 10), 1922 => to_unsigned(248, 10), 1923 => to_unsigned(911, 10), 1924 => to_unsigned(157, 10), 1925 => to_unsigned(511, 10), 1926 => to_unsigned(230, 10), 1927 => to_unsigned(208, 10), 1928 => to_unsigned(829, 10), 1929 => to_unsigned(562, 10), 1930 => to_unsigned(771, 10), 1931 => to_unsigned(689, 10), 1932 => to_unsigned(453, 10), 1933 => to_unsigned(485, 10), 1934 => to_unsigned(602, 10), 1935 => to_unsigned(674, 10), 1936 => to_unsigned(353, 10), 1937 => to_unsigned(216, 10), 1938 => to_unsigned(437, 10), 1939 => to_unsigned(298, 10), 1940 => to_unsigned(674, 10), 1941 => to_unsigned(202, 10), 1942 => to_unsigned(834, 10), 1943 => to_unsigned(577, 10), 1944 => to_unsigned(960, 10), 1945 => to_unsigned(939, 10), 1946 => to_unsigned(505, 10), 1947 => to_unsigned(267, 10), 1948 => to_unsigned(886, 10), 1949 => to_unsigned(839, 10), 1950 => to_unsigned(419, 10), 1951 => to_unsigned(657, 10), 1952 => to_unsigned(872, 10), 1953 => to_unsigned(456, 10), 1954 => to_unsigned(37, 10), 1955 => to_unsigned(288, 10), 1956 => to_unsigned(193, 10), 1957 => to_unsigned(617, 10), 1958 => to_unsigned(516, 10), 1959 => to_unsigned(750, 10), 1960 => to_unsigned(209, 10), 1961 => to_unsigned(476, 10), 1962 => to_unsigned(443, 10), 1963 => to_unsigned(863, 10), 1964 => to_unsigned(209, 10), 1965 => to_unsigned(164, 10), 1966 => to_unsigned(448, 10), 1967 => to_unsigned(237, 10), 1968 => to_unsigned(83, 10), 1969 => to_unsigned(281, 10), 1970 => to_unsigned(29, 10), 1971 => to_unsigned(255, 10), 1972 => to_unsigned(263, 10), 1973 => to_unsigned(602, 10), 1974 => to_unsigned(390, 10), 1975 => to_unsigned(159, 10), 1976 => to_unsigned(443, 10), 1977 => to_unsigned(1005, 10), 1978 => to_unsigned(67, 10), 1979 => to_unsigned(260, 10), 1980 => to_unsigned(769, 10), 1981 => to_unsigned(588, 10), 1982 => to_unsigned(1011, 10), 1983 => to_unsigned(648, 10), 1984 => to_unsigned(831, 10), 1985 => to_unsigned(289, 10), 1986 => to_unsigned(161, 10), 1987 => to_unsigned(375, 10), 1988 => to_unsigned(29, 10), 1989 => to_unsigned(925, 10), 1990 => to_unsigned(726, 10), 1991 => to_unsigned(831, 10), 1992 => to_unsigned(409, 10), 1993 => to_unsigned(93, 10), 1994 => to_unsigned(568, 10), 1995 => to_unsigned(195, 10), 1996 => to_unsigned(362, 10), 1997 => to_unsigned(347, 10), 1998 => to_unsigned(296, 10), 1999 => to_unsigned(756, 10), 2000 => to_unsigned(108, 10), 2001 => to_unsigned(269, 10), 2002 => to_unsigned(90, 10), 2003 => to_unsigned(172, 10), 2004 => to_unsigned(536, 10), 2005 => to_unsigned(354, 10), 2006 => to_unsigned(176, 10), 2007 => to_unsigned(665, 10), 2008 => to_unsigned(700, 10), 2009 => to_unsigned(421, 10), 2010 => to_unsigned(503, 10), 2011 => to_unsigned(31, 10), 2012 => to_unsigned(527, 10), 2013 => to_unsigned(214, 10), 2014 => to_unsigned(481, 10), 2015 => to_unsigned(139, 10), 2016 => to_unsigned(998, 10), 2017 => to_unsigned(998, 10), 2018 => to_unsigned(145, 10), 2019 => to_unsigned(284, 10), 2020 => to_unsigned(299, 10), 2021 => to_unsigned(639, 10), 2022 => to_unsigned(788, 10), 2023 => to_unsigned(364, 10), 2024 => to_unsigned(36, 10), 2025 => to_unsigned(264, 10), 2026 => to_unsigned(303, 10), 2027 => to_unsigned(773, 10), 2028 => to_unsigned(542, 10), 2029 => to_unsigned(700, 10), 2030 => to_unsigned(947, 10), 2031 => to_unsigned(175, 10), 2032 => to_unsigned(819, 10), 2033 => to_unsigned(514, 10), 2034 => to_unsigned(212, 10), 2035 => to_unsigned(856, 10), 2036 => to_unsigned(492, 10), 2037 => to_unsigned(909, 10), 2038 => to_unsigned(702, 10), 2039 => to_unsigned(339, 10), 2040 => to_unsigned(545, 10), 2041 => to_unsigned(806, 10), 2042 => to_unsigned(988, 10), 2043 => to_unsigned(80, 10), 2044 => to_unsigned(275, 10), 2045 => to_unsigned(676, 10), 2046 => to_unsigned(271, 10), 2047 => to_unsigned(677, 10)),
            5 => (0 => to_unsigned(118, 10), 1 => to_unsigned(870, 10), 2 => to_unsigned(266, 10), 3 => to_unsigned(745, 10), 4 => to_unsigned(502, 10), 5 => to_unsigned(307, 10), 6 => to_unsigned(1018, 10), 7 => to_unsigned(147, 10), 8 => to_unsigned(693, 10), 9 => to_unsigned(425, 10), 10 => to_unsigned(890, 10), 11 => to_unsigned(1002, 10), 12 => to_unsigned(777, 10), 13 => to_unsigned(973, 10), 14 => to_unsigned(73, 10), 15 => to_unsigned(669, 10), 16 => to_unsigned(65, 10), 17 => to_unsigned(891, 10), 18 => to_unsigned(373, 10), 19 => to_unsigned(311, 10), 20 => to_unsigned(83, 10), 21 => to_unsigned(96, 10), 22 => to_unsigned(418, 10), 23 => to_unsigned(570, 10), 24 => to_unsigned(158, 10), 25 => to_unsigned(949, 10), 26 => to_unsigned(804, 10), 27 => to_unsigned(410, 10), 28 => to_unsigned(680, 10), 29 => to_unsigned(128, 10), 30 => to_unsigned(401, 10), 31 => to_unsigned(826, 10), 32 => to_unsigned(479, 10), 33 => to_unsigned(983, 10), 34 => to_unsigned(32, 10), 35 => to_unsigned(17, 10), 36 => to_unsigned(455, 10), 37 => to_unsigned(263, 10), 38 => to_unsigned(374, 10), 39 => to_unsigned(949, 10), 40 => to_unsigned(656, 10), 41 => to_unsigned(639, 10), 42 => to_unsigned(874, 10), 43 => to_unsigned(30, 10), 44 => to_unsigned(286, 10), 45 => to_unsigned(502, 10), 46 => to_unsigned(930, 10), 47 => to_unsigned(409, 10), 48 => to_unsigned(850, 10), 49 => to_unsigned(713, 10), 50 => to_unsigned(978, 10), 51 => to_unsigned(660, 10), 52 => to_unsigned(185, 10), 53 => to_unsigned(204, 10), 54 => to_unsigned(783, 10), 55 => to_unsigned(725, 10), 56 => to_unsigned(682, 10), 57 => to_unsigned(678, 10), 58 => to_unsigned(405, 10), 59 => to_unsigned(139, 10), 60 => to_unsigned(242, 10), 61 => to_unsigned(325, 10), 62 => to_unsigned(85, 10), 63 => to_unsigned(118, 10), 64 => to_unsigned(470, 10), 65 => to_unsigned(107, 10), 66 => to_unsigned(474, 10), 67 => to_unsigned(913, 10), 68 => to_unsigned(968, 10), 69 => to_unsigned(785, 10), 70 => to_unsigned(661, 10), 71 => to_unsigned(819, 10), 72 => to_unsigned(258, 10), 73 => to_unsigned(570, 10), 74 => to_unsigned(1007, 10), 75 => to_unsigned(954, 10), 76 => to_unsigned(560, 10), 77 => to_unsigned(496, 10), 78 => to_unsigned(553, 10), 79 => to_unsigned(797, 10), 80 => to_unsigned(729, 10), 81 => to_unsigned(979, 10), 82 => to_unsigned(864, 10), 83 => to_unsigned(76, 10), 84 => to_unsigned(561, 10), 85 => to_unsigned(687, 10), 86 => to_unsigned(117, 10), 87 => to_unsigned(550, 10), 88 => to_unsigned(812, 10), 89 => to_unsigned(593, 10), 90 => to_unsigned(383, 10), 91 => to_unsigned(669, 10), 92 => to_unsigned(324, 10), 93 => to_unsigned(918, 10), 94 => to_unsigned(206, 10), 95 => to_unsigned(164, 10), 96 => to_unsigned(177, 10), 97 => to_unsigned(464, 10), 98 => to_unsigned(79, 10), 99 => to_unsigned(415, 10), 100 => to_unsigned(913, 10), 101 => to_unsigned(64, 10), 102 => to_unsigned(527, 10), 103 => to_unsigned(450, 10), 104 => to_unsigned(861, 10), 105 => to_unsigned(871, 10), 106 => to_unsigned(941, 10), 107 => to_unsigned(186, 10), 108 => to_unsigned(802, 10), 109 => to_unsigned(894, 10), 110 => to_unsigned(77, 10), 111 => to_unsigned(434, 10), 112 => to_unsigned(123, 10), 113 => to_unsigned(734, 10), 114 => to_unsigned(963, 10), 115 => to_unsigned(353, 10), 116 => to_unsigned(822, 10), 117 => to_unsigned(116, 10), 118 => to_unsigned(227, 10), 119 => to_unsigned(315, 10), 120 => to_unsigned(636, 10), 121 => to_unsigned(403, 10), 122 => to_unsigned(4, 10), 123 => to_unsigned(203, 10), 124 => to_unsigned(178, 10), 125 => to_unsigned(933, 10), 126 => to_unsigned(590, 10), 127 => to_unsigned(175, 10), 128 => to_unsigned(460, 10), 129 => to_unsigned(870, 10), 130 => to_unsigned(682, 10), 131 => to_unsigned(817, 10), 132 => to_unsigned(540, 10), 133 => to_unsigned(596, 10), 134 => to_unsigned(224, 10), 135 => to_unsigned(875, 10), 136 => to_unsigned(902, 10), 137 => to_unsigned(636, 10), 138 => to_unsigned(462, 10), 139 => to_unsigned(752, 10), 140 => to_unsigned(229, 10), 141 => to_unsigned(440, 10), 142 => to_unsigned(312, 10), 143 => to_unsigned(685, 10), 144 => to_unsigned(770, 10), 145 => to_unsigned(1016, 10), 146 => to_unsigned(948, 10), 147 => to_unsigned(841, 10), 148 => to_unsigned(539, 10), 149 => to_unsigned(879, 10), 150 => to_unsigned(861, 10), 151 => to_unsigned(290, 10), 152 => to_unsigned(901, 10), 153 => to_unsigned(312, 10), 154 => to_unsigned(280, 10), 155 => to_unsigned(170, 10), 156 => to_unsigned(557, 10), 157 => to_unsigned(202, 10), 158 => to_unsigned(493, 10), 159 => to_unsigned(524, 10), 160 => to_unsigned(4, 10), 161 => to_unsigned(758, 10), 162 => to_unsigned(737, 10), 163 => to_unsigned(100, 10), 164 => to_unsigned(676, 10), 165 => to_unsigned(93, 10), 166 => to_unsigned(678, 10), 167 => to_unsigned(330, 10), 168 => to_unsigned(554, 10), 169 => to_unsigned(803, 10), 170 => to_unsigned(866, 10), 171 => to_unsigned(570, 10), 172 => to_unsigned(716, 10), 173 => to_unsigned(533, 10), 174 => to_unsigned(582, 10), 175 => to_unsigned(479, 10), 176 => to_unsigned(652, 10), 177 => to_unsigned(298, 10), 178 => to_unsigned(706, 10), 179 => to_unsigned(947, 10), 180 => to_unsigned(151, 10), 181 => to_unsigned(920, 10), 182 => to_unsigned(383, 10), 183 => to_unsigned(842, 10), 184 => to_unsigned(241, 10), 185 => to_unsigned(715, 10), 186 => to_unsigned(54, 10), 187 => to_unsigned(104, 10), 188 => to_unsigned(437, 10), 189 => to_unsigned(964, 10), 190 => to_unsigned(226, 10), 191 => to_unsigned(593, 10), 192 => to_unsigned(580, 10), 193 => to_unsigned(154, 10), 194 => to_unsigned(552, 10), 195 => to_unsigned(775, 10), 196 => to_unsigned(130, 10), 197 => to_unsigned(1013, 10), 198 => to_unsigned(98, 10), 199 => to_unsigned(97, 10), 200 => to_unsigned(171, 10), 201 => to_unsigned(468, 10), 202 => to_unsigned(285, 10), 203 => to_unsigned(748, 10), 204 => to_unsigned(834, 10), 205 => to_unsigned(462, 10), 206 => to_unsigned(753, 10), 207 => to_unsigned(883, 10), 208 => to_unsigned(202, 10), 209 => to_unsigned(204, 10), 210 => to_unsigned(474, 10), 211 => to_unsigned(814, 10), 212 => to_unsigned(935, 10), 213 => to_unsigned(880, 10), 214 => to_unsigned(309, 10), 215 => to_unsigned(1014, 10), 216 => to_unsigned(14, 10), 217 => to_unsigned(158, 10), 218 => to_unsigned(963, 10), 219 => to_unsigned(718, 10), 220 => to_unsigned(1002, 10), 221 => to_unsigned(241, 10), 222 => to_unsigned(917, 10), 223 => to_unsigned(932, 10), 224 => to_unsigned(69, 10), 225 => to_unsigned(424, 10), 226 => to_unsigned(241, 10), 227 => to_unsigned(620, 10), 228 => to_unsigned(144, 10), 229 => to_unsigned(766, 10), 230 => to_unsigned(775, 10), 231 => to_unsigned(980, 10), 232 => to_unsigned(659, 10), 233 => to_unsigned(258, 10), 234 => to_unsigned(316, 10), 235 => to_unsigned(672, 10), 236 => to_unsigned(611, 10), 237 => to_unsigned(658, 10), 238 => to_unsigned(51, 10), 239 => to_unsigned(559, 10), 240 => to_unsigned(889, 10), 241 => to_unsigned(573, 10), 242 => to_unsigned(913, 10), 243 => to_unsigned(834, 10), 244 => to_unsigned(694, 10), 245 => to_unsigned(777, 10), 246 => to_unsigned(682, 10), 247 => to_unsigned(326, 10), 248 => to_unsigned(21, 10), 249 => to_unsigned(433, 10), 250 => to_unsigned(301, 10), 251 => to_unsigned(263, 10), 252 => to_unsigned(469, 10), 253 => to_unsigned(585, 10), 254 => to_unsigned(111, 10), 255 => to_unsigned(729, 10), 256 => to_unsigned(914, 10), 257 => to_unsigned(502, 10), 258 => to_unsigned(444, 10), 259 => to_unsigned(711, 10), 260 => to_unsigned(974, 10), 261 => to_unsigned(260, 10), 262 => to_unsigned(113, 10), 263 => to_unsigned(988, 10), 264 => to_unsigned(211, 10), 265 => to_unsigned(713, 10), 266 => to_unsigned(731, 10), 267 => to_unsigned(660, 10), 268 => to_unsigned(962, 10), 269 => to_unsigned(781, 10), 270 => to_unsigned(445, 10), 271 => to_unsigned(886, 10), 272 => to_unsigned(224, 10), 273 => to_unsigned(655, 10), 274 => to_unsigned(634, 10), 275 => to_unsigned(690, 10), 276 => to_unsigned(53, 10), 277 => to_unsigned(837, 10), 278 => to_unsigned(716, 10), 279 => to_unsigned(170, 10), 280 => to_unsigned(933, 10), 281 => to_unsigned(645, 10), 282 => to_unsigned(820, 10), 283 => to_unsigned(624, 10), 284 => to_unsigned(572, 10), 285 => to_unsigned(827, 10), 286 => to_unsigned(798, 10), 287 => to_unsigned(135, 10), 288 => to_unsigned(212, 10), 289 => to_unsigned(851, 10), 290 => to_unsigned(290, 10), 291 => to_unsigned(538, 10), 292 => to_unsigned(295, 10), 293 => to_unsigned(971, 10), 294 => to_unsigned(594, 10), 295 => to_unsigned(657, 10), 296 => to_unsigned(383, 10), 297 => to_unsigned(704, 10), 298 => to_unsigned(110, 10), 299 => to_unsigned(701, 10), 300 => to_unsigned(566, 10), 301 => to_unsigned(644, 10), 302 => to_unsigned(976, 10), 303 => to_unsigned(1002, 10), 304 => to_unsigned(56, 10), 305 => to_unsigned(729, 10), 306 => to_unsigned(737, 10), 307 => to_unsigned(412, 10), 308 => to_unsigned(378, 10), 309 => to_unsigned(366, 10), 310 => to_unsigned(226, 10), 311 => to_unsigned(913, 10), 312 => to_unsigned(135, 10), 313 => to_unsigned(171, 10), 314 => to_unsigned(192, 10), 315 => to_unsigned(305, 10), 316 => to_unsigned(456, 10), 317 => to_unsigned(468, 10), 318 => to_unsigned(513, 10), 319 => to_unsigned(741, 10), 320 => to_unsigned(508, 10), 321 => to_unsigned(667, 10), 322 => to_unsigned(171, 10), 323 => to_unsigned(314, 10), 324 => to_unsigned(783, 10), 325 => to_unsigned(948, 10), 326 => to_unsigned(521, 10), 327 => to_unsigned(792, 10), 328 => to_unsigned(968, 10), 329 => to_unsigned(876, 10), 330 => to_unsigned(89, 10), 331 => to_unsigned(754, 10), 332 => to_unsigned(995, 10), 333 => to_unsigned(686, 10), 334 => to_unsigned(475, 10), 335 => to_unsigned(354, 10), 336 => to_unsigned(45, 10), 337 => to_unsigned(577, 10), 338 => to_unsigned(950, 10), 339 => to_unsigned(200, 10), 340 => to_unsigned(719, 10), 341 => to_unsigned(664, 10), 342 => to_unsigned(125, 10), 343 => to_unsigned(629, 10), 344 => to_unsigned(8, 10), 345 => to_unsigned(913, 10), 346 => to_unsigned(633, 10), 347 => to_unsigned(295, 10), 348 => to_unsigned(596, 10), 349 => to_unsigned(6, 10), 350 => to_unsigned(228, 10), 351 => to_unsigned(302, 10), 352 => to_unsigned(978, 10), 353 => to_unsigned(666, 10), 354 => to_unsigned(240, 10), 355 => to_unsigned(591, 10), 356 => to_unsigned(7, 10), 357 => to_unsigned(385, 10), 358 => to_unsigned(284, 10), 359 => to_unsigned(272, 10), 360 => to_unsigned(157, 10), 361 => to_unsigned(844, 10), 362 => to_unsigned(353, 10), 363 => to_unsigned(129, 10), 364 => to_unsigned(498, 10), 365 => to_unsigned(669, 10), 366 => to_unsigned(174, 10), 367 => to_unsigned(606, 10), 368 => to_unsigned(977, 10), 369 => to_unsigned(369, 10), 370 => to_unsigned(389, 10), 371 => to_unsigned(405, 10), 372 => to_unsigned(901, 10), 373 => to_unsigned(1015, 10), 374 => to_unsigned(600, 10), 375 => to_unsigned(1001, 10), 376 => to_unsigned(399, 10), 377 => to_unsigned(310, 10), 378 => to_unsigned(999, 10), 379 => to_unsigned(1003, 10), 380 => to_unsigned(872, 10), 381 => to_unsigned(301, 10), 382 => to_unsigned(599, 10), 383 => to_unsigned(559, 10), 384 => to_unsigned(469, 10), 385 => to_unsigned(42, 10), 386 => to_unsigned(150, 10), 387 => to_unsigned(744, 10), 388 => to_unsigned(32, 10), 389 => to_unsigned(969, 10), 390 => to_unsigned(360, 10), 391 => to_unsigned(220, 10), 392 => to_unsigned(571, 10), 393 => to_unsigned(303, 10), 394 => to_unsigned(877, 10), 395 => to_unsigned(668, 10), 396 => to_unsigned(650, 10), 397 => to_unsigned(789, 10), 398 => to_unsigned(715, 10), 399 => to_unsigned(377, 10), 400 => to_unsigned(403, 10), 401 => to_unsigned(847, 10), 402 => to_unsigned(137, 10), 403 => to_unsigned(24, 10), 404 => to_unsigned(305, 10), 405 => to_unsigned(818, 10), 406 => to_unsigned(436, 10), 407 => to_unsigned(979, 10), 408 => to_unsigned(270, 10), 409 => to_unsigned(356, 10), 410 => to_unsigned(287, 10), 411 => to_unsigned(966, 10), 412 => to_unsigned(357, 10), 413 => to_unsigned(797, 10), 414 => to_unsigned(228, 10), 415 => to_unsigned(933, 10), 416 => to_unsigned(636, 10), 417 => to_unsigned(173, 10), 418 => to_unsigned(988, 10), 419 => to_unsigned(80, 10), 420 => to_unsigned(570, 10), 421 => to_unsigned(261, 10), 422 => to_unsigned(594, 10), 423 => to_unsigned(689, 10), 424 => to_unsigned(209, 10), 425 => to_unsigned(161, 10), 426 => to_unsigned(474, 10), 427 => to_unsigned(983, 10), 428 => to_unsigned(106, 10), 429 => to_unsigned(306, 10), 430 => to_unsigned(505, 10), 431 => to_unsigned(16, 10), 432 => to_unsigned(597, 10), 433 => to_unsigned(301, 10), 434 => to_unsigned(428, 10), 435 => to_unsigned(149, 10), 436 => to_unsigned(431, 10), 437 => to_unsigned(794, 10), 438 => to_unsigned(46, 10), 439 => to_unsigned(370, 10), 440 => to_unsigned(491, 10), 441 => to_unsigned(730, 10), 442 => to_unsigned(260, 10), 443 => to_unsigned(550, 10), 444 => to_unsigned(333, 10), 445 => to_unsigned(585, 10), 446 => to_unsigned(326, 10), 447 => to_unsigned(291, 10), 448 => to_unsigned(12, 10), 449 => to_unsigned(645, 10), 450 => to_unsigned(991, 10), 451 => to_unsigned(56, 10), 452 => to_unsigned(796, 10), 453 => to_unsigned(210, 10), 454 => to_unsigned(958, 10), 455 => to_unsigned(729, 10), 456 => to_unsigned(988, 10), 457 => to_unsigned(227, 10), 458 => to_unsigned(876, 10), 459 => to_unsigned(15, 10), 460 => to_unsigned(351, 10), 461 => to_unsigned(943, 10), 462 => to_unsigned(291, 10), 463 => to_unsigned(507, 10), 464 => to_unsigned(766, 10), 465 => to_unsigned(732, 10), 466 => to_unsigned(607, 10), 467 => to_unsigned(139, 10), 468 => to_unsigned(153, 10), 469 => to_unsigned(530, 10), 470 => to_unsigned(608, 10), 471 => to_unsigned(60, 10), 472 => to_unsigned(483, 10), 473 => to_unsigned(90, 10), 474 => to_unsigned(819, 10), 475 => to_unsigned(890, 10), 476 => to_unsigned(478, 10), 477 => to_unsigned(68, 10), 478 => to_unsigned(939, 10), 479 => to_unsigned(270, 10), 480 => to_unsigned(261, 10), 481 => to_unsigned(992, 10), 482 => to_unsigned(128, 10), 483 => to_unsigned(174, 10), 484 => to_unsigned(260, 10), 485 => to_unsigned(829, 10), 486 => to_unsigned(789, 10), 487 => to_unsigned(763, 10), 488 => to_unsigned(212, 10), 489 => to_unsigned(562, 10), 490 => to_unsigned(383, 10), 491 => to_unsigned(111, 10), 492 => to_unsigned(615, 10), 493 => to_unsigned(14, 10), 494 => to_unsigned(183, 10), 495 => to_unsigned(709, 10), 496 => to_unsigned(396, 10), 497 => to_unsigned(624, 10), 498 => to_unsigned(441, 10), 499 => to_unsigned(515, 10), 500 => to_unsigned(797, 10), 501 => to_unsigned(801, 10), 502 => to_unsigned(816, 10), 503 => to_unsigned(889, 10), 504 => to_unsigned(677, 10), 505 => to_unsigned(786, 10), 506 => to_unsigned(201, 10), 507 => to_unsigned(164, 10), 508 => to_unsigned(624, 10), 509 => to_unsigned(67, 10), 510 => to_unsigned(752, 10), 511 => to_unsigned(133, 10), 512 => to_unsigned(956, 10), 513 => to_unsigned(575, 10), 514 => to_unsigned(200, 10), 515 => to_unsigned(713, 10), 516 => to_unsigned(401, 10), 517 => to_unsigned(362, 10), 518 => to_unsigned(870, 10), 519 => to_unsigned(111, 10), 520 => to_unsigned(471, 10), 521 => to_unsigned(876, 10), 522 => to_unsigned(1012, 10), 523 => to_unsigned(451, 10), 524 => to_unsigned(615, 10), 525 => to_unsigned(515, 10), 526 => to_unsigned(747, 10), 527 => to_unsigned(581, 10), 528 => to_unsigned(684, 10), 529 => to_unsigned(506, 10), 530 => to_unsigned(459, 10), 531 => to_unsigned(553, 10), 532 => to_unsigned(958, 10), 533 => to_unsigned(299, 10), 534 => to_unsigned(891, 10), 535 => to_unsigned(996, 10), 536 => to_unsigned(79, 10), 537 => to_unsigned(862, 10), 538 => to_unsigned(384, 10), 539 => to_unsigned(656, 10), 540 => to_unsigned(502, 10), 541 => to_unsigned(161, 10), 542 => to_unsigned(173, 10), 543 => to_unsigned(555, 10), 544 => to_unsigned(583, 10), 545 => to_unsigned(81, 10), 546 => to_unsigned(421, 10), 547 => to_unsigned(169, 10), 548 => to_unsigned(294, 10), 549 => to_unsigned(35, 10), 550 => to_unsigned(305, 10), 551 => to_unsigned(209, 10), 552 => to_unsigned(527, 10), 553 => to_unsigned(54, 10), 554 => to_unsigned(554, 10), 555 => to_unsigned(345, 10), 556 => to_unsigned(328, 10), 557 => to_unsigned(685, 10), 558 => to_unsigned(941, 10), 559 => to_unsigned(143, 10), 560 => to_unsigned(958, 10), 561 => to_unsigned(239, 10), 562 => to_unsigned(122, 10), 563 => to_unsigned(564, 10), 564 => to_unsigned(363, 10), 565 => to_unsigned(740, 10), 566 => to_unsigned(291, 10), 567 => to_unsigned(610, 10), 568 => to_unsigned(108, 10), 569 => to_unsigned(824, 10), 570 => to_unsigned(897, 10), 571 => to_unsigned(1014, 10), 572 => to_unsigned(739, 10), 573 => to_unsigned(951, 10), 574 => to_unsigned(92, 10), 575 => to_unsigned(539, 10), 576 => to_unsigned(253, 10), 577 => to_unsigned(895, 10), 578 => to_unsigned(169, 10), 579 => to_unsigned(242, 10), 580 => to_unsigned(514, 10), 581 => to_unsigned(142, 10), 582 => to_unsigned(280, 10), 583 => to_unsigned(984, 10), 584 => to_unsigned(490, 10), 585 => to_unsigned(1023, 10), 586 => to_unsigned(19, 10), 587 => to_unsigned(901, 10), 588 => to_unsigned(99, 10), 589 => to_unsigned(123, 10), 590 => to_unsigned(291, 10), 591 => to_unsigned(929, 10), 592 => to_unsigned(218, 10), 593 => to_unsigned(204, 10), 594 => to_unsigned(666, 10), 595 => to_unsigned(878, 10), 596 => to_unsigned(783, 10), 597 => to_unsigned(424, 10), 598 => to_unsigned(101, 10), 599 => to_unsigned(15, 10), 600 => to_unsigned(931, 10), 601 => to_unsigned(853, 10), 602 => to_unsigned(925, 10), 603 => to_unsigned(150, 10), 604 => to_unsigned(698, 10), 605 => to_unsigned(123, 10), 606 => to_unsigned(941, 10), 607 => to_unsigned(742, 10), 608 => to_unsigned(3, 10), 609 => to_unsigned(601, 10), 610 => to_unsigned(847, 10), 611 => to_unsigned(217, 10), 612 => to_unsigned(707, 10), 613 => to_unsigned(58, 10), 614 => to_unsigned(237, 10), 615 => to_unsigned(916, 10), 616 => to_unsigned(953, 10), 617 => to_unsigned(188, 10), 618 => to_unsigned(748, 10), 619 => to_unsigned(279, 10), 620 => to_unsigned(643, 10), 621 => to_unsigned(855, 10), 622 => to_unsigned(865, 10), 623 => to_unsigned(963, 10), 624 => to_unsigned(649, 10), 625 => to_unsigned(414, 10), 626 => to_unsigned(399, 10), 627 => to_unsigned(640, 10), 628 => to_unsigned(463, 10), 629 => to_unsigned(935, 10), 630 => to_unsigned(282, 10), 631 => to_unsigned(573, 10), 632 => to_unsigned(472, 10), 633 => to_unsigned(431, 10), 634 => to_unsigned(317, 10), 635 => to_unsigned(602, 10), 636 => to_unsigned(626, 10), 637 => to_unsigned(2, 10), 638 => to_unsigned(201, 10), 639 => to_unsigned(377, 10), 640 => to_unsigned(674, 10), 641 => to_unsigned(800, 10), 642 => to_unsigned(460, 10), 643 => to_unsigned(597, 10), 644 => to_unsigned(578, 10), 645 => to_unsigned(700, 10), 646 => to_unsigned(29, 10), 647 => to_unsigned(8, 10), 648 => to_unsigned(84, 10), 649 => to_unsigned(1017, 10), 650 => to_unsigned(736, 10), 651 => to_unsigned(57, 10), 652 => to_unsigned(156, 10), 653 => to_unsigned(419, 10), 654 => to_unsigned(256, 10), 655 => to_unsigned(949, 10), 656 => to_unsigned(750, 10), 657 => to_unsigned(243, 10), 658 => to_unsigned(714, 10), 659 => to_unsigned(387, 10), 660 => to_unsigned(110, 10), 661 => to_unsigned(321, 10), 662 => to_unsigned(409, 10), 663 => to_unsigned(396, 10), 664 => to_unsigned(572, 10), 665 => to_unsigned(74, 10), 666 => to_unsigned(697, 10), 667 => to_unsigned(496, 10), 668 => to_unsigned(406, 10), 669 => to_unsigned(877, 10), 670 => to_unsigned(733, 10), 671 => to_unsigned(586, 10), 672 => to_unsigned(315, 10), 673 => to_unsigned(56, 10), 674 => to_unsigned(50, 10), 675 => to_unsigned(111, 10), 676 => to_unsigned(579, 10), 677 => to_unsigned(759, 10), 678 => to_unsigned(288, 10), 679 => to_unsigned(804, 10), 680 => to_unsigned(457, 10), 681 => to_unsigned(115, 10), 682 => to_unsigned(225, 10), 683 => to_unsigned(291, 10), 684 => to_unsigned(489, 10), 685 => to_unsigned(517, 10), 686 => to_unsigned(222, 10), 687 => to_unsigned(171, 10), 688 => to_unsigned(97, 10), 689 => to_unsigned(965, 10), 690 => to_unsigned(284, 10), 691 => to_unsigned(393, 10), 692 => to_unsigned(101, 10), 693 => to_unsigned(766, 10), 694 => to_unsigned(875, 10), 695 => to_unsigned(829, 10), 696 => to_unsigned(109, 10), 697 => to_unsigned(94, 10), 698 => to_unsigned(479, 10), 699 => to_unsigned(57, 10), 700 => to_unsigned(449, 10), 701 => to_unsigned(146, 10), 702 => to_unsigned(766, 10), 703 => to_unsigned(183, 10), 704 => to_unsigned(963, 10), 705 => to_unsigned(901, 10), 706 => to_unsigned(721, 10), 707 => to_unsigned(166, 10), 708 => to_unsigned(155, 10), 709 => to_unsigned(746, 10), 710 => to_unsigned(263, 10), 711 => to_unsigned(247, 10), 712 => to_unsigned(491, 10), 713 => to_unsigned(747, 10), 714 => to_unsigned(118, 10), 715 => to_unsigned(699, 10), 716 => to_unsigned(872, 10), 717 => to_unsigned(991, 10), 718 => to_unsigned(761, 10), 719 => to_unsigned(246, 10), 720 => to_unsigned(224, 10), 721 => to_unsigned(865, 10), 722 => to_unsigned(745, 10), 723 => to_unsigned(730, 10), 724 => to_unsigned(688, 10), 725 => to_unsigned(670, 10), 726 => to_unsigned(88, 10), 727 => to_unsigned(359, 10), 728 => to_unsigned(556, 10), 729 => to_unsigned(698, 10), 730 => to_unsigned(437, 10), 731 => to_unsigned(849, 10), 732 => to_unsigned(721, 10), 733 => to_unsigned(556, 10), 734 => to_unsigned(161, 10), 735 => to_unsigned(824, 10), 736 => to_unsigned(645, 10), 737 => to_unsigned(430, 10), 738 => to_unsigned(262, 10), 739 => to_unsigned(231, 10), 740 => to_unsigned(988, 10), 741 => to_unsigned(148, 10), 742 => to_unsigned(897, 10), 743 => to_unsigned(721, 10), 744 => to_unsigned(583, 10), 745 => to_unsigned(548, 10), 746 => to_unsigned(917, 10), 747 => to_unsigned(360, 10), 748 => to_unsigned(553, 10), 749 => to_unsigned(169, 10), 750 => to_unsigned(916, 10), 751 => to_unsigned(830, 10), 752 => to_unsigned(714, 10), 753 => to_unsigned(519, 10), 754 => to_unsigned(951, 10), 755 => to_unsigned(829, 10), 756 => to_unsigned(72, 10), 757 => to_unsigned(881, 10), 758 => to_unsigned(981, 10), 759 => to_unsigned(438, 10), 760 => to_unsigned(439, 10), 761 => to_unsigned(662, 10), 762 => to_unsigned(271, 10), 763 => to_unsigned(217, 10), 764 => to_unsigned(426, 10), 765 => to_unsigned(545, 10), 766 => to_unsigned(739, 10), 767 => to_unsigned(166, 10), 768 => to_unsigned(885, 10), 769 => to_unsigned(286, 10), 770 => to_unsigned(876, 10), 771 => to_unsigned(297, 10), 772 => to_unsigned(333, 10), 773 => to_unsigned(470, 10), 774 => to_unsigned(675, 10), 775 => to_unsigned(585, 10), 776 => to_unsigned(364, 10), 777 => to_unsigned(987, 10), 778 => to_unsigned(763, 10), 779 => to_unsigned(926, 10), 780 => to_unsigned(268, 10), 781 => to_unsigned(62, 10), 782 => to_unsigned(654, 10), 783 => to_unsigned(482, 10), 784 => to_unsigned(511, 10), 785 => to_unsigned(994, 10), 786 => to_unsigned(716, 10), 787 => to_unsigned(361, 10), 788 => to_unsigned(624, 10), 789 => to_unsigned(353, 10), 790 => to_unsigned(331, 10), 791 => to_unsigned(248, 10), 792 => to_unsigned(699, 10), 793 => to_unsigned(987, 10), 794 => to_unsigned(566, 10), 795 => to_unsigned(726, 10), 796 => to_unsigned(868, 10), 797 => to_unsigned(181, 10), 798 => to_unsigned(1002, 10), 799 => to_unsigned(823, 10), 800 => to_unsigned(450, 10), 801 => to_unsigned(986, 10), 802 => to_unsigned(66, 10), 803 => to_unsigned(64, 10), 804 => to_unsigned(335, 10), 805 => to_unsigned(570, 10), 806 => to_unsigned(916, 10), 807 => to_unsigned(497, 10), 808 => to_unsigned(811, 10), 809 => to_unsigned(729, 10), 810 => to_unsigned(911, 10), 811 => to_unsigned(664, 10), 812 => to_unsigned(700, 10), 813 => to_unsigned(515, 10), 814 => to_unsigned(904, 10), 815 => to_unsigned(365, 10), 816 => to_unsigned(276, 10), 817 => to_unsigned(835, 10), 818 => to_unsigned(47, 10), 819 => to_unsigned(558, 10), 820 => to_unsigned(762, 10), 821 => to_unsigned(830, 10), 822 => to_unsigned(915, 10), 823 => to_unsigned(736, 10), 824 => to_unsigned(112, 10), 825 => to_unsigned(685, 10), 826 => to_unsigned(443, 10), 827 => to_unsigned(444, 10), 828 => to_unsigned(628, 10), 829 => to_unsigned(698, 10), 830 => to_unsigned(518, 10), 831 => to_unsigned(80, 10), 832 => to_unsigned(626, 10), 833 => to_unsigned(63, 10), 834 => to_unsigned(882, 10), 835 => to_unsigned(455, 10), 836 => to_unsigned(599, 10), 837 => to_unsigned(404, 10), 838 => to_unsigned(893, 10), 839 => to_unsigned(962, 10), 840 => to_unsigned(313, 10), 841 => to_unsigned(863, 10), 842 => to_unsigned(538, 10), 843 => to_unsigned(942, 10), 844 => to_unsigned(710, 10), 845 => to_unsigned(1002, 10), 846 => to_unsigned(205, 10), 847 => to_unsigned(816, 10), 848 => to_unsigned(699, 10), 849 => to_unsigned(186, 10), 850 => to_unsigned(562, 10), 851 => to_unsigned(350, 10), 852 => to_unsigned(102, 10), 853 => to_unsigned(235, 10), 854 => to_unsigned(568, 10), 855 => to_unsigned(509, 10), 856 => to_unsigned(357, 10), 857 => to_unsigned(557, 10), 858 => to_unsigned(816, 10), 859 => to_unsigned(637, 10), 860 => to_unsigned(225, 10), 861 => to_unsigned(407, 10), 862 => to_unsigned(68, 10), 863 => to_unsigned(840, 10), 864 => to_unsigned(784, 10), 865 => to_unsigned(118, 10), 866 => to_unsigned(769, 10), 867 => to_unsigned(179, 10), 868 => to_unsigned(685, 10), 869 => to_unsigned(592, 10), 870 => to_unsigned(294, 10), 871 => to_unsigned(496, 10), 872 => to_unsigned(506, 10), 873 => to_unsigned(260, 10), 874 => to_unsigned(627, 10), 875 => to_unsigned(794, 10), 876 => to_unsigned(748, 10), 877 => to_unsigned(75, 10), 878 => to_unsigned(773, 10), 879 => to_unsigned(372, 10), 880 => to_unsigned(166, 10), 881 => to_unsigned(491, 10), 882 => to_unsigned(670, 10), 883 => to_unsigned(24, 10), 884 => to_unsigned(971, 10), 885 => to_unsigned(45, 10), 886 => to_unsigned(145, 10), 887 => to_unsigned(485, 10), 888 => to_unsigned(709, 10), 889 => to_unsigned(695, 10), 890 => to_unsigned(318, 10), 891 => to_unsigned(90, 10), 892 => to_unsigned(409, 10), 893 => to_unsigned(781, 10), 894 => to_unsigned(276, 10), 895 => to_unsigned(125, 10), 896 => to_unsigned(516, 10), 897 => to_unsigned(207, 10), 898 => to_unsigned(1017, 10), 899 => to_unsigned(931, 10), 900 => to_unsigned(314, 10), 901 => to_unsigned(189, 10), 902 => to_unsigned(40, 10), 903 => to_unsigned(898, 10), 904 => to_unsigned(967, 10), 905 => to_unsigned(330, 10), 906 => to_unsigned(347, 10), 907 => to_unsigned(653, 10), 908 => to_unsigned(396, 10), 909 => to_unsigned(867, 10), 910 => to_unsigned(587, 10), 911 => to_unsigned(704, 10), 912 => to_unsigned(420, 10), 913 => to_unsigned(670, 10), 914 => to_unsigned(134, 10), 915 => to_unsigned(765, 10), 916 => to_unsigned(991, 10), 917 => to_unsigned(892, 10), 918 => to_unsigned(112, 10), 919 => to_unsigned(490, 10), 920 => to_unsigned(383, 10), 921 => to_unsigned(502, 10), 922 => to_unsigned(500, 10), 923 => to_unsigned(487, 10), 924 => to_unsigned(897, 10), 925 => to_unsigned(657, 10), 926 => to_unsigned(553, 10), 927 => to_unsigned(610, 10), 928 => to_unsigned(641, 10), 929 => to_unsigned(934, 10), 930 => to_unsigned(336, 10), 931 => to_unsigned(908, 10), 932 => to_unsigned(64, 10), 933 => to_unsigned(948, 10), 934 => to_unsigned(214, 10), 935 => to_unsigned(928, 10), 936 => to_unsigned(976, 10), 937 => to_unsigned(795, 10), 938 => to_unsigned(117, 10), 939 => to_unsigned(930, 10), 940 => to_unsigned(152, 10), 941 => to_unsigned(226, 10), 942 => to_unsigned(642, 10), 943 => to_unsigned(798, 10), 944 => to_unsigned(511, 10), 945 => to_unsigned(286, 10), 946 => to_unsigned(837, 10), 947 => to_unsigned(319, 10), 948 => to_unsigned(507, 10), 949 => to_unsigned(880, 10), 950 => to_unsigned(728, 10), 951 => to_unsigned(902, 10), 952 => to_unsigned(461, 10), 953 => to_unsigned(401, 10), 954 => to_unsigned(549, 10), 955 => to_unsigned(466, 10), 956 => to_unsigned(275, 10), 957 => to_unsigned(322, 10), 958 => to_unsigned(696, 10), 959 => to_unsigned(407, 10), 960 => to_unsigned(529, 10), 961 => to_unsigned(352, 10), 962 => to_unsigned(828, 10), 963 => to_unsigned(545, 10), 964 => to_unsigned(1003, 10), 965 => to_unsigned(435, 10), 966 => to_unsigned(786, 10), 967 => to_unsigned(426, 10), 968 => to_unsigned(609, 10), 969 => to_unsigned(968, 10), 970 => to_unsigned(809, 10), 971 => to_unsigned(972, 10), 972 => to_unsigned(493, 10), 973 => to_unsigned(129, 10), 974 => to_unsigned(989, 10), 975 => to_unsigned(953, 10), 976 => to_unsigned(110, 10), 977 => to_unsigned(1021, 10), 978 => to_unsigned(76, 10), 979 => to_unsigned(64, 10), 980 => to_unsigned(316, 10), 981 => to_unsigned(929, 10), 982 => to_unsigned(858, 10), 983 => to_unsigned(555, 10), 984 => to_unsigned(167, 10), 985 => to_unsigned(312, 10), 986 => to_unsigned(222, 10), 987 => to_unsigned(407, 10), 988 => to_unsigned(104, 10), 989 => to_unsigned(790, 10), 990 => to_unsigned(972, 10), 991 => to_unsigned(66, 10), 992 => to_unsigned(473, 10), 993 => to_unsigned(698, 10), 994 => to_unsigned(636, 10), 995 => to_unsigned(144, 10), 996 => to_unsigned(353, 10), 997 => to_unsigned(980, 10), 998 => to_unsigned(691, 10), 999 => to_unsigned(955, 10), 1000 => to_unsigned(115, 10), 1001 => to_unsigned(590, 10), 1002 => to_unsigned(901, 10), 1003 => to_unsigned(735, 10), 1004 => to_unsigned(47, 10), 1005 => to_unsigned(912, 10), 1006 => to_unsigned(896, 10), 1007 => to_unsigned(559, 10), 1008 => to_unsigned(506, 10), 1009 => to_unsigned(110, 10), 1010 => to_unsigned(22, 10), 1011 => to_unsigned(466, 10), 1012 => to_unsigned(995, 10), 1013 => to_unsigned(28, 10), 1014 => to_unsigned(331, 10), 1015 => to_unsigned(422, 10), 1016 => to_unsigned(73, 10), 1017 => to_unsigned(897, 10), 1018 => to_unsigned(399, 10), 1019 => to_unsigned(611, 10), 1020 => to_unsigned(788, 10), 1021 => to_unsigned(858, 10), 1022 => to_unsigned(635, 10), 1023 => to_unsigned(172, 10), 1024 => to_unsigned(396, 10), 1025 => to_unsigned(239, 10), 1026 => to_unsigned(617, 10), 1027 => to_unsigned(682, 10), 1028 => to_unsigned(79, 10), 1029 => to_unsigned(820, 10), 1030 => to_unsigned(1019, 10), 1031 => to_unsigned(709, 10), 1032 => to_unsigned(725, 10), 1033 => to_unsigned(796, 10), 1034 => to_unsigned(294, 10), 1035 => to_unsigned(391, 10), 1036 => to_unsigned(531, 10), 1037 => to_unsigned(390, 10), 1038 => to_unsigned(588, 10), 1039 => to_unsigned(137, 10), 1040 => to_unsigned(26, 10), 1041 => to_unsigned(148, 10), 1042 => to_unsigned(358, 10), 1043 => to_unsigned(548, 10), 1044 => to_unsigned(886, 10), 1045 => to_unsigned(159, 10), 1046 => to_unsigned(297, 10), 1047 => to_unsigned(212, 10), 1048 => to_unsigned(656, 10), 1049 => to_unsigned(416, 10), 1050 => to_unsigned(475, 10), 1051 => to_unsigned(460, 10), 1052 => to_unsigned(159, 10), 1053 => to_unsigned(47, 10), 1054 => to_unsigned(243, 10), 1055 => to_unsigned(614, 10), 1056 => to_unsigned(548, 10), 1057 => to_unsigned(753, 10), 1058 => to_unsigned(151, 10), 1059 => to_unsigned(914, 10), 1060 => to_unsigned(282, 10), 1061 => to_unsigned(307, 10), 1062 => to_unsigned(560, 10), 1063 => to_unsigned(511, 10), 1064 => to_unsigned(845, 10), 1065 => to_unsigned(117, 10), 1066 => to_unsigned(670, 10), 1067 => to_unsigned(119, 10), 1068 => to_unsigned(372, 10), 1069 => to_unsigned(79, 10), 1070 => to_unsigned(706, 10), 1071 => to_unsigned(843, 10), 1072 => to_unsigned(388, 10), 1073 => to_unsigned(967, 10), 1074 => to_unsigned(465, 10), 1075 => to_unsigned(979, 10), 1076 => to_unsigned(576, 10), 1077 => to_unsigned(156, 10), 1078 => to_unsigned(740, 10), 1079 => to_unsigned(439, 10), 1080 => to_unsigned(103, 10), 1081 => to_unsigned(318, 10), 1082 => to_unsigned(238, 10), 1083 => to_unsigned(698, 10), 1084 => to_unsigned(463, 10), 1085 => to_unsigned(226, 10), 1086 => to_unsigned(326, 10), 1087 => to_unsigned(557, 10), 1088 => to_unsigned(163, 10), 1089 => to_unsigned(565, 10), 1090 => to_unsigned(392, 10), 1091 => to_unsigned(205, 10), 1092 => to_unsigned(399, 10), 1093 => to_unsigned(719, 10), 1094 => to_unsigned(754, 10), 1095 => to_unsigned(236, 10), 1096 => to_unsigned(509, 10), 1097 => to_unsigned(731, 10), 1098 => to_unsigned(915, 10), 1099 => to_unsigned(448, 10), 1100 => to_unsigned(842, 10), 1101 => to_unsigned(266, 10), 1102 => to_unsigned(949, 10), 1103 => to_unsigned(494, 10), 1104 => to_unsigned(480, 10), 1105 => to_unsigned(900, 10), 1106 => to_unsigned(195, 10), 1107 => to_unsigned(680, 10), 1108 => to_unsigned(905, 10), 1109 => to_unsigned(311, 10), 1110 => to_unsigned(896, 10), 1111 => to_unsigned(803, 10), 1112 => to_unsigned(668, 10), 1113 => to_unsigned(350, 10), 1114 => to_unsigned(697, 10), 1115 => to_unsigned(81, 10), 1116 => to_unsigned(69, 10), 1117 => to_unsigned(737, 10), 1118 => to_unsigned(886, 10), 1119 => to_unsigned(235, 10), 1120 => to_unsigned(813, 10), 1121 => to_unsigned(261, 10), 1122 => to_unsigned(792, 10), 1123 => to_unsigned(751, 10), 1124 => to_unsigned(469, 10), 1125 => to_unsigned(525, 10), 1126 => to_unsigned(511, 10), 1127 => to_unsigned(663, 10), 1128 => to_unsigned(930, 10), 1129 => to_unsigned(349, 10), 1130 => to_unsigned(971, 10), 1131 => to_unsigned(203, 10), 1132 => to_unsigned(981, 10), 1133 => to_unsigned(475, 10), 1134 => to_unsigned(954, 10), 1135 => to_unsigned(510, 10), 1136 => to_unsigned(685, 10), 1137 => to_unsigned(235, 10), 1138 => to_unsigned(194, 10), 1139 => to_unsigned(425, 10), 1140 => to_unsigned(519, 10), 1141 => to_unsigned(655, 10), 1142 => to_unsigned(384, 10), 1143 => to_unsigned(478, 10), 1144 => to_unsigned(431, 10), 1145 => to_unsigned(123, 10), 1146 => to_unsigned(42, 10), 1147 => to_unsigned(742, 10), 1148 => to_unsigned(241, 10), 1149 => to_unsigned(332, 10), 1150 => to_unsigned(464, 10), 1151 => to_unsigned(157, 10), 1152 => to_unsigned(855, 10), 1153 => to_unsigned(839, 10), 1154 => to_unsigned(622, 10), 1155 => to_unsigned(836, 10), 1156 => to_unsigned(543, 10), 1157 => to_unsigned(160, 10), 1158 => to_unsigned(899, 10), 1159 => to_unsigned(101, 10), 1160 => to_unsigned(398, 10), 1161 => to_unsigned(322, 10), 1162 => to_unsigned(16, 10), 1163 => to_unsigned(159, 10), 1164 => to_unsigned(126, 10), 1165 => to_unsigned(115, 10), 1166 => to_unsigned(23, 10), 1167 => to_unsigned(729, 10), 1168 => to_unsigned(283, 10), 1169 => to_unsigned(733, 10), 1170 => to_unsigned(279, 10), 1171 => to_unsigned(844, 10), 1172 => to_unsigned(741, 10), 1173 => to_unsigned(808, 10), 1174 => to_unsigned(999, 10), 1175 => to_unsigned(434, 10), 1176 => to_unsigned(268, 10), 1177 => to_unsigned(313, 10), 1178 => to_unsigned(675, 10), 1179 => to_unsigned(704, 10), 1180 => to_unsigned(350, 10), 1181 => to_unsigned(529, 10), 1182 => to_unsigned(1010, 10), 1183 => to_unsigned(55, 10), 1184 => to_unsigned(284, 10), 1185 => to_unsigned(176, 10), 1186 => to_unsigned(841, 10), 1187 => to_unsigned(130, 10), 1188 => to_unsigned(803, 10), 1189 => to_unsigned(778, 10), 1190 => to_unsigned(924, 10), 1191 => to_unsigned(553, 10), 1192 => to_unsigned(386, 10), 1193 => to_unsigned(72, 10), 1194 => to_unsigned(108, 10), 1195 => to_unsigned(976, 10), 1196 => to_unsigned(26, 10), 1197 => to_unsigned(210, 10), 1198 => to_unsigned(996, 10), 1199 => to_unsigned(660, 10), 1200 => to_unsigned(443, 10), 1201 => to_unsigned(490, 10), 1202 => to_unsigned(461, 10), 1203 => to_unsigned(13, 10), 1204 => to_unsigned(14, 10), 1205 => to_unsigned(1018, 10), 1206 => to_unsigned(480, 10), 1207 => to_unsigned(949, 10), 1208 => to_unsigned(139, 10), 1209 => to_unsigned(367, 10), 1210 => to_unsigned(816, 10), 1211 => to_unsigned(186, 10), 1212 => to_unsigned(264, 10), 1213 => to_unsigned(497, 10), 1214 => to_unsigned(492, 10), 1215 => to_unsigned(40, 10), 1216 => to_unsigned(48, 10), 1217 => to_unsigned(162, 10), 1218 => to_unsigned(165, 10), 1219 => to_unsigned(867, 10), 1220 => to_unsigned(621, 10), 1221 => to_unsigned(808, 10), 1222 => to_unsigned(633, 10), 1223 => to_unsigned(522, 10), 1224 => to_unsigned(47, 10), 1225 => to_unsigned(891, 10), 1226 => to_unsigned(535, 10), 1227 => to_unsigned(56, 10), 1228 => to_unsigned(678, 10), 1229 => to_unsigned(132, 10), 1230 => to_unsigned(948, 10), 1231 => to_unsigned(830, 10), 1232 => to_unsigned(1020, 10), 1233 => to_unsigned(1015, 10), 1234 => to_unsigned(687, 10), 1235 => to_unsigned(794, 10), 1236 => to_unsigned(711, 10), 1237 => to_unsigned(244, 10), 1238 => to_unsigned(243, 10), 1239 => to_unsigned(90, 10), 1240 => to_unsigned(25, 10), 1241 => to_unsigned(297, 10), 1242 => to_unsigned(20, 10), 1243 => to_unsigned(1021, 10), 1244 => to_unsigned(159, 10), 1245 => to_unsigned(366, 10), 1246 => to_unsigned(759, 10), 1247 => to_unsigned(182, 10), 1248 => to_unsigned(130, 10), 1249 => to_unsigned(446, 10), 1250 => to_unsigned(823, 10), 1251 => to_unsigned(644, 10), 1252 => to_unsigned(990, 10), 1253 => to_unsigned(540, 10), 1254 => to_unsigned(269, 10), 1255 => to_unsigned(25, 10), 1256 => to_unsigned(861, 10), 1257 => to_unsigned(113, 10), 1258 => to_unsigned(82, 10), 1259 => to_unsigned(534, 10), 1260 => to_unsigned(900, 10), 1261 => to_unsigned(434, 10), 1262 => to_unsigned(375, 10), 1263 => to_unsigned(891, 10), 1264 => to_unsigned(499, 10), 1265 => to_unsigned(109, 10), 1266 => to_unsigned(352, 10), 1267 => to_unsigned(551, 10), 1268 => to_unsigned(657, 10), 1269 => to_unsigned(578, 10), 1270 => to_unsigned(988, 10), 1271 => to_unsigned(312, 10), 1272 => to_unsigned(667, 10), 1273 => to_unsigned(78, 10), 1274 => to_unsigned(340, 10), 1275 => to_unsigned(160, 10), 1276 => to_unsigned(631, 10), 1277 => to_unsigned(152, 10), 1278 => to_unsigned(331, 10), 1279 => to_unsigned(78, 10), 1280 => to_unsigned(14, 10), 1281 => to_unsigned(1005, 10), 1282 => to_unsigned(748, 10), 1283 => to_unsigned(932, 10), 1284 => to_unsigned(392, 10), 1285 => to_unsigned(813, 10), 1286 => to_unsigned(501, 10), 1287 => to_unsigned(217, 10), 1288 => to_unsigned(881, 10), 1289 => to_unsigned(433, 10), 1290 => to_unsigned(87, 10), 1291 => to_unsigned(936, 10), 1292 => to_unsigned(265, 10), 1293 => to_unsigned(819, 10), 1294 => to_unsigned(616, 10), 1295 => to_unsigned(941, 10), 1296 => to_unsigned(473, 10), 1297 => to_unsigned(62, 10), 1298 => to_unsigned(10, 10), 1299 => to_unsigned(500, 10), 1300 => to_unsigned(79, 10), 1301 => to_unsigned(1000, 10), 1302 => to_unsigned(423, 10), 1303 => to_unsigned(934, 10), 1304 => to_unsigned(380, 10), 1305 => to_unsigned(772, 10), 1306 => to_unsigned(767, 10), 1307 => to_unsigned(673, 10), 1308 => to_unsigned(202, 10), 1309 => to_unsigned(889, 10), 1310 => to_unsigned(565, 10), 1311 => to_unsigned(162, 10), 1312 => to_unsigned(322, 10), 1313 => to_unsigned(175, 10), 1314 => to_unsigned(829, 10), 1315 => to_unsigned(452, 10), 1316 => to_unsigned(484, 10), 1317 => to_unsigned(418, 10), 1318 => to_unsigned(1013, 10), 1319 => to_unsigned(34, 10), 1320 => to_unsigned(274, 10), 1321 => to_unsigned(364, 10), 1322 => to_unsigned(517, 10), 1323 => to_unsigned(1013, 10), 1324 => to_unsigned(283, 10), 1325 => to_unsigned(147, 10), 1326 => to_unsigned(117, 10), 1327 => to_unsigned(80, 10), 1328 => to_unsigned(611, 10), 1329 => to_unsigned(809, 10), 1330 => to_unsigned(422, 10), 1331 => to_unsigned(988, 10), 1332 => to_unsigned(651, 10), 1333 => to_unsigned(378, 10), 1334 => to_unsigned(239, 10), 1335 => to_unsigned(1018, 10), 1336 => to_unsigned(313, 10), 1337 => to_unsigned(448, 10), 1338 => to_unsigned(402, 10), 1339 => to_unsigned(293, 10), 1340 => to_unsigned(550, 10), 1341 => to_unsigned(782, 10), 1342 => to_unsigned(715, 10), 1343 => to_unsigned(933, 10), 1344 => to_unsigned(778, 10), 1345 => to_unsigned(727, 10), 1346 => to_unsigned(135, 10), 1347 => to_unsigned(215, 10), 1348 => to_unsigned(88, 10), 1349 => to_unsigned(145, 10), 1350 => to_unsigned(784, 10), 1351 => to_unsigned(120, 10), 1352 => to_unsigned(796, 10), 1353 => to_unsigned(370, 10), 1354 => to_unsigned(439, 10), 1355 => to_unsigned(21, 10), 1356 => to_unsigned(722, 10), 1357 => to_unsigned(523, 10), 1358 => to_unsigned(216, 10), 1359 => to_unsigned(89, 10), 1360 => to_unsigned(346, 10), 1361 => to_unsigned(230, 10), 1362 => to_unsigned(1006, 10), 1363 => to_unsigned(15, 10), 1364 => to_unsigned(890, 10), 1365 => to_unsigned(503, 10), 1366 => to_unsigned(805, 10), 1367 => to_unsigned(609, 10), 1368 => to_unsigned(21, 10), 1369 => to_unsigned(77, 10), 1370 => to_unsigned(606, 10), 1371 => to_unsigned(84, 10), 1372 => to_unsigned(990, 10), 1373 => to_unsigned(667, 10), 1374 => to_unsigned(738, 10), 1375 => to_unsigned(605, 10), 1376 => to_unsigned(514, 10), 1377 => to_unsigned(395, 10), 1378 => to_unsigned(987, 10), 1379 => to_unsigned(290, 10), 1380 => to_unsigned(886, 10), 1381 => to_unsigned(891, 10), 1382 => to_unsigned(1019, 10), 1383 => to_unsigned(321, 10), 1384 => to_unsigned(243, 10), 1385 => to_unsigned(73, 10), 1386 => to_unsigned(86, 10), 1387 => to_unsigned(407, 10), 1388 => to_unsigned(344, 10), 1389 => to_unsigned(323, 10), 1390 => to_unsigned(189, 10), 1391 => to_unsigned(609, 10), 1392 => to_unsigned(856, 10), 1393 => to_unsigned(895, 10), 1394 => to_unsigned(155, 10), 1395 => to_unsigned(371, 10), 1396 => to_unsigned(460, 10), 1397 => to_unsigned(1022, 10), 1398 => to_unsigned(103, 10), 1399 => to_unsigned(90, 10), 1400 => to_unsigned(101, 10), 1401 => to_unsigned(628, 10), 1402 => to_unsigned(159, 10), 1403 => to_unsigned(806, 10), 1404 => to_unsigned(571, 10), 1405 => to_unsigned(156, 10), 1406 => to_unsigned(420, 10), 1407 => to_unsigned(979, 10), 1408 => to_unsigned(453, 10), 1409 => to_unsigned(943, 10), 1410 => to_unsigned(647, 10), 1411 => to_unsigned(783, 10), 1412 => to_unsigned(546, 10), 1413 => to_unsigned(141, 10), 1414 => to_unsigned(88, 10), 1415 => to_unsigned(693, 10), 1416 => to_unsigned(759, 10), 1417 => to_unsigned(367, 10), 1418 => to_unsigned(171, 10), 1419 => to_unsigned(467, 10), 1420 => to_unsigned(57, 10), 1421 => to_unsigned(432, 10), 1422 => to_unsigned(395, 10), 1423 => to_unsigned(738, 10), 1424 => to_unsigned(88, 10), 1425 => to_unsigned(661, 10), 1426 => to_unsigned(881, 10), 1427 => to_unsigned(470, 10), 1428 => to_unsigned(952, 10), 1429 => to_unsigned(481, 10), 1430 => to_unsigned(755, 10), 1431 => to_unsigned(39, 10), 1432 => to_unsigned(683, 10), 1433 => to_unsigned(864, 10), 1434 => to_unsigned(402, 10), 1435 => to_unsigned(124, 10), 1436 => to_unsigned(144, 10), 1437 => to_unsigned(5, 10), 1438 => to_unsigned(415, 10), 1439 => to_unsigned(20, 10), 1440 => to_unsigned(283, 10), 1441 => to_unsigned(1002, 10), 1442 => to_unsigned(213, 10), 1443 => to_unsigned(710, 10), 1444 => to_unsigned(791, 10), 1445 => to_unsigned(752, 10), 1446 => to_unsigned(743, 10), 1447 => to_unsigned(695, 10), 1448 => to_unsigned(543, 10), 1449 => to_unsigned(52, 10), 1450 => to_unsigned(637, 10), 1451 => to_unsigned(904, 10), 1452 => to_unsigned(824, 10), 1453 => to_unsigned(170, 10), 1454 => to_unsigned(756, 10), 1455 => to_unsigned(1023, 10), 1456 => to_unsigned(739, 10), 1457 => to_unsigned(731, 10), 1458 => to_unsigned(739, 10), 1459 => to_unsigned(769, 10), 1460 => to_unsigned(633, 10), 1461 => to_unsigned(294, 10), 1462 => to_unsigned(482, 10), 1463 => to_unsigned(476, 10), 1464 => to_unsigned(484, 10), 1465 => to_unsigned(662, 10), 1466 => to_unsigned(905, 10), 1467 => to_unsigned(159, 10), 1468 => to_unsigned(878, 10), 1469 => to_unsigned(889, 10), 1470 => to_unsigned(89, 10), 1471 => to_unsigned(258, 10), 1472 => to_unsigned(133, 10), 1473 => to_unsigned(735, 10), 1474 => to_unsigned(157, 10), 1475 => to_unsigned(872, 10), 1476 => to_unsigned(472, 10), 1477 => to_unsigned(501, 10), 1478 => to_unsigned(944, 10), 1479 => to_unsigned(990, 10), 1480 => to_unsigned(340, 10), 1481 => to_unsigned(205, 10), 1482 => to_unsigned(440, 10), 1483 => to_unsigned(482, 10), 1484 => to_unsigned(665, 10), 1485 => to_unsigned(44, 10), 1486 => to_unsigned(901, 10), 1487 => to_unsigned(736, 10), 1488 => to_unsigned(617, 10), 1489 => to_unsigned(388, 10), 1490 => to_unsigned(803, 10), 1491 => to_unsigned(87, 10), 1492 => to_unsigned(490, 10), 1493 => to_unsigned(890, 10), 1494 => to_unsigned(2, 10), 1495 => to_unsigned(338, 10), 1496 => to_unsigned(778, 10), 1497 => to_unsigned(688, 10), 1498 => to_unsigned(816, 10), 1499 => to_unsigned(539, 10), 1500 => to_unsigned(28, 10), 1501 => to_unsigned(120, 10), 1502 => to_unsigned(470, 10), 1503 => to_unsigned(498, 10), 1504 => to_unsigned(613, 10), 1505 => to_unsigned(225, 10), 1506 => to_unsigned(631, 10), 1507 => to_unsigned(649, 10), 1508 => to_unsigned(878, 10), 1509 => to_unsigned(788, 10), 1510 => to_unsigned(1003, 10), 1511 => to_unsigned(411, 10), 1512 => to_unsigned(1008, 10), 1513 => to_unsigned(483, 10), 1514 => to_unsigned(5, 10), 1515 => to_unsigned(219, 10), 1516 => to_unsigned(438, 10), 1517 => to_unsigned(714, 10), 1518 => to_unsigned(229, 10), 1519 => to_unsigned(933, 10), 1520 => to_unsigned(929, 10), 1521 => to_unsigned(496, 10), 1522 => to_unsigned(791, 10), 1523 => to_unsigned(499, 10), 1524 => to_unsigned(355, 10), 1525 => to_unsigned(49, 10), 1526 => to_unsigned(356, 10), 1527 => to_unsigned(62, 10), 1528 => to_unsigned(456, 10), 1529 => to_unsigned(373, 10), 1530 => to_unsigned(523, 10), 1531 => to_unsigned(248, 10), 1532 => to_unsigned(502, 10), 1533 => to_unsigned(333, 10), 1534 => to_unsigned(759, 10), 1535 => to_unsigned(13, 10), 1536 => to_unsigned(750, 10), 1537 => to_unsigned(917, 10), 1538 => to_unsigned(223, 10), 1539 => to_unsigned(400, 10), 1540 => to_unsigned(820, 10), 1541 => to_unsigned(382, 10), 1542 => to_unsigned(835, 10), 1543 => to_unsigned(301, 10), 1544 => to_unsigned(600, 10), 1545 => to_unsigned(491, 10), 1546 => to_unsigned(293, 10), 1547 => to_unsigned(630, 10), 1548 => to_unsigned(341, 10), 1549 => to_unsigned(725, 10), 1550 => to_unsigned(779, 10), 1551 => to_unsigned(554, 10), 1552 => to_unsigned(252, 10), 1553 => to_unsigned(815, 10), 1554 => to_unsigned(688, 10), 1555 => to_unsigned(13, 10), 1556 => to_unsigned(160, 10), 1557 => to_unsigned(711, 10), 1558 => to_unsigned(203, 10), 1559 => to_unsigned(231, 10), 1560 => to_unsigned(872, 10), 1561 => to_unsigned(962, 10), 1562 => to_unsigned(686, 10), 1563 => to_unsigned(74, 10), 1564 => to_unsigned(945, 10), 1565 => to_unsigned(599, 10), 1566 => to_unsigned(351, 10), 1567 => to_unsigned(550, 10), 1568 => to_unsigned(672, 10), 1569 => to_unsigned(47, 10), 1570 => to_unsigned(94, 10), 1571 => to_unsigned(448, 10), 1572 => to_unsigned(886, 10), 1573 => to_unsigned(821, 10), 1574 => to_unsigned(716, 10), 1575 => to_unsigned(917, 10), 1576 => to_unsigned(651, 10), 1577 => to_unsigned(284, 10), 1578 => to_unsigned(330, 10), 1579 => to_unsigned(279, 10), 1580 => to_unsigned(13, 10), 1581 => to_unsigned(256, 10), 1582 => to_unsigned(525, 10), 1583 => to_unsigned(656, 10), 1584 => to_unsigned(540, 10), 1585 => to_unsigned(533, 10), 1586 => to_unsigned(844, 10), 1587 => to_unsigned(421, 10), 1588 => to_unsigned(81, 10), 1589 => to_unsigned(229, 10), 1590 => to_unsigned(545, 10), 1591 => to_unsigned(302, 10), 1592 => to_unsigned(709, 10), 1593 => to_unsigned(73, 10), 1594 => to_unsigned(855, 10), 1595 => to_unsigned(468, 10), 1596 => to_unsigned(347, 10), 1597 => to_unsigned(93, 10), 1598 => to_unsigned(599, 10), 1599 => to_unsigned(412, 10), 1600 => to_unsigned(1021, 10), 1601 => to_unsigned(290, 10), 1602 => to_unsigned(0, 10), 1603 => to_unsigned(787, 10), 1604 => to_unsigned(552, 10), 1605 => to_unsigned(923, 10), 1606 => to_unsigned(555, 10), 1607 => to_unsigned(866, 10), 1608 => to_unsigned(941, 10), 1609 => to_unsigned(206, 10), 1610 => to_unsigned(666, 10), 1611 => to_unsigned(626, 10), 1612 => to_unsigned(912, 10), 1613 => to_unsigned(538, 10), 1614 => to_unsigned(643, 10), 1615 => to_unsigned(544, 10), 1616 => to_unsigned(199, 10), 1617 => to_unsigned(547, 10), 1618 => to_unsigned(695, 10), 1619 => to_unsigned(225, 10), 1620 => to_unsigned(629, 10), 1621 => to_unsigned(373, 10), 1622 => to_unsigned(471, 10), 1623 => to_unsigned(688, 10), 1624 => to_unsigned(99, 10), 1625 => to_unsigned(451, 10), 1626 => to_unsigned(422, 10), 1627 => to_unsigned(704, 10), 1628 => to_unsigned(433, 10), 1629 => to_unsigned(439, 10), 1630 => to_unsigned(614, 10), 1631 => to_unsigned(40, 10), 1632 => to_unsigned(634, 10), 1633 => to_unsigned(711, 10), 1634 => to_unsigned(922, 10), 1635 => to_unsigned(914, 10), 1636 => to_unsigned(652, 10), 1637 => to_unsigned(6, 10), 1638 => to_unsigned(225, 10), 1639 => to_unsigned(648, 10), 1640 => to_unsigned(36, 10), 1641 => to_unsigned(985, 10), 1642 => to_unsigned(517, 10), 1643 => to_unsigned(987, 10), 1644 => to_unsigned(280, 10), 1645 => to_unsigned(338, 10), 1646 => to_unsigned(825, 10), 1647 => to_unsigned(763, 10), 1648 => to_unsigned(287, 10), 1649 => to_unsigned(97, 10), 1650 => to_unsigned(691, 10), 1651 => to_unsigned(737, 10), 1652 => to_unsigned(666, 10), 1653 => to_unsigned(351, 10), 1654 => to_unsigned(14, 10), 1655 => to_unsigned(12, 10), 1656 => to_unsigned(382, 10), 1657 => to_unsigned(803, 10), 1658 => to_unsigned(792, 10), 1659 => to_unsigned(584, 10), 1660 => to_unsigned(119, 10), 1661 => to_unsigned(393, 10), 1662 => to_unsigned(180, 10), 1663 => to_unsigned(615, 10), 1664 => to_unsigned(331, 10), 1665 => to_unsigned(972, 10), 1666 => to_unsigned(913, 10), 1667 => to_unsigned(867, 10), 1668 => to_unsigned(864, 10), 1669 => to_unsigned(896, 10), 1670 => to_unsigned(750, 10), 1671 => to_unsigned(267, 10), 1672 => to_unsigned(723, 10), 1673 => to_unsigned(699, 10), 1674 => to_unsigned(600, 10), 1675 => to_unsigned(907, 10), 1676 => to_unsigned(766, 10), 1677 => to_unsigned(883, 10), 1678 => to_unsigned(860, 10), 1679 => to_unsigned(849, 10), 1680 => to_unsigned(644, 10), 1681 => to_unsigned(697, 10), 1682 => to_unsigned(278, 10), 1683 => to_unsigned(598, 10), 1684 => to_unsigned(182, 10), 1685 => to_unsigned(1, 10), 1686 => to_unsigned(749, 10), 1687 => to_unsigned(129, 10), 1688 => to_unsigned(136, 10), 1689 => to_unsigned(279, 10), 1690 => to_unsigned(879, 10), 1691 => to_unsigned(848, 10), 1692 => to_unsigned(358, 10), 1693 => to_unsigned(726, 10), 1694 => to_unsigned(971, 10), 1695 => to_unsigned(447, 10), 1696 => to_unsigned(236, 10), 1697 => to_unsigned(92, 10), 1698 => to_unsigned(931, 10), 1699 => to_unsigned(460, 10), 1700 => to_unsigned(323, 10), 1701 => to_unsigned(1002, 10), 1702 => to_unsigned(460, 10), 1703 => to_unsigned(952, 10), 1704 => to_unsigned(258, 10), 1705 => to_unsigned(11, 10), 1706 => to_unsigned(200, 10), 1707 => to_unsigned(636, 10), 1708 => to_unsigned(961, 10), 1709 => to_unsigned(147, 10), 1710 => to_unsigned(996, 10), 1711 => to_unsigned(116, 10), 1712 => to_unsigned(926, 10), 1713 => to_unsigned(851, 10), 1714 => to_unsigned(147, 10), 1715 => to_unsigned(867, 10), 1716 => to_unsigned(884, 10), 1717 => to_unsigned(455, 10), 1718 => to_unsigned(394, 10), 1719 => to_unsigned(493, 10), 1720 => to_unsigned(377, 10), 1721 => to_unsigned(28, 10), 1722 => to_unsigned(803, 10), 1723 => to_unsigned(690, 10), 1724 => to_unsigned(879, 10), 1725 => to_unsigned(689, 10), 1726 => to_unsigned(946, 10), 1727 => to_unsigned(131, 10), 1728 => to_unsigned(329, 10), 1729 => to_unsigned(618, 10), 1730 => to_unsigned(82, 10), 1731 => to_unsigned(639, 10), 1732 => to_unsigned(438, 10), 1733 => to_unsigned(69, 10), 1734 => to_unsigned(922, 10), 1735 => to_unsigned(189, 10), 1736 => to_unsigned(951, 10), 1737 => to_unsigned(847, 10), 1738 => to_unsigned(893, 10), 1739 => to_unsigned(662, 10), 1740 => to_unsigned(375, 10), 1741 => to_unsigned(269, 10), 1742 => to_unsigned(254, 10), 1743 => to_unsigned(721, 10), 1744 => to_unsigned(43, 10), 1745 => to_unsigned(825, 10), 1746 => to_unsigned(930, 10), 1747 => to_unsigned(782, 10), 1748 => to_unsigned(522, 10), 1749 => to_unsigned(835, 10), 1750 => to_unsigned(328, 10), 1751 => to_unsigned(987, 10), 1752 => to_unsigned(65, 10), 1753 => to_unsigned(871, 10), 1754 => to_unsigned(690, 10), 1755 => to_unsigned(492, 10), 1756 => to_unsigned(658, 10), 1757 => to_unsigned(695, 10), 1758 => to_unsigned(1022, 10), 1759 => to_unsigned(328, 10), 1760 => to_unsigned(0, 10), 1761 => to_unsigned(243, 10), 1762 => to_unsigned(332, 10), 1763 => to_unsigned(381, 10), 1764 => to_unsigned(127, 10), 1765 => to_unsigned(425, 10), 1766 => to_unsigned(715, 10), 1767 => to_unsigned(138, 10), 1768 => to_unsigned(44, 10), 1769 => to_unsigned(618, 10), 1770 => to_unsigned(6, 10), 1771 => to_unsigned(214, 10), 1772 => to_unsigned(1004, 10), 1773 => to_unsigned(455, 10), 1774 => to_unsigned(524, 10), 1775 => to_unsigned(852, 10), 1776 => to_unsigned(553, 10), 1777 => to_unsigned(605, 10), 1778 => to_unsigned(356, 10), 1779 => to_unsigned(387, 10), 1780 => to_unsigned(376, 10), 1781 => to_unsigned(876, 10), 1782 => to_unsigned(775, 10), 1783 => to_unsigned(461, 10), 1784 => to_unsigned(313, 10), 1785 => to_unsigned(658, 10), 1786 => to_unsigned(444, 10), 1787 => to_unsigned(600, 10), 1788 => to_unsigned(1017, 10), 1789 => to_unsigned(225, 10), 1790 => to_unsigned(98, 10), 1791 => to_unsigned(876, 10), 1792 => to_unsigned(469, 10), 1793 => to_unsigned(35, 10), 1794 => to_unsigned(604, 10), 1795 => to_unsigned(241, 10), 1796 => to_unsigned(383, 10), 1797 => to_unsigned(614, 10), 1798 => to_unsigned(236, 10), 1799 => to_unsigned(795, 10), 1800 => to_unsigned(606, 10), 1801 => to_unsigned(731, 10), 1802 => to_unsigned(833, 10), 1803 => to_unsigned(8, 10), 1804 => to_unsigned(885, 10), 1805 => to_unsigned(857, 10), 1806 => to_unsigned(285, 10), 1807 => to_unsigned(655, 10), 1808 => to_unsigned(259, 10), 1809 => to_unsigned(435, 10), 1810 => to_unsigned(663, 10), 1811 => to_unsigned(863, 10), 1812 => to_unsigned(886, 10), 1813 => to_unsigned(228, 10), 1814 => to_unsigned(21, 10), 1815 => to_unsigned(341, 10), 1816 => to_unsigned(962, 10), 1817 => to_unsigned(371, 10), 1818 => to_unsigned(991, 10), 1819 => to_unsigned(200, 10), 1820 => to_unsigned(709, 10), 1821 => to_unsigned(441, 10), 1822 => to_unsigned(563, 10), 1823 => to_unsigned(524, 10), 1824 => to_unsigned(612, 10), 1825 => to_unsigned(138, 10), 1826 => to_unsigned(185, 10), 1827 => to_unsigned(870, 10), 1828 => to_unsigned(187, 10), 1829 => to_unsigned(306, 10), 1830 => to_unsigned(232, 10), 1831 => to_unsigned(203, 10), 1832 => to_unsigned(42, 10), 1833 => to_unsigned(767, 10), 1834 => to_unsigned(413, 10), 1835 => to_unsigned(357, 10), 1836 => to_unsigned(565, 10), 1837 => to_unsigned(424, 10), 1838 => to_unsigned(428, 10), 1839 => to_unsigned(329, 10), 1840 => to_unsigned(425, 10), 1841 => to_unsigned(88, 10), 1842 => to_unsigned(811, 10), 1843 => to_unsigned(935, 10), 1844 => to_unsigned(481, 10), 1845 => to_unsigned(969, 10), 1846 => to_unsigned(518, 10), 1847 => to_unsigned(600, 10), 1848 => to_unsigned(663, 10), 1849 => to_unsigned(808, 10), 1850 => to_unsigned(517, 10), 1851 => to_unsigned(654, 10), 1852 => to_unsigned(1020, 10), 1853 => to_unsigned(983, 10), 1854 => to_unsigned(656, 10), 1855 => to_unsigned(168, 10), 1856 => to_unsigned(282, 10), 1857 => to_unsigned(526, 10), 1858 => to_unsigned(459, 10), 1859 => to_unsigned(314, 10), 1860 => to_unsigned(719, 10), 1861 => to_unsigned(744, 10), 1862 => to_unsigned(271, 10), 1863 => to_unsigned(700, 10), 1864 => to_unsigned(659, 10), 1865 => to_unsigned(122, 10), 1866 => to_unsigned(338, 10), 1867 => to_unsigned(190, 10), 1868 => to_unsigned(319, 10), 1869 => to_unsigned(379, 10), 1870 => to_unsigned(591, 10), 1871 => to_unsigned(645, 10), 1872 => to_unsigned(327, 10), 1873 => to_unsigned(583, 10), 1874 => to_unsigned(918, 10), 1875 => to_unsigned(560, 10), 1876 => to_unsigned(851, 10), 1877 => to_unsigned(782, 10), 1878 => to_unsigned(770, 10), 1879 => to_unsigned(1017, 10), 1880 => to_unsigned(875, 10), 1881 => to_unsigned(975, 10), 1882 => to_unsigned(916, 10), 1883 => to_unsigned(394, 10), 1884 => to_unsigned(341, 10), 1885 => to_unsigned(362, 10), 1886 => to_unsigned(297, 10), 1887 => to_unsigned(561, 10), 1888 => to_unsigned(953, 10), 1889 => to_unsigned(945, 10), 1890 => to_unsigned(496, 10), 1891 => to_unsigned(413, 10), 1892 => to_unsigned(619, 10), 1893 => to_unsigned(324, 10), 1894 => to_unsigned(676, 10), 1895 => to_unsigned(714, 10), 1896 => to_unsigned(320, 10), 1897 => to_unsigned(146, 10), 1898 => to_unsigned(44, 10), 1899 => to_unsigned(387, 10), 1900 => to_unsigned(560, 10), 1901 => to_unsigned(856, 10), 1902 => to_unsigned(156, 10), 1903 => to_unsigned(802, 10), 1904 => to_unsigned(747, 10), 1905 => to_unsigned(840, 10), 1906 => to_unsigned(122, 10), 1907 => to_unsigned(312, 10), 1908 => to_unsigned(805, 10), 1909 => to_unsigned(234, 10), 1910 => to_unsigned(735, 10), 1911 => to_unsigned(361, 10), 1912 => to_unsigned(882, 10), 1913 => to_unsigned(908, 10), 1914 => to_unsigned(299, 10), 1915 => to_unsigned(294, 10), 1916 => to_unsigned(688, 10), 1917 => to_unsigned(474, 10), 1918 => to_unsigned(772, 10), 1919 => to_unsigned(934, 10), 1920 => to_unsigned(207, 10), 1921 => to_unsigned(667, 10), 1922 => to_unsigned(245, 10), 1923 => to_unsigned(10, 10), 1924 => to_unsigned(106, 10), 1925 => to_unsigned(775, 10), 1926 => to_unsigned(694, 10), 1927 => to_unsigned(728, 10), 1928 => to_unsigned(929, 10), 1929 => to_unsigned(736, 10), 1930 => to_unsigned(313, 10), 1931 => to_unsigned(446, 10), 1932 => to_unsigned(763, 10), 1933 => to_unsigned(216, 10), 1934 => to_unsigned(212, 10), 1935 => to_unsigned(734, 10), 1936 => to_unsigned(260, 10), 1937 => to_unsigned(53, 10), 1938 => to_unsigned(908, 10), 1939 => to_unsigned(158, 10), 1940 => to_unsigned(302, 10), 1941 => to_unsigned(20, 10), 1942 => to_unsigned(481, 10), 1943 => to_unsigned(570, 10), 1944 => to_unsigned(563, 10), 1945 => to_unsigned(901, 10), 1946 => to_unsigned(60, 10), 1947 => to_unsigned(339, 10), 1948 => to_unsigned(903, 10), 1949 => to_unsigned(430, 10), 1950 => to_unsigned(472, 10), 1951 => to_unsigned(393, 10), 1952 => to_unsigned(49, 10), 1953 => to_unsigned(785, 10), 1954 => to_unsigned(866, 10), 1955 => to_unsigned(910, 10), 1956 => to_unsigned(194, 10), 1957 => to_unsigned(103, 10), 1958 => to_unsigned(393, 10), 1959 => to_unsigned(442, 10), 1960 => to_unsigned(411, 10), 1961 => to_unsigned(971, 10), 1962 => to_unsigned(59, 10), 1963 => to_unsigned(107, 10), 1964 => to_unsigned(559, 10), 1965 => to_unsigned(501, 10), 1966 => to_unsigned(815, 10), 1967 => to_unsigned(726, 10), 1968 => to_unsigned(416, 10), 1969 => to_unsigned(360, 10), 1970 => to_unsigned(489, 10), 1971 => to_unsigned(309, 10), 1972 => to_unsigned(388, 10), 1973 => to_unsigned(541, 10), 1974 => to_unsigned(165, 10), 1975 => to_unsigned(42, 10), 1976 => to_unsigned(226, 10), 1977 => to_unsigned(239, 10), 1978 => to_unsigned(102, 10), 1979 => to_unsigned(789, 10), 1980 => to_unsigned(662, 10), 1981 => to_unsigned(822, 10), 1982 => to_unsigned(318, 10), 1983 => to_unsigned(401, 10), 1984 => to_unsigned(370, 10), 1985 => to_unsigned(3, 10), 1986 => to_unsigned(786, 10), 1987 => to_unsigned(965, 10), 1988 => to_unsigned(41, 10), 1989 => to_unsigned(546, 10), 1990 => to_unsigned(649, 10), 1991 => to_unsigned(114, 10), 1992 => to_unsigned(371, 10), 1993 => to_unsigned(860, 10), 1994 => to_unsigned(800, 10), 1995 => to_unsigned(541, 10), 1996 => to_unsigned(224, 10), 1997 => to_unsigned(351, 10), 1998 => to_unsigned(251, 10), 1999 => to_unsigned(330, 10), 2000 => to_unsigned(137, 10), 2001 => to_unsigned(405, 10), 2002 => to_unsigned(317, 10), 2003 => to_unsigned(570, 10), 2004 => to_unsigned(695, 10), 2005 => to_unsigned(99, 10), 2006 => to_unsigned(889, 10), 2007 => to_unsigned(254, 10), 2008 => to_unsigned(860, 10), 2009 => to_unsigned(905, 10), 2010 => to_unsigned(432, 10), 2011 => to_unsigned(298, 10), 2012 => to_unsigned(348, 10), 2013 => to_unsigned(581, 10), 2014 => to_unsigned(836, 10), 2015 => to_unsigned(529, 10), 2016 => to_unsigned(560, 10), 2017 => to_unsigned(240, 10), 2018 => to_unsigned(192, 10), 2019 => to_unsigned(308, 10), 2020 => to_unsigned(889, 10), 2021 => to_unsigned(772, 10), 2022 => to_unsigned(176, 10), 2023 => to_unsigned(895, 10), 2024 => to_unsigned(904, 10), 2025 => to_unsigned(231, 10), 2026 => to_unsigned(945, 10), 2027 => to_unsigned(856, 10), 2028 => to_unsigned(28, 10), 2029 => to_unsigned(57, 10), 2030 => to_unsigned(556, 10), 2031 => to_unsigned(731, 10), 2032 => to_unsigned(875, 10), 2033 => to_unsigned(678, 10), 2034 => to_unsigned(68, 10), 2035 => to_unsigned(602, 10), 2036 => to_unsigned(152, 10), 2037 => to_unsigned(75, 10), 2038 => to_unsigned(300, 10), 2039 => to_unsigned(281, 10), 2040 => to_unsigned(950, 10), 2041 => to_unsigned(52, 10), 2042 => to_unsigned(215, 10), 2043 => to_unsigned(347, 10), 2044 => to_unsigned(304, 10), 2045 => to_unsigned(831, 10), 2046 => to_unsigned(276, 10), 2047 => to_unsigned(531, 10)),
            6 => (0 => to_unsigned(828, 10), 1 => to_unsigned(884, 10), 2 => to_unsigned(651, 10), 3 => to_unsigned(218, 10), 4 => to_unsigned(297, 10), 5 => to_unsigned(41, 10), 6 => to_unsigned(774, 10), 7 => to_unsigned(609, 10), 8 => to_unsigned(141, 10), 9 => to_unsigned(627, 10), 10 => to_unsigned(130, 10), 11 => to_unsigned(813, 10), 12 => to_unsigned(456, 10), 13 => to_unsigned(541, 10), 14 => to_unsigned(341, 10), 15 => to_unsigned(240, 10), 16 => to_unsigned(479, 10), 17 => to_unsigned(310, 10), 18 => to_unsigned(567, 10), 19 => to_unsigned(328, 10), 20 => to_unsigned(434, 10), 21 => to_unsigned(815, 10), 22 => to_unsigned(312, 10), 23 => to_unsigned(870, 10), 24 => to_unsigned(891, 10), 25 => to_unsigned(852, 10), 26 => to_unsigned(280, 10), 27 => to_unsigned(988, 10), 28 => to_unsigned(430, 10), 29 => to_unsigned(239, 10), 30 => to_unsigned(618, 10), 31 => to_unsigned(142, 10), 32 => to_unsigned(149, 10), 33 => to_unsigned(857, 10), 34 => to_unsigned(980, 10), 35 => to_unsigned(183, 10), 36 => to_unsigned(252, 10), 37 => to_unsigned(224, 10), 38 => to_unsigned(596, 10), 39 => to_unsigned(1000, 10), 40 => to_unsigned(289, 10), 41 => to_unsigned(140, 10), 42 => to_unsigned(97, 10), 43 => to_unsigned(327, 10), 44 => to_unsigned(649, 10), 45 => to_unsigned(856, 10), 46 => to_unsigned(654, 10), 47 => to_unsigned(87, 10), 48 => to_unsigned(357, 10), 49 => to_unsigned(901, 10), 50 => to_unsigned(302, 10), 51 => to_unsigned(233, 10), 52 => to_unsigned(750, 10), 53 => to_unsigned(644, 10), 54 => to_unsigned(268, 10), 55 => to_unsigned(344, 10), 56 => to_unsigned(81, 10), 57 => to_unsigned(462, 10), 58 => to_unsigned(695, 10), 59 => to_unsigned(78, 10), 60 => to_unsigned(849, 10), 61 => to_unsigned(350, 10), 62 => to_unsigned(9, 10), 63 => to_unsigned(677, 10), 64 => to_unsigned(257, 10), 65 => to_unsigned(947, 10), 66 => to_unsigned(448, 10), 67 => to_unsigned(751, 10), 68 => to_unsigned(1010, 10), 69 => to_unsigned(538, 10), 70 => to_unsigned(395, 10), 71 => to_unsigned(807, 10), 72 => to_unsigned(169, 10), 73 => to_unsigned(468, 10), 74 => to_unsigned(153, 10), 75 => to_unsigned(109, 10), 76 => to_unsigned(801, 10), 77 => to_unsigned(498, 10), 78 => to_unsigned(307, 10), 79 => to_unsigned(758, 10), 80 => to_unsigned(120, 10), 81 => to_unsigned(277, 10), 82 => to_unsigned(637, 10), 83 => to_unsigned(566, 10), 84 => to_unsigned(591, 10), 85 => to_unsigned(353, 10), 86 => to_unsigned(368, 10), 87 => to_unsigned(896, 10), 88 => to_unsigned(779, 10), 89 => to_unsigned(220, 10), 90 => to_unsigned(801, 10), 91 => to_unsigned(1018, 10), 92 => to_unsigned(266, 10), 93 => to_unsigned(397, 10), 94 => to_unsigned(981, 10), 95 => to_unsigned(10, 10), 96 => to_unsigned(231, 10), 97 => to_unsigned(807, 10), 98 => to_unsigned(800, 10), 99 => to_unsigned(356, 10), 100 => to_unsigned(964, 10), 101 => to_unsigned(163, 10), 102 => to_unsigned(712, 10), 103 => to_unsigned(343, 10), 104 => to_unsigned(87, 10), 105 => to_unsigned(205, 10), 106 => to_unsigned(612, 10), 107 => to_unsigned(594, 10), 108 => to_unsigned(959, 10), 109 => to_unsigned(174, 10), 110 => to_unsigned(738, 10), 111 => to_unsigned(338, 10), 112 => to_unsigned(20, 10), 113 => to_unsigned(26, 10), 114 => to_unsigned(412, 10), 115 => to_unsigned(780, 10), 116 => to_unsigned(785, 10), 117 => to_unsigned(386, 10), 118 => to_unsigned(1012, 10), 119 => to_unsigned(804, 10), 120 => to_unsigned(970, 10), 121 => to_unsigned(546, 10), 122 => to_unsigned(935, 10), 123 => to_unsigned(10, 10), 124 => to_unsigned(563, 10), 125 => to_unsigned(130, 10), 126 => to_unsigned(193, 10), 127 => to_unsigned(919, 10), 128 => to_unsigned(384, 10), 129 => to_unsigned(380, 10), 130 => to_unsigned(842, 10), 131 => to_unsigned(507, 10), 132 => to_unsigned(68, 10), 133 => to_unsigned(404, 10), 134 => to_unsigned(697, 10), 135 => to_unsigned(261, 10), 136 => to_unsigned(747, 10), 137 => to_unsigned(868, 10), 138 => to_unsigned(761, 10), 139 => to_unsigned(750, 10), 140 => to_unsigned(515, 10), 141 => to_unsigned(365, 10), 142 => to_unsigned(781, 10), 143 => to_unsigned(606, 10), 144 => to_unsigned(171, 10), 145 => to_unsigned(258, 10), 146 => to_unsigned(379, 10), 147 => to_unsigned(929, 10), 148 => to_unsigned(379, 10), 149 => to_unsigned(411, 10), 150 => to_unsigned(517, 10), 151 => to_unsigned(563, 10), 152 => to_unsigned(461, 10), 153 => to_unsigned(933, 10), 154 => to_unsigned(791, 10), 155 => to_unsigned(143, 10), 156 => to_unsigned(586, 10), 157 => to_unsigned(732, 10), 158 => to_unsigned(419, 10), 159 => to_unsigned(920, 10), 160 => to_unsigned(606, 10), 161 => to_unsigned(445, 10), 162 => to_unsigned(309, 10), 163 => to_unsigned(255, 10), 164 => to_unsigned(876, 10), 165 => to_unsigned(87, 10), 166 => to_unsigned(392, 10), 167 => to_unsigned(925, 10), 168 => to_unsigned(350, 10), 169 => to_unsigned(99, 10), 170 => to_unsigned(458, 10), 171 => to_unsigned(878, 10), 172 => to_unsigned(921, 10), 173 => to_unsigned(389, 10), 174 => to_unsigned(493, 10), 175 => to_unsigned(645, 10), 176 => to_unsigned(100, 10), 177 => to_unsigned(670, 10), 178 => to_unsigned(771, 10), 179 => to_unsigned(376, 10), 180 => to_unsigned(11, 10), 181 => to_unsigned(185, 10), 182 => to_unsigned(27, 10), 183 => to_unsigned(1000, 10), 184 => to_unsigned(640, 10), 185 => to_unsigned(987, 10), 186 => to_unsigned(139, 10), 187 => to_unsigned(164, 10), 188 => to_unsigned(66, 10), 189 => to_unsigned(917, 10), 190 => to_unsigned(969, 10), 191 => to_unsigned(606, 10), 192 => to_unsigned(826, 10), 193 => to_unsigned(254, 10), 194 => to_unsigned(795, 10), 195 => to_unsigned(914, 10), 196 => to_unsigned(117, 10), 197 => to_unsigned(622, 10), 198 => to_unsigned(433, 10), 199 => to_unsigned(890, 10), 200 => to_unsigned(825, 10), 201 => to_unsigned(984, 10), 202 => to_unsigned(552, 10), 203 => to_unsigned(51, 10), 204 => to_unsigned(406, 10), 205 => to_unsigned(626, 10), 206 => to_unsigned(797, 10), 207 => to_unsigned(437, 10), 208 => to_unsigned(680, 10), 209 => to_unsigned(813, 10), 210 => to_unsigned(50, 10), 211 => to_unsigned(949, 10), 212 => to_unsigned(592, 10), 213 => to_unsigned(231, 10), 214 => to_unsigned(523, 10), 215 => to_unsigned(800, 10), 216 => to_unsigned(616, 10), 217 => to_unsigned(825, 10), 218 => to_unsigned(895, 10), 219 => to_unsigned(667, 10), 220 => to_unsigned(908, 10), 221 => to_unsigned(334, 10), 222 => to_unsigned(690, 10), 223 => to_unsigned(956, 10), 224 => to_unsigned(845, 10), 225 => to_unsigned(958, 10), 226 => to_unsigned(436, 10), 227 => to_unsigned(449, 10), 228 => to_unsigned(188, 10), 229 => to_unsigned(159, 10), 230 => to_unsigned(112, 10), 231 => to_unsigned(305, 10), 232 => to_unsigned(713, 10), 233 => to_unsigned(509, 10), 234 => to_unsigned(233, 10), 235 => to_unsigned(910, 10), 236 => to_unsigned(207, 10), 237 => to_unsigned(523, 10), 238 => to_unsigned(708, 10), 239 => to_unsigned(801, 10), 240 => to_unsigned(1005, 10), 241 => to_unsigned(184, 10), 242 => to_unsigned(760, 10), 243 => to_unsigned(425, 10), 244 => to_unsigned(667, 10), 245 => to_unsigned(434, 10), 246 => to_unsigned(607, 10), 247 => to_unsigned(145, 10), 248 => to_unsigned(399, 10), 249 => to_unsigned(422, 10), 250 => to_unsigned(898, 10), 251 => to_unsigned(853, 10), 252 => to_unsigned(675, 10), 253 => to_unsigned(529, 10), 254 => to_unsigned(423, 10), 255 => to_unsigned(734, 10), 256 => to_unsigned(703, 10), 257 => to_unsigned(505, 10), 258 => to_unsigned(120, 10), 259 => to_unsigned(305, 10), 260 => to_unsigned(137, 10), 261 => to_unsigned(25, 10), 262 => to_unsigned(669, 10), 263 => to_unsigned(240, 10), 264 => to_unsigned(450, 10), 265 => to_unsigned(624, 10), 266 => to_unsigned(512, 10), 267 => to_unsigned(433, 10), 268 => to_unsigned(217, 10), 269 => to_unsigned(239, 10), 270 => to_unsigned(773, 10), 271 => to_unsigned(852, 10), 272 => to_unsigned(653, 10), 273 => to_unsigned(805, 10), 274 => to_unsigned(84, 10), 275 => to_unsigned(619, 10), 276 => to_unsigned(798, 10), 277 => to_unsigned(444, 10), 278 => to_unsigned(313, 10), 279 => to_unsigned(507, 10), 280 => to_unsigned(642, 10), 281 => to_unsigned(421, 10), 282 => to_unsigned(436, 10), 283 => to_unsigned(406, 10), 284 => to_unsigned(93, 10), 285 => to_unsigned(852, 10), 286 => to_unsigned(65, 10), 287 => to_unsigned(41, 10), 288 => to_unsigned(376, 10), 289 => to_unsigned(86, 10), 290 => to_unsigned(950, 10), 291 => to_unsigned(455, 10), 292 => to_unsigned(38, 10), 293 => to_unsigned(400, 10), 294 => to_unsigned(948, 10), 295 => to_unsigned(604, 10), 296 => to_unsigned(179, 10), 297 => to_unsigned(237, 10), 298 => to_unsigned(87, 10), 299 => to_unsigned(540, 10), 300 => to_unsigned(174, 10), 301 => to_unsigned(137, 10), 302 => to_unsigned(425, 10), 303 => to_unsigned(667, 10), 304 => to_unsigned(911, 10), 305 => to_unsigned(282, 10), 306 => to_unsigned(975, 10), 307 => to_unsigned(1010, 10), 308 => to_unsigned(494, 10), 309 => to_unsigned(1017, 10), 310 => to_unsigned(654, 10), 311 => to_unsigned(998, 10), 312 => to_unsigned(656, 10), 313 => to_unsigned(669, 10), 314 => to_unsigned(445, 10), 315 => to_unsigned(978, 10), 316 => to_unsigned(518, 10), 317 => to_unsigned(504, 10), 318 => to_unsigned(55, 10), 319 => to_unsigned(577, 10), 320 => to_unsigned(81, 10), 321 => to_unsigned(640, 10), 322 => to_unsigned(414, 10), 323 => to_unsigned(49, 10), 324 => to_unsigned(1012, 10), 325 => to_unsigned(318, 10), 326 => to_unsigned(1, 10), 327 => to_unsigned(508, 10), 328 => to_unsigned(971, 10), 329 => to_unsigned(671, 10), 330 => to_unsigned(544, 10), 331 => to_unsigned(330, 10), 332 => to_unsigned(387, 10), 333 => to_unsigned(829, 10), 334 => to_unsigned(856, 10), 335 => to_unsigned(122, 10), 336 => to_unsigned(396, 10), 337 => to_unsigned(538, 10), 338 => to_unsigned(772, 10), 339 => to_unsigned(681, 10), 340 => to_unsigned(177, 10), 341 => to_unsigned(974, 10), 342 => to_unsigned(916, 10), 343 => to_unsigned(699, 10), 344 => to_unsigned(42, 10), 345 => to_unsigned(654, 10), 346 => to_unsigned(310, 10), 347 => to_unsigned(388, 10), 348 => to_unsigned(59, 10), 349 => to_unsigned(306, 10), 350 => to_unsigned(727, 10), 351 => to_unsigned(251, 10), 352 => to_unsigned(372, 10), 353 => to_unsigned(522, 10), 354 => to_unsigned(370, 10), 355 => to_unsigned(267, 10), 356 => to_unsigned(341, 10), 357 => to_unsigned(441, 10), 358 => to_unsigned(962, 10), 359 => to_unsigned(637, 10), 360 => to_unsigned(574, 10), 361 => to_unsigned(651, 10), 362 => to_unsigned(895, 10), 363 => to_unsigned(329, 10), 364 => to_unsigned(182, 10), 365 => to_unsigned(437, 10), 366 => to_unsigned(184, 10), 367 => to_unsigned(414, 10), 368 => to_unsigned(491, 10), 369 => to_unsigned(186, 10), 370 => to_unsigned(936, 10), 371 => to_unsigned(439, 10), 372 => to_unsigned(620, 10), 373 => to_unsigned(223, 10), 374 => to_unsigned(856, 10), 375 => to_unsigned(776, 10), 376 => to_unsigned(976, 10), 377 => to_unsigned(209, 10), 378 => to_unsigned(989, 10), 379 => to_unsigned(221, 10), 380 => to_unsigned(271, 10), 381 => to_unsigned(441, 10), 382 => to_unsigned(889, 10), 383 => to_unsigned(647, 10), 384 => to_unsigned(24, 10), 385 => to_unsigned(202, 10), 386 => to_unsigned(309, 10), 387 => to_unsigned(178, 10), 388 => to_unsigned(584, 10), 389 => to_unsigned(766, 10), 390 => to_unsigned(424, 10), 391 => to_unsigned(586, 10), 392 => to_unsigned(679, 10), 393 => to_unsigned(739, 10), 394 => to_unsigned(918, 10), 395 => to_unsigned(511, 10), 396 => to_unsigned(300, 10), 397 => to_unsigned(944, 10), 398 => to_unsigned(693, 10), 399 => to_unsigned(896, 10), 400 => to_unsigned(233, 10), 401 => to_unsigned(977, 10), 402 => to_unsigned(456, 10), 403 => to_unsigned(115, 10), 404 => to_unsigned(534, 10), 405 => to_unsigned(587, 10), 406 => to_unsigned(221, 10), 407 => to_unsigned(509, 10), 408 => to_unsigned(105, 10), 409 => to_unsigned(692, 10), 410 => to_unsigned(160, 10), 411 => to_unsigned(814, 10), 412 => to_unsigned(403, 10), 413 => to_unsigned(243, 10), 414 => to_unsigned(373, 10), 415 => to_unsigned(550, 10), 416 => to_unsigned(96, 10), 417 => to_unsigned(229, 10), 418 => to_unsigned(47, 10), 419 => to_unsigned(500, 10), 420 => to_unsigned(303, 10), 421 => to_unsigned(713, 10), 422 => to_unsigned(176, 10), 423 => to_unsigned(412, 10), 424 => to_unsigned(210, 10), 425 => to_unsigned(362, 10), 426 => to_unsigned(244, 10), 427 => to_unsigned(661, 10), 428 => to_unsigned(542, 10), 429 => to_unsigned(609, 10), 430 => to_unsigned(672, 10), 431 => to_unsigned(711, 10), 432 => to_unsigned(742, 10), 433 => to_unsigned(99, 10), 434 => to_unsigned(408, 10), 435 => to_unsigned(577, 10), 436 => to_unsigned(722, 10), 437 => to_unsigned(822, 10), 438 => to_unsigned(701, 10), 439 => to_unsigned(128, 10), 440 => to_unsigned(53, 10), 441 => to_unsigned(596, 10), 442 => to_unsigned(448, 10), 443 => to_unsigned(53, 10), 444 => to_unsigned(136, 10), 445 => to_unsigned(590, 10), 446 => to_unsigned(294, 10), 447 => to_unsigned(978, 10), 448 => to_unsigned(258, 10), 449 => to_unsigned(771, 10), 450 => to_unsigned(438, 10), 451 => to_unsigned(658, 10), 452 => to_unsigned(814, 10), 453 => to_unsigned(754, 10), 454 => to_unsigned(263, 10), 455 => to_unsigned(760, 10), 456 => to_unsigned(506, 10), 457 => to_unsigned(262, 10), 458 => to_unsigned(512, 10), 459 => to_unsigned(456, 10), 460 => to_unsigned(28, 10), 461 => to_unsigned(16, 10), 462 => to_unsigned(43, 10), 463 => to_unsigned(223, 10), 464 => to_unsigned(824, 10), 465 => to_unsigned(624, 10), 466 => to_unsigned(489, 10), 467 => to_unsigned(859, 10), 468 => to_unsigned(329, 10), 469 => to_unsigned(548, 10), 470 => to_unsigned(359, 10), 471 => to_unsigned(679, 10), 472 => to_unsigned(775, 10), 473 => to_unsigned(672, 10), 474 => to_unsigned(782, 10), 475 => to_unsigned(398, 10), 476 => to_unsigned(383, 10), 477 => to_unsigned(867, 10), 478 => to_unsigned(607, 10), 479 => to_unsigned(891, 10), 480 => to_unsigned(524, 10), 481 => to_unsigned(498, 10), 482 => to_unsigned(635, 10), 483 => to_unsigned(522, 10), 484 => to_unsigned(420, 10), 485 => to_unsigned(974, 10), 486 => to_unsigned(517, 10), 487 => to_unsigned(143, 10), 488 => to_unsigned(117, 10), 489 => to_unsigned(626, 10), 490 => to_unsigned(845, 10), 491 => to_unsigned(84, 10), 492 => to_unsigned(744, 10), 493 => to_unsigned(400, 10), 494 => to_unsigned(80, 10), 495 => to_unsigned(689, 10), 496 => to_unsigned(475, 10), 497 => to_unsigned(876, 10), 498 => to_unsigned(26, 10), 499 => to_unsigned(660, 10), 500 => to_unsigned(425, 10), 501 => to_unsigned(938, 10), 502 => to_unsigned(686, 10), 503 => to_unsigned(542, 10), 504 => to_unsigned(929, 10), 505 => to_unsigned(767, 10), 506 => to_unsigned(186, 10), 507 => to_unsigned(947, 10), 508 => to_unsigned(968, 10), 509 => to_unsigned(392, 10), 510 => to_unsigned(27, 10), 511 => to_unsigned(605, 10), 512 => to_unsigned(323, 10), 513 => to_unsigned(549, 10), 514 => to_unsigned(824, 10), 515 => to_unsigned(332, 10), 516 => to_unsigned(2, 10), 517 => to_unsigned(972, 10), 518 => to_unsigned(796, 10), 519 => to_unsigned(883, 10), 520 => to_unsigned(207, 10), 521 => to_unsigned(136, 10), 522 => to_unsigned(158, 10), 523 => to_unsigned(602, 10), 524 => to_unsigned(253, 10), 525 => to_unsigned(30, 10), 526 => to_unsigned(304, 10), 527 => to_unsigned(101, 10), 528 => to_unsigned(40, 10), 529 => to_unsigned(0, 10), 530 => to_unsigned(875, 10), 531 => to_unsigned(912, 10), 532 => to_unsigned(784, 10), 533 => to_unsigned(341, 10), 534 => to_unsigned(453, 10), 535 => to_unsigned(618, 10), 536 => to_unsigned(142, 10), 537 => to_unsigned(203, 10), 538 => to_unsigned(620, 10), 539 => to_unsigned(633, 10), 540 => to_unsigned(7, 10), 541 => to_unsigned(541, 10), 542 => to_unsigned(167, 10), 543 => to_unsigned(200, 10), 544 => to_unsigned(944, 10), 545 => to_unsigned(167, 10), 546 => to_unsigned(399, 10), 547 => to_unsigned(98, 10), 548 => to_unsigned(564, 10), 549 => to_unsigned(465, 10), 550 => to_unsigned(458, 10), 551 => to_unsigned(326, 10), 552 => to_unsigned(615, 10), 553 => to_unsigned(681, 10), 554 => to_unsigned(650, 10), 555 => to_unsigned(847, 10), 556 => to_unsigned(591, 10), 557 => to_unsigned(370, 10), 558 => to_unsigned(237, 10), 559 => to_unsigned(1014, 10), 560 => to_unsigned(147, 10), 561 => to_unsigned(554, 10), 562 => to_unsigned(941, 10), 563 => to_unsigned(860, 10), 564 => to_unsigned(323, 10), 565 => to_unsigned(361, 10), 566 => to_unsigned(814, 10), 567 => to_unsigned(214, 10), 568 => to_unsigned(429, 10), 569 => to_unsigned(539, 10), 570 => to_unsigned(429, 10), 571 => to_unsigned(585, 10), 572 => to_unsigned(281, 10), 573 => to_unsigned(145, 10), 574 => to_unsigned(826, 10), 575 => to_unsigned(293, 10), 576 => to_unsigned(68, 10), 577 => to_unsigned(275, 10), 578 => to_unsigned(697, 10), 579 => to_unsigned(132, 10), 580 => to_unsigned(574, 10), 581 => to_unsigned(369, 10), 582 => to_unsigned(617, 10), 583 => to_unsigned(144, 10), 584 => to_unsigned(849, 10), 585 => to_unsigned(384, 10), 586 => to_unsigned(432, 10), 587 => to_unsigned(287, 10), 588 => to_unsigned(1013, 10), 589 => to_unsigned(809, 10), 590 => to_unsigned(927, 10), 591 => to_unsigned(836, 10), 592 => to_unsigned(613, 10), 593 => to_unsigned(924, 10), 594 => to_unsigned(146, 10), 595 => to_unsigned(863, 10), 596 => to_unsigned(639, 10), 597 => to_unsigned(912, 10), 598 => to_unsigned(838, 10), 599 => to_unsigned(116, 10), 600 => to_unsigned(878, 10), 601 => to_unsigned(724, 10), 602 => to_unsigned(546, 10), 603 => to_unsigned(168, 10), 604 => to_unsigned(718, 10), 605 => to_unsigned(601, 10), 606 => to_unsigned(614, 10), 607 => to_unsigned(439, 10), 608 => to_unsigned(535, 10), 609 => to_unsigned(854, 10), 610 => to_unsigned(342, 10), 611 => to_unsigned(575, 10), 612 => to_unsigned(175, 10), 613 => to_unsigned(544, 10), 614 => to_unsigned(631, 10), 615 => to_unsigned(301, 10), 616 => to_unsigned(85, 10), 617 => to_unsigned(379, 10), 618 => to_unsigned(492, 10), 619 => to_unsigned(394, 10), 620 => to_unsigned(728, 10), 621 => to_unsigned(842, 10), 622 => to_unsigned(939, 10), 623 => to_unsigned(489, 10), 624 => to_unsigned(191, 10), 625 => to_unsigned(441, 10), 626 => to_unsigned(620, 10), 627 => to_unsigned(840, 10), 628 => to_unsigned(923, 10), 629 => to_unsigned(304, 10), 630 => to_unsigned(824, 10), 631 => to_unsigned(807, 10), 632 => to_unsigned(490, 10), 633 => to_unsigned(668, 10), 634 => to_unsigned(654, 10), 635 => to_unsigned(116, 10), 636 => to_unsigned(30, 10), 637 => to_unsigned(415, 10), 638 => to_unsigned(382, 10), 639 => to_unsigned(64, 10), 640 => to_unsigned(832, 10), 641 => to_unsigned(139, 10), 642 => to_unsigned(1015, 10), 643 => to_unsigned(293, 10), 644 => to_unsigned(640, 10), 645 => to_unsigned(631, 10), 646 => to_unsigned(876, 10), 647 => to_unsigned(290, 10), 648 => to_unsigned(891, 10), 649 => to_unsigned(18, 10), 650 => to_unsigned(800, 10), 651 => to_unsigned(422, 10), 652 => to_unsigned(927, 10), 653 => to_unsigned(395, 10), 654 => to_unsigned(893, 10), 655 => to_unsigned(118, 10), 656 => to_unsigned(215, 10), 657 => to_unsigned(210, 10), 658 => to_unsigned(923, 10), 659 => to_unsigned(801, 10), 660 => to_unsigned(777, 10), 661 => to_unsigned(901, 10), 662 => to_unsigned(708, 10), 663 => to_unsigned(510, 10), 664 => to_unsigned(643, 10), 665 => to_unsigned(109, 10), 666 => to_unsigned(459, 10), 667 => to_unsigned(524, 10), 668 => to_unsigned(841, 10), 669 => to_unsigned(139, 10), 670 => to_unsigned(909, 10), 671 => to_unsigned(1015, 10), 672 => to_unsigned(255, 10), 673 => to_unsigned(933, 10), 674 => to_unsigned(741, 10), 675 => to_unsigned(628, 10), 676 => to_unsigned(148, 10), 677 => to_unsigned(307, 10), 678 => to_unsigned(201, 10), 679 => to_unsigned(933, 10), 680 => to_unsigned(485, 10), 681 => to_unsigned(762, 10), 682 => to_unsigned(537, 10), 683 => to_unsigned(557, 10), 684 => to_unsigned(771, 10), 685 => to_unsigned(531, 10), 686 => to_unsigned(910, 10), 687 => to_unsigned(179, 10), 688 => to_unsigned(374, 10), 689 => to_unsigned(857, 10), 690 => to_unsigned(386, 10), 691 => to_unsigned(74, 10), 692 => to_unsigned(566, 10), 693 => to_unsigned(391, 10), 694 => to_unsigned(708, 10), 695 => to_unsigned(134, 10), 696 => to_unsigned(68, 10), 697 => to_unsigned(552, 10), 698 => to_unsigned(96, 10), 699 => to_unsigned(152, 10), 700 => to_unsigned(911, 10), 701 => to_unsigned(1016, 10), 702 => to_unsigned(50, 10), 703 => to_unsigned(918, 10), 704 => to_unsigned(867, 10), 705 => to_unsigned(335, 10), 706 => to_unsigned(982, 10), 707 => to_unsigned(494, 10), 708 => to_unsigned(714, 10), 709 => to_unsigned(178, 10), 710 => to_unsigned(164, 10), 711 => to_unsigned(146, 10), 712 => to_unsigned(622, 10), 713 => to_unsigned(693, 10), 714 => to_unsigned(384, 10), 715 => to_unsigned(325, 10), 716 => to_unsigned(893, 10), 717 => to_unsigned(580, 10), 718 => to_unsigned(168, 10), 719 => to_unsigned(172, 10), 720 => to_unsigned(12, 10), 721 => to_unsigned(5, 10), 722 => to_unsigned(521, 10), 723 => to_unsigned(796, 10), 724 => to_unsigned(769, 10), 725 => to_unsigned(123, 10), 726 => to_unsigned(478, 10), 727 => to_unsigned(279, 10), 728 => to_unsigned(208, 10), 729 => to_unsigned(527, 10), 730 => to_unsigned(38, 10), 731 => to_unsigned(450, 10), 732 => to_unsigned(351, 10), 733 => to_unsigned(987, 10), 734 => to_unsigned(610, 10), 735 => to_unsigned(694, 10), 736 => to_unsigned(62, 10), 737 => to_unsigned(224, 10), 738 => to_unsigned(402, 10), 739 => to_unsigned(844, 10), 740 => to_unsigned(411, 10), 741 => to_unsigned(559, 10), 742 => to_unsigned(469, 10), 743 => to_unsigned(601, 10), 744 => to_unsigned(938, 10), 745 => to_unsigned(219, 10), 746 => to_unsigned(49, 10), 747 => to_unsigned(127, 10), 748 => to_unsigned(168, 10), 749 => to_unsigned(1008, 10), 750 => to_unsigned(827, 10), 751 => to_unsigned(518, 10), 752 => to_unsigned(297, 10), 753 => to_unsigned(774, 10), 754 => to_unsigned(229, 10), 755 => to_unsigned(131, 10), 756 => to_unsigned(723, 10), 757 => to_unsigned(854, 10), 758 => to_unsigned(129, 10), 759 => to_unsigned(820, 10), 760 => to_unsigned(598, 10), 761 => to_unsigned(738, 10), 762 => to_unsigned(61, 10), 763 => to_unsigned(182, 10), 764 => to_unsigned(445, 10), 765 => to_unsigned(674, 10), 766 => to_unsigned(978, 10), 767 => to_unsigned(707, 10), 768 => to_unsigned(258, 10), 769 => to_unsigned(235, 10), 770 => to_unsigned(619, 10), 771 => to_unsigned(417, 10), 772 => to_unsigned(384, 10), 773 => to_unsigned(631, 10), 774 => to_unsigned(977, 10), 775 => to_unsigned(740, 10), 776 => to_unsigned(791, 10), 777 => to_unsigned(762, 10), 778 => to_unsigned(833, 10), 779 => to_unsigned(321, 10), 780 => to_unsigned(257, 10), 781 => to_unsigned(503, 10), 782 => to_unsigned(532, 10), 783 => to_unsigned(76, 10), 784 => to_unsigned(202, 10), 785 => to_unsigned(863, 10), 786 => to_unsigned(38, 10), 787 => to_unsigned(453, 10), 788 => to_unsigned(184, 10), 789 => to_unsigned(789, 10), 790 => to_unsigned(858, 10), 791 => to_unsigned(189, 10), 792 => to_unsigned(357, 10), 793 => to_unsigned(840, 10), 794 => to_unsigned(392, 10), 795 => to_unsigned(636, 10), 796 => to_unsigned(924, 10), 797 => to_unsigned(255, 10), 798 => to_unsigned(101, 10), 799 => to_unsigned(910, 10), 800 => to_unsigned(767, 10), 801 => to_unsigned(593, 10), 802 => to_unsigned(434, 10), 803 => to_unsigned(32, 10), 804 => to_unsigned(248, 10), 805 => to_unsigned(567, 10), 806 => to_unsigned(728, 10), 807 => to_unsigned(774, 10), 808 => to_unsigned(1013, 10), 809 => to_unsigned(255, 10), 810 => to_unsigned(15, 10), 811 => to_unsigned(233, 10), 812 => to_unsigned(356, 10), 813 => to_unsigned(783, 10), 814 => to_unsigned(604, 10), 815 => to_unsigned(729, 10), 816 => to_unsigned(398, 10), 817 => to_unsigned(790, 10), 818 => to_unsigned(706, 10), 819 => to_unsigned(986, 10), 820 => to_unsigned(529, 10), 821 => to_unsigned(492, 10), 822 => to_unsigned(47, 10), 823 => to_unsigned(658, 10), 824 => to_unsigned(88, 10), 825 => to_unsigned(776, 10), 826 => to_unsigned(884, 10), 827 => to_unsigned(662, 10), 828 => to_unsigned(217, 10), 829 => to_unsigned(329, 10), 830 => to_unsigned(783, 10), 831 => to_unsigned(735, 10), 832 => to_unsigned(754, 10), 833 => to_unsigned(1004, 10), 834 => to_unsigned(444, 10), 835 => to_unsigned(813, 10), 836 => to_unsigned(538, 10), 837 => to_unsigned(911, 10), 838 => to_unsigned(196, 10), 839 => to_unsigned(383, 10), 840 => to_unsigned(236, 10), 841 => to_unsigned(125, 10), 842 => to_unsigned(650, 10), 843 => to_unsigned(852, 10), 844 => to_unsigned(175, 10), 845 => to_unsigned(942, 10), 846 => to_unsigned(885, 10), 847 => to_unsigned(303, 10), 848 => to_unsigned(581, 10), 849 => to_unsigned(558, 10), 850 => to_unsigned(794, 10), 851 => to_unsigned(605, 10), 852 => to_unsigned(501, 10), 853 => to_unsigned(429, 10), 854 => to_unsigned(519, 10), 855 => to_unsigned(771, 10), 856 => to_unsigned(921, 10), 857 => to_unsigned(705, 10), 858 => to_unsigned(284, 10), 859 => to_unsigned(847, 10), 860 => to_unsigned(880, 10), 861 => to_unsigned(583, 10), 862 => to_unsigned(48, 10), 863 => to_unsigned(255, 10), 864 => to_unsigned(870, 10), 865 => to_unsigned(711, 10), 866 => to_unsigned(353, 10), 867 => to_unsigned(774, 10), 868 => to_unsigned(504, 10), 869 => to_unsigned(338, 10), 870 => to_unsigned(546, 10), 871 => to_unsigned(165, 10), 872 => to_unsigned(869, 10), 873 => to_unsigned(611, 10), 874 => to_unsigned(744, 10), 875 => to_unsigned(785, 10), 876 => to_unsigned(107, 10), 877 => to_unsigned(447, 10), 878 => to_unsigned(406, 10), 879 => to_unsigned(932, 10), 880 => to_unsigned(18, 10), 881 => to_unsigned(585, 10), 882 => to_unsigned(133, 10), 883 => to_unsigned(135, 10), 884 => to_unsigned(534, 10), 885 => to_unsigned(273, 10), 886 => to_unsigned(168, 10), 887 => to_unsigned(81, 10), 888 => to_unsigned(92, 10), 889 => to_unsigned(830, 10), 890 => to_unsigned(216, 10), 891 => to_unsigned(672, 10), 892 => to_unsigned(891, 10), 893 => to_unsigned(688, 10), 894 => to_unsigned(739, 10), 895 => to_unsigned(924, 10), 896 => to_unsigned(409, 10), 897 => to_unsigned(669, 10), 898 => to_unsigned(156, 10), 899 => to_unsigned(215, 10), 900 => to_unsigned(504, 10), 901 => to_unsigned(958, 10), 902 => to_unsigned(585, 10), 903 => to_unsigned(877, 10), 904 => to_unsigned(585, 10), 905 => to_unsigned(202, 10), 906 => to_unsigned(277, 10), 907 => to_unsigned(918, 10), 908 => to_unsigned(636, 10), 909 => to_unsigned(475, 10), 910 => to_unsigned(516, 10), 911 => to_unsigned(822, 10), 912 => to_unsigned(231, 10), 913 => to_unsigned(780, 10), 914 => to_unsigned(193, 10), 915 => to_unsigned(652, 10), 916 => to_unsigned(148, 10), 917 => to_unsigned(141, 10), 918 => to_unsigned(756, 10), 919 => to_unsigned(26, 10), 920 => to_unsigned(705, 10), 921 => to_unsigned(883, 10), 922 => to_unsigned(1008, 10), 923 => to_unsigned(353, 10), 924 => to_unsigned(517, 10), 925 => to_unsigned(686, 10), 926 => to_unsigned(970, 10), 927 => to_unsigned(291, 10), 928 => to_unsigned(104, 10), 929 => to_unsigned(409, 10), 930 => to_unsigned(47, 10), 931 => to_unsigned(512, 10), 932 => to_unsigned(149, 10), 933 => to_unsigned(647, 10), 934 => to_unsigned(770, 10), 935 => to_unsigned(644, 10), 936 => to_unsigned(696, 10), 937 => to_unsigned(369, 10), 938 => to_unsigned(890, 10), 939 => to_unsigned(34, 10), 940 => to_unsigned(510, 10), 941 => to_unsigned(54, 10), 942 => to_unsigned(22, 10), 943 => to_unsigned(207, 10), 944 => to_unsigned(405, 10), 945 => to_unsigned(1005, 10), 946 => to_unsigned(386, 10), 947 => to_unsigned(847, 10), 948 => to_unsigned(820, 10), 949 => to_unsigned(279, 10), 950 => to_unsigned(350, 10), 951 => to_unsigned(173, 10), 952 => to_unsigned(764, 10), 953 => to_unsigned(829, 10), 954 => to_unsigned(246, 10), 955 => to_unsigned(753, 10), 956 => to_unsigned(786, 10), 957 => to_unsigned(283, 10), 958 => to_unsigned(210, 10), 959 => to_unsigned(649, 10), 960 => to_unsigned(453, 10), 961 => to_unsigned(482, 10), 962 => to_unsigned(122, 10), 963 => to_unsigned(23, 10), 964 => to_unsigned(839, 10), 965 => to_unsigned(414, 10), 966 => to_unsigned(359, 10), 967 => to_unsigned(363, 10), 968 => to_unsigned(137, 10), 969 => to_unsigned(466, 10), 970 => to_unsigned(276, 10), 971 => to_unsigned(592, 10), 972 => to_unsigned(243, 10), 973 => to_unsigned(109, 10), 974 => to_unsigned(619, 10), 975 => to_unsigned(982, 10), 976 => to_unsigned(913, 10), 977 => to_unsigned(476, 10), 978 => to_unsigned(476, 10), 979 => to_unsigned(812, 10), 980 => to_unsigned(401, 10), 981 => to_unsigned(553, 10), 982 => to_unsigned(777, 10), 983 => to_unsigned(23, 10), 984 => to_unsigned(205, 10), 985 => to_unsigned(455, 10), 986 => to_unsigned(1023, 10), 987 => to_unsigned(474, 10), 988 => to_unsigned(410, 10), 989 => to_unsigned(147, 10), 990 => to_unsigned(323, 10), 991 => to_unsigned(696, 10), 992 => to_unsigned(264, 10), 993 => to_unsigned(46, 10), 994 => to_unsigned(251, 10), 995 => to_unsigned(456, 10), 996 => to_unsigned(642, 10), 997 => to_unsigned(891, 10), 998 => to_unsigned(517, 10), 999 => to_unsigned(398, 10), 1000 => to_unsigned(161, 10), 1001 => to_unsigned(68, 10), 1002 => to_unsigned(246, 10), 1003 => to_unsigned(737, 10), 1004 => to_unsigned(360, 10), 1005 => to_unsigned(65, 10), 1006 => to_unsigned(819, 10), 1007 => to_unsigned(811, 10), 1008 => to_unsigned(248, 10), 1009 => to_unsigned(878, 10), 1010 => to_unsigned(387, 10), 1011 => to_unsigned(361, 10), 1012 => to_unsigned(52, 10), 1013 => to_unsigned(472, 10), 1014 => to_unsigned(4, 10), 1015 => to_unsigned(538, 10), 1016 => to_unsigned(414, 10), 1017 => to_unsigned(164, 10), 1018 => to_unsigned(686, 10), 1019 => to_unsigned(891, 10), 1020 => to_unsigned(969, 10), 1021 => to_unsigned(519, 10), 1022 => to_unsigned(412, 10), 1023 => to_unsigned(108, 10), 1024 => to_unsigned(270, 10), 1025 => to_unsigned(697, 10), 1026 => to_unsigned(126, 10), 1027 => to_unsigned(415, 10), 1028 => to_unsigned(808, 10), 1029 => to_unsigned(705, 10), 1030 => to_unsigned(725, 10), 1031 => to_unsigned(405, 10), 1032 => to_unsigned(102, 10), 1033 => to_unsigned(479, 10), 1034 => to_unsigned(722, 10), 1035 => to_unsigned(1020, 10), 1036 => to_unsigned(31, 10), 1037 => to_unsigned(737, 10), 1038 => to_unsigned(902, 10), 1039 => to_unsigned(924, 10), 1040 => to_unsigned(728, 10), 1041 => to_unsigned(980, 10), 1042 => to_unsigned(284, 10), 1043 => to_unsigned(17, 10), 1044 => to_unsigned(39, 10), 1045 => to_unsigned(144, 10), 1046 => to_unsigned(58, 10), 1047 => to_unsigned(1, 10), 1048 => to_unsigned(873, 10), 1049 => to_unsigned(309, 10), 1050 => to_unsigned(837, 10), 1051 => to_unsigned(311, 10), 1052 => to_unsigned(824, 10), 1053 => to_unsigned(99, 10), 1054 => to_unsigned(420, 10), 1055 => to_unsigned(505, 10), 1056 => to_unsigned(671, 10), 1057 => to_unsigned(616, 10), 1058 => to_unsigned(893, 10), 1059 => to_unsigned(577, 10), 1060 => to_unsigned(360, 10), 1061 => to_unsigned(735, 10), 1062 => to_unsigned(224, 10), 1063 => to_unsigned(658, 10), 1064 => to_unsigned(232, 10), 1065 => to_unsigned(798, 10), 1066 => to_unsigned(782, 10), 1067 => to_unsigned(725, 10), 1068 => to_unsigned(223, 10), 1069 => to_unsigned(416, 10), 1070 => to_unsigned(139, 10), 1071 => to_unsigned(870, 10), 1072 => to_unsigned(236, 10), 1073 => to_unsigned(78, 10), 1074 => to_unsigned(783, 10), 1075 => to_unsigned(647, 10), 1076 => to_unsigned(967, 10), 1077 => to_unsigned(330, 10), 1078 => to_unsigned(446, 10), 1079 => to_unsigned(852, 10), 1080 => to_unsigned(161, 10), 1081 => to_unsigned(503, 10), 1082 => to_unsigned(18, 10), 1083 => to_unsigned(511, 10), 1084 => to_unsigned(170, 10), 1085 => to_unsigned(1000, 10), 1086 => to_unsigned(155, 10), 1087 => to_unsigned(792, 10), 1088 => to_unsigned(69, 10), 1089 => to_unsigned(195, 10), 1090 => to_unsigned(925, 10), 1091 => to_unsigned(670, 10), 1092 => to_unsigned(95, 10), 1093 => to_unsigned(802, 10), 1094 => to_unsigned(26, 10), 1095 => to_unsigned(963, 10), 1096 => to_unsigned(496, 10), 1097 => to_unsigned(23, 10), 1098 => to_unsigned(200, 10), 1099 => to_unsigned(490, 10), 1100 => to_unsigned(920, 10), 1101 => to_unsigned(1002, 10), 1102 => to_unsigned(390, 10), 1103 => to_unsigned(842, 10), 1104 => to_unsigned(893, 10), 1105 => to_unsigned(889, 10), 1106 => to_unsigned(1007, 10), 1107 => to_unsigned(611, 10), 1108 => to_unsigned(427, 10), 1109 => to_unsigned(622, 10), 1110 => to_unsigned(249, 10), 1111 => to_unsigned(231, 10), 1112 => to_unsigned(751, 10), 1113 => to_unsigned(241, 10), 1114 => to_unsigned(564, 10), 1115 => to_unsigned(730, 10), 1116 => to_unsigned(45, 10), 1117 => to_unsigned(484, 10), 1118 => to_unsigned(463, 10), 1119 => to_unsigned(914, 10), 1120 => to_unsigned(771, 10), 1121 => to_unsigned(988, 10), 1122 => to_unsigned(319, 10), 1123 => to_unsigned(186, 10), 1124 => to_unsigned(447, 10), 1125 => to_unsigned(423, 10), 1126 => to_unsigned(478, 10), 1127 => to_unsigned(389, 10), 1128 => to_unsigned(431, 10), 1129 => to_unsigned(662, 10), 1130 => to_unsigned(619, 10), 1131 => to_unsigned(51, 10), 1132 => to_unsigned(561, 10), 1133 => to_unsigned(585, 10), 1134 => to_unsigned(908, 10), 1135 => to_unsigned(416, 10), 1136 => to_unsigned(335, 10), 1137 => to_unsigned(1014, 10), 1138 => to_unsigned(800, 10), 1139 => to_unsigned(803, 10), 1140 => to_unsigned(498, 10), 1141 => to_unsigned(764, 10), 1142 => to_unsigned(510, 10), 1143 => to_unsigned(572, 10), 1144 => to_unsigned(830, 10), 1145 => to_unsigned(495, 10), 1146 => to_unsigned(348, 10), 1147 => to_unsigned(383, 10), 1148 => to_unsigned(474, 10), 1149 => to_unsigned(739, 10), 1150 => to_unsigned(594, 10), 1151 => to_unsigned(428, 10), 1152 => to_unsigned(234, 10), 1153 => to_unsigned(435, 10), 1154 => to_unsigned(568, 10), 1155 => to_unsigned(476, 10), 1156 => to_unsigned(264, 10), 1157 => to_unsigned(945, 10), 1158 => to_unsigned(560, 10), 1159 => to_unsigned(1021, 10), 1160 => to_unsigned(183, 10), 1161 => to_unsigned(662, 10), 1162 => to_unsigned(574, 10), 1163 => to_unsigned(479, 10), 1164 => to_unsigned(825, 10), 1165 => to_unsigned(725, 10), 1166 => to_unsigned(290, 10), 1167 => to_unsigned(951, 10), 1168 => to_unsigned(809, 10), 1169 => to_unsigned(704, 10), 1170 => to_unsigned(299, 10), 1171 => to_unsigned(11, 10), 1172 => to_unsigned(136, 10), 1173 => to_unsigned(919, 10), 1174 => to_unsigned(568, 10), 1175 => to_unsigned(981, 10), 1176 => to_unsigned(1017, 10), 1177 => to_unsigned(568, 10), 1178 => to_unsigned(240, 10), 1179 => to_unsigned(311, 10), 1180 => to_unsigned(878, 10), 1181 => to_unsigned(93, 10), 1182 => to_unsigned(381, 10), 1183 => to_unsigned(136, 10), 1184 => to_unsigned(277, 10), 1185 => to_unsigned(888, 10), 1186 => to_unsigned(244, 10), 1187 => to_unsigned(716, 10), 1188 => to_unsigned(493, 10), 1189 => to_unsigned(683, 10), 1190 => to_unsigned(393, 10), 1191 => to_unsigned(251, 10), 1192 => to_unsigned(203, 10), 1193 => to_unsigned(33, 10), 1194 => to_unsigned(45, 10), 1195 => to_unsigned(1001, 10), 1196 => to_unsigned(51, 10), 1197 => to_unsigned(752, 10), 1198 => to_unsigned(728, 10), 1199 => to_unsigned(327, 10), 1200 => to_unsigned(725, 10), 1201 => to_unsigned(797, 10), 1202 => to_unsigned(746, 10), 1203 => to_unsigned(231, 10), 1204 => to_unsigned(358, 10), 1205 => to_unsigned(983, 10), 1206 => to_unsigned(66, 10), 1207 => to_unsigned(170, 10), 1208 => to_unsigned(37, 10), 1209 => to_unsigned(883, 10), 1210 => to_unsigned(753, 10), 1211 => to_unsigned(326, 10), 1212 => to_unsigned(916, 10), 1213 => to_unsigned(49, 10), 1214 => to_unsigned(740, 10), 1215 => to_unsigned(550, 10), 1216 => to_unsigned(725, 10), 1217 => to_unsigned(681, 10), 1218 => to_unsigned(381, 10), 1219 => to_unsigned(337, 10), 1220 => to_unsigned(380, 10), 1221 => to_unsigned(160, 10), 1222 => to_unsigned(47, 10), 1223 => to_unsigned(594, 10), 1224 => to_unsigned(795, 10), 1225 => to_unsigned(843, 10), 1226 => to_unsigned(725, 10), 1227 => to_unsigned(328, 10), 1228 => to_unsigned(574, 10), 1229 => to_unsigned(855, 10), 1230 => to_unsigned(680, 10), 1231 => to_unsigned(211, 10), 1232 => to_unsigned(660, 10), 1233 => to_unsigned(731, 10), 1234 => to_unsigned(253, 10), 1235 => to_unsigned(902, 10), 1236 => to_unsigned(937, 10), 1237 => to_unsigned(92, 10), 1238 => to_unsigned(112, 10), 1239 => to_unsigned(331, 10), 1240 => to_unsigned(6, 10), 1241 => to_unsigned(336, 10), 1242 => to_unsigned(671, 10), 1243 => to_unsigned(941, 10), 1244 => to_unsigned(967, 10), 1245 => to_unsigned(420, 10), 1246 => to_unsigned(25, 10), 1247 => to_unsigned(541, 10), 1248 => to_unsigned(502, 10), 1249 => to_unsigned(126, 10), 1250 => to_unsigned(639, 10), 1251 => to_unsigned(430, 10), 1252 => to_unsigned(581, 10), 1253 => to_unsigned(185, 10), 1254 => to_unsigned(191, 10), 1255 => to_unsigned(584, 10), 1256 => to_unsigned(324, 10), 1257 => to_unsigned(289, 10), 1258 => to_unsigned(421, 10), 1259 => to_unsigned(897, 10), 1260 => to_unsigned(663, 10), 1261 => to_unsigned(49, 10), 1262 => to_unsigned(524, 10), 1263 => to_unsigned(1, 10), 1264 => to_unsigned(583, 10), 1265 => to_unsigned(348, 10), 1266 => to_unsigned(648, 10), 1267 => to_unsigned(174, 10), 1268 => to_unsigned(932, 10), 1269 => to_unsigned(816, 10), 1270 => to_unsigned(440, 10), 1271 => to_unsigned(169, 10), 1272 => to_unsigned(600, 10), 1273 => to_unsigned(576, 10), 1274 => to_unsigned(738, 10), 1275 => to_unsigned(45, 10), 1276 => to_unsigned(429, 10), 1277 => to_unsigned(271, 10), 1278 => to_unsigned(551, 10), 1279 => to_unsigned(770, 10), 1280 => to_unsigned(810, 10), 1281 => to_unsigned(267, 10), 1282 => to_unsigned(879, 10), 1283 => to_unsigned(964, 10), 1284 => to_unsigned(863, 10), 1285 => to_unsigned(494, 10), 1286 => to_unsigned(710, 10), 1287 => to_unsigned(700, 10), 1288 => to_unsigned(450, 10), 1289 => to_unsigned(57, 10), 1290 => to_unsigned(714, 10), 1291 => to_unsigned(484, 10), 1292 => to_unsigned(170, 10), 1293 => to_unsigned(685, 10), 1294 => to_unsigned(721, 10), 1295 => to_unsigned(110, 10), 1296 => to_unsigned(460, 10), 1297 => to_unsigned(232, 10), 1298 => to_unsigned(785, 10), 1299 => to_unsigned(943, 10), 1300 => to_unsigned(693, 10), 1301 => to_unsigned(391, 10), 1302 => to_unsigned(843, 10), 1303 => to_unsigned(410, 10), 1304 => to_unsigned(278, 10), 1305 => to_unsigned(228, 10), 1306 => to_unsigned(625, 10), 1307 => to_unsigned(475, 10), 1308 => to_unsigned(636, 10), 1309 => to_unsigned(76, 10), 1310 => to_unsigned(199, 10), 1311 => to_unsigned(978, 10), 1312 => to_unsigned(831, 10), 1313 => to_unsigned(593, 10), 1314 => to_unsigned(566, 10), 1315 => to_unsigned(135, 10), 1316 => to_unsigned(182, 10), 1317 => to_unsigned(199, 10), 1318 => to_unsigned(904, 10), 1319 => to_unsigned(84, 10), 1320 => to_unsigned(561, 10), 1321 => to_unsigned(11, 10), 1322 => to_unsigned(472, 10), 1323 => to_unsigned(124, 10), 1324 => to_unsigned(434, 10), 1325 => to_unsigned(410, 10), 1326 => to_unsigned(781, 10), 1327 => to_unsigned(112, 10), 1328 => to_unsigned(556, 10), 1329 => to_unsigned(140, 10), 1330 => to_unsigned(587, 10), 1331 => to_unsigned(206, 10), 1332 => to_unsigned(275, 10), 1333 => to_unsigned(162, 10), 1334 => to_unsigned(786, 10), 1335 => to_unsigned(614, 10), 1336 => to_unsigned(956, 10), 1337 => to_unsigned(449, 10), 1338 => to_unsigned(543, 10), 1339 => to_unsigned(581, 10), 1340 => to_unsigned(307, 10), 1341 => to_unsigned(231, 10), 1342 => to_unsigned(240, 10), 1343 => to_unsigned(904, 10), 1344 => to_unsigned(416, 10), 1345 => to_unsigned(122, 10), 1346 => to_unsigned(262, 10), 1347 => to_unsigned(929, 10), 1348 => to_unsigned(512, 10), 1349 => to_unsigned(634, 10), 1350 => to_unsigned(131, 10), 1351 => to_unsigned(63, 10), 1352 => to_unsigned(507, 10), 1353 => to_unsigned(425, 10), 1354 => to_unsigned(181, 10), 1355 => to_unsigned(815, 10), 1356 => to_unsigned(570, 10), 1357 => to_unsigned(965, 10), 1358 => to_unsigned(44, 10), 1359 => to_unsigned(635, 10), 1360 => to_unsigned(98, 10), 1361 => to_unsigned(385, 10), 1362 => to_unsigned(103, 10), 1363 => to_unsigned(651, 10), 1364 => to_unsigned(754, 10), 1365 => to_unsigned(909, 10), 1366 => to_unsigned(524, 10), 1367 => to_unsigned(76, 10), 1368 => to_unsigned(17, 10), 1369 => to_unsigned(443, 10), 1370 => to_unsigned(425, 10), 1371 => to_unsigned(308, 10), 1372 => to_unsigned(345, 10), 1373 => to_unsigned(235, 10), 1374 => to_unsigned(291, 10), 1375 => to_unsigned(666, 10), 1376 => to_unsigned(311, 10), 1377 => to_unsigned(446, 10), 1378 => to_unsigned(994, 10), 1379 => to_unsigned(693, 10), 1380 => to_unsigned(328, 10), 1381 => to_unsigned(170, 10), 1382 => to_unsigned(455, 10), 1383 => to_unsigned(13, 10), 1384 => to_unsigned(392, 10), 1385 => to_unsigned(538, 10), 1386 => to_unsigned(83, 10), 1387 => to_unsigned(687, 10), 1388 => to_unsigned(371, 10), 1389 => to_unsigned(697, 10), 1390 => to_unsigned(414, 10), 1391 => to_unsigned(203, 10), 1392 => to_unsigned(694, 10), 1393 => to_unsigned(627, 10), 1394 => to_unsigned(440, 10), 1395 => to_unsigned(49, 10), 1396 => to_unsigned(995, 10), 1397 => to_unsigned(659, 10), 1398 => to_unsigned(150, 10), 1399 => to_unsigned(612, 10), 1400 => to_unsigned(915, 10), 1401 => to_unsigned(884, 10), 1402 => to_unsigned(943, 10), 1403 => to_unsigned(434, 10), 1404 => to_unsigned(482, 10), 1405 => to_unsigned(1019, 10), 1406 => to_unsigned(73, 10), 1407 => to_unsigned(299, 10), 1408 => to_unsigned(18, 10), 1409 => to_unsigned(564, 10), 1410 => to_unsigned(108, 10), 1411 => to_unsigned(517, 10), 1412 => to_unsigned(538, 10), 1413 => to_unsigned(271, 10), 1414 => to_unsigned(415, 10), 1415 => to_unsigned(11, 10), 1416 => to_unsigned(2, 10), 1417 => to_unsigned(183, 10), 1418 => to_unsigned(170, 10), 1419 => to_unsigned(636, 10), 1420 => to_unsigned(206, 10), 1421 => to_unsigned(652, 10), 1422 => to_unsigned(458, 10), 1423 => to_unsigned(711, 10), 1424 => to_unsigned(406, 10), 1425 => to_unsigned(55, 10), 1426 => to_unsigned(463, 10), 1427 => to_unsigned(948, 10), 1428 => to_unsigned(323, 10), 1429 => to_unsigned(975, 10), 1430 => to_unsigned(107, 10), 1431 => to_unsigned(480, 10), 1432 => to_unsigned(386, 10), 1433 => to_unsigned(1023, 10), 1434 => to_unsigned(1023, 10), 1435 => to_unsigned(878, 10), 1436 => to_unsigned(665, 10), 1437 => to_unsigned(621, 10), 1438 => to_unsigned(827, 10), 1439 => to_unsigned(774, 10), 1440 => to_unsigned(909, 10), 1441 => to_unsigned(366, 10), 1442 => to_unsigned(716, 10), 1443 => to_unsigned(754, 10), 1444 => to_unsigned(121, 10), 1445 => to_unsigned(633, 10), 1446 => to_unsigned(606, 10), 1447 => to_unsigned(985, 10), 1448 => to_unsigned(302, 10), 1449 => to_unsigned(641, 10), 1450 => to_unsigned(823, 10), 1451 => to_unsigned(79, 10), 1452 => to_unsigned(435, 10), 1453 => to_unsigned(456, 10), 1454 => to_unsigned(620, 10), 1455 => to_unsigned(219, 10), 1456 => to_unsigned(64, 10), 1457 => to_unsigned(43, 10), 1458 => to_unsigned(36, 10), 1459 => to_unsigned(315, 10), 1460 => to_unsigned(92, 10), 1461 => to_unsigned(298, 10), 1462 => to_unsigned(427, 10), 1463 => to_unsigned(234, 10), 1464 => to_unsigned(211, 10), 1465 => to_unsigned(802, 10), 1466 => to_unsigned(837, 10), 1467 => to_unsigned(98, 10), 1468 => to_unsigned(290, 10), 1469 => to_unsigned(961, 10), 1470 => to_unsigned(224, 10), 1471 => to_unsigned(768, 10), 1472 => to_unsigned(575, 10), 1473 => to_unsigned(869, 10), 1474 => to_unsigned(130, 10), 1475 => to_unsigned(127, 10), 1476 => to_unsigned(581, 10), 1477 => to_unsigned(569, 10), 1478 => to_unsigned(633, 10), 1479 => to_unsigned(204, 10), 1480 => to_unsigned(129, 10), 1481 => to_unsigned(775, 10), 1482 => to_unsigned(807, 10), 1483 => to_unsigned(930, 10), 1484 => to_unsigned(876, 10), 1485 => to_unsigned(351, 10), 1486 => to_unsigned(728, 10), 1487 => to_unsigned(590, 10), 1488 => to_unsigned(696, 10), 1489 => to_unsigned(51, 10), 1490 => to_unsigned(882, 10), 1491 => to_unsigned(479, 10), 1492 => to_unsigned(374, 10), 1493 => to_unsigned(789, 10), 1494 => to_unsigned(979, 10), 1495 => to_unsigned(543, 10), 1496 => to_unsigned(471, 10), 1497 => to_unsigned(560, 10), 1498 => to_unsigned(561, 10), 1499 => to_unsigned(956, 10), 1500 => to_unsigned(829, 10), 1501 => to_unsigned(227, 10), 1502 => to_unsigned(50, 10), 1503 => to_unsigned(32, 10), 1504 => to_unsigned(320, 10), 1505 => to_unsigned(357, 10), 1506 => to_unsigned(276, 10), 1507 => to_unsigned(968, 10), 1508 => to_unsigned(381, 10), 1509 => to_unsigned(683, 10), 1510 => to_unsigned(453, 10), 1511 => to_unsigned(424, 10), 1512 => to_unsigned(368, 10), 1513 => to_unsigned(380, 10), 1514 => to_unsigned(921, 10), 1515 => to_unsigned(119, 10), 1516 => to_unsigned(966, 10), 1517 => to_unsigned(765, 10), 1518 => to_unsigned(274, 10), 1519 => to_unsigned(471, 10), 1520 => to_unsigned(69, 10), 1521 => to_unsigned(970, 10), 1522 => to_unsigned(867, 10), 1523 => to_unsigned(821, 10), 1524 => to_unsigned(306, 10), 1525 => to_unsigned(276, 10), 1526 => to_unsigned(508, 10), 1527 => to_unsigned(64, 10), 1528 => to_unsigned(429, 10), 1529 => to_unsigned(607, 10), 1530 => to_unsigned(7, 10), 1531 => to_unsigned(592, 10), 1532 => to_unsigned(611, 10), 1533 => to_unsigned(613, 10), 1534 => to_unsigned(337, 10), 1535 => to_unsigned(958, 10), 1536 => to_unsigned(183, 10), 1537 => to_unsigned(848, 10), 1538 => to_unsigned(916, 10), 1539 => to_unsigned(632, 10), 1540 => to_unsigned(291, 10), 1541 => to_unsigned(163, 10), 1542 => to_unsigned(23, 10), 1543 => to_unsigned(472, 10), 1544 => to_unsigned(825, 10), 1545 => to_unsigned(138, 10), 1546 => to_unsigned(661, 10), 1547 => to_unsigned(596, 10), 1548 => to_unsigned(873, 10), 1549 => to_unsigned(219, 10), 1550 => to_unsigned(148, 10), 1551 => to_unsigned(357, 10), 1552 => to_unsigned(367, 10), 1553 => to_unsigned(468, 10), 1554 => to_unsigned(594, 10), 1555 => to_unsigned(19, 10), 1556 => to_unsigned(330, 10), 1557 => to_unsigned(71, 10), 1558 => to_unsigned(426, 10), 1559 => to_unsigned(447, 10), 1560 => to_unsigned(617, 10), 1561 => to_unsigned(479, 10), 1562 => to_unsigned(462, 10), 1563 => to_unsigned(349, 10), 1564 => to_unsigned(691, 10), 1565 => to_unsigned(115, 10), 1566 => to_unsigned(31, 10), 1567 => to_unsigned(929, 10), 1568 => to_unsigned(990, 10), 1569 => to_unsigned(103, 10), 1570 => to_unsigned(374, 10), 1571 => to_unsigned(1003, 10), 1572 => to_unsigned(417, 10), 1573 => to_unsigned(635, 10), 1574 => to_unsigned(29, 10), 1575 => to_unsigned(904, 10), 1576 => to_unsigned(419, 10), 1577 => to_unsigned(646, 10), 1578 => to_unsigned(328, 10), 1579 => to_unsigned(255, 10), 1580 => to_unsigned(365, 10), 1581 => to_unsigned(162, 10), 1582 => to_unsigned(202, 10), 1583 => to_unsigned(446, 10), 1584 => to_unsigned(954, 10), 1585 => to_unsigned(244, 10), 1586 => to_unsigned(818, 10), 1587 => to_unsigned(614, 10), 1588 => to_unsigned(792, 10), 1589 => to_unsigned(573, 10), 1590 => to_unsigned(921, 10), 1591 => to_unsigned(222, 10), 1592 => to_unsigned(585, 10), 1593 => to_unsigned(692, 10), 1594 => to_unsigned(670, 10), 1595 => to_unsigned(299, 10), 1596 => to_unsigned(482, 10), 1597 => to_unsigned(155, 10), 1598 => to_unsigned(255, 10), 1599 => to_unsigned(775, 10), 1600 => to_unsigned(409, 10), 1601 => to_unsigned(976, 10), 1602 => to_unsigned(692, 10), 1603 => to_unsigned(820, 10), 1604 => to_unsigned(364, 10), 1605 => to_unsigned(962, 10), 1606 => to_unsigned(438, 10), 1607 => to_unsigned(414, 10), 1608 => to_unsigned(772, 10), 1609 => to_unsigned(584, 10), 1610 => to_unsigned(880, 10), 1611 => to_unsigned(788, 10), 1612 => to_unsigned(431, 10), 1613 => to_unsigned(225, 10), 1614 => to_unsigned(701, 10), 1615 => to_unsigned(838, 10), 1616 => to_unsigned(503, 10), 1617 => to_unsigned(797, 10), 1618 => to_unsigned(454, 10), 1619 => to_unsigned(249, 10), 1620 => to_unsigned(676, 10), 1621 => to_unsigned(474, 10), 1622 => to_unsigned(545, 10), 1623 => to_unsigned(468, 10), 1624 => to_unsigned(975, 10), 1625 => to_unsigned(824, 10), 1626 => to_unsigned(523, 10), 1627 => to_unsigned(527, 10), 1628 => to_unsigned(633, 10), 1629 => to_unsigned(746, 10), 1630 => to_unsigned(405, 10), 1631 => to_unsigned(91, 10), 1632 => to_unsigned(43, 10), 1633 => to_unsigned(850, 10), 1634 => to_unsigned(650, 10), 1635 => to_unsigned(268, 10), 1636 => to_unsigned(688, 10), 1637 => to_unsigned(758, 10), 1638 => to_unsigned(374, 10), 1639 => to_unsigned(626, 10), 1640 => to_unsigned(2, 10), 1641 => to_unsigned(459, 10), 1642 => to_unsigned(390, 10), 1643 => to_unsigned(865, 10), 1644 => to_unsigned(215, 10), 1645 => to_unsigned(885, 10), 1646 => to_unsigned(233, 10), 1647 => to_unsigned(222, 10), 1648 => to_unsigned(189, 10), 1649 => to_unsigned(703, 10), 1650 => to_unsigned(666, 10), 1651 => to_unsigned(248, 10), 1652 => to_unsigned(42, 10), 1653 => to_unsigned(728, 10), 1654 => to_unsigned(899, 10), 1655 => to_unsigned(84, 10), 1656 => to_unsigned(343, 10), 1657 => to_unsigned(383, 10), 1658 => to_unsigned(843, 10), 1659 => to_unsigned(516, 10), 1660 => to_unsigned(949, 10), 1661 => to_unsigned(683, 10), 1662 => to_unsigned(754, 10), 1663 => to_unsigned(326, 10), 1664 => to_unsigned(221, 10), 1665 => to_unsigned(74, 10), 1666 => to_unsigned(88, 10), 1667 => to_unsigned(1023, 10), 1668 => to_unsigned(186, 10), 1669 => to_unsigned(213, 10), 1670 => to_unsigned(713, 10), 1671 => to_unsigned(934, 10), 1672 => to_unsigned(330, 10), 1673 => to_unsigned(201, 10), 1674 => to_unsigned(293, 10), 1675 => to_unsigned(587, 10), 1676 => to_unsigned(531, 10), 1677 => to_unsigned(484, 10), 1678 => to_unsigned(815, 10), 1679 => to_unsigned(821, 10), 1680 => to_unsigned(572, 10), 1681 => to_unsigned(242, 10), 1682 => to_unsigned(430, 10), 1683 => to_unsigned(506, 10), 1684 => to_unsigned(157, 10), 1685 => to_unsigned(28, 10), 1686 => to_unsigned(935, 10), 1687 => to_unsigned(710, 10), 1688 => to_unsigned(386, 10), 1689 => to_unsigned(521, 10), 1690 => to_unsigned(227, 10), 1691 => to_unsigned(8, 10), 1692 => to_unsigned(520, 10), 1693 => to_unsigned(259, 10), 1694 => to_unsigned(208, 10), 1695 => to_unsigned(456, 10), 1696 => to_unsigned(201, 10), 1697 => to_unsigned(27, 10), 1698 => to_unsigned(758, 10), 1699 => to_unsigned(279, 10), 1700 => to_unsigned(765, 10), 1701 => to_unsigned(244, 10), 1702 => to_unsigned(283, 10), 1703 => to_unsigned(58, 10), 1704 => to_unsigned(794, 10), 1705 => to_unsigned(155, 10), 1706 => to_unsigned(64, 10), 1707 => to_unsigned(833, 10), 1708 => to_unsigned(918, 10), 1709 => to_unsigned(799, 10), 1710 => to_unsigned(658, 10), 1711 => to_unsigned(884, 10), 1712 => to_unsigned(537, 10), 1713 => to_unsigned(580, 10), 1714 => to_unsigned(432, 10), 1715 => to_unsigned(588, 10), 1716 => to_unsigned(764, 10), 1717 => to_unsigned(946, 10), 1718 => to_unsigned(640, 10), 1719 => to_unsigned(428, 10), 1720 => to_unsigned(633, 10), 1721 => to_unsigned(979, 10), 1722 => to_unsigned(629, 10), 1723 => to_unsigned(891, 10), 1724 => to_unsigned(1018, 10), 1725 => to_unsigned(54, 10), 1726 => to_unsigned(415, 10), 1727 => to_unsigned(772, 10), 1728 => to_unsigned(103, 10), 1729 => to_unsigned(105, 10), 1730 => to_unsigned(729, 10), 1731 => to_unsigned(557, 10), 1732 => to_unsigned(348, 10), 1733 => to_unsigned(789, 10), 1734 => to_unsigned(678, 10), 1735 => to_unsigned(919, 10), 1736 => to_unsigned(439, 10), 1737 => to_unsigned(286, 10), 1738 => to_unsigned(740, 10), 1739 => to_unsigned(736, 10), 1740 => to_unsigned(427, 10), 1741 => to_unsigned(996, 10), 1742 => to_unsigned(143, 10), 1743 => to_unsigned(540, 10), 1744 => to_unsigned(247, 10), 1745 => to_unsigned(649, 10), 1746 => to_unsigned(934, 10), 1747 => to_unsigned(493, 10), 1748 => to_unsigned(589, 10), 1749 => to_unsigned(794, 10), 1750 => to_unsigned(125, 10), 1751 => to_unsigned(451, 10), 1752 => to_unsigned(363, 10), 1753 => to_unsigned(807, 10), 1754 => to_unsigned(611, 10), 1755 => to_unsigned(24, 10), 1756 => to_unsigned(483, 10), 1757 => to_unsigned(281, 10), 1758 => to_unsigned(356, 10), 1759 => to_unsigned(841, 10), 1760 => to_unsigned(280, 10), 1761 => to_unsigned(472, 10), 1762 => to_unsigned(273, 10), 1763 => to_unsigned(802, 10), 1764 => to_unsigned(831, 10), 1765 => to_unsigned(826, 10), 1766 => to_unsigned(533, 10), 1767 => to_unsigned(597, 10), 1768 => to_unsigned(248, 10), 1769 => to_unsigned(279, 10), 1770 => to_unsigned(109, 10), 1771 => to_unsigned(330, 10), 1772 => to_unsigned(655, 10), 1773 => to_unsigned(741, 10), 1774 => to_unsigned(421, 10), 1775 => to_unsigned(94, 10), 1776 => to_unsigned(646, 10), 1777 => to_unsigned(478, 10), 1778 => to_unsigned(742, 10), 1779 => to_unsigned(1021, 10), 1780 => to_unsigned(929, 10), 1781 => to_unsigned(840, 10), 1782 => to_unsigned(759, 10), 1783 => to_unsigned(459, 10), 1784 => to_unsigned(671, 10), 1785 => to_unsigned(362, 10), 1786 => to_unsigned(245, 10), 1787 => to_unsigned(29, 10), 1788 => to_unsigned(126, 10), 1789 => to_unsigned(474, 10), 1790 => to_unsigned(677, 10), 1791 => to_unsigned(265, 10), 1792 => to_unsigned(991, 10), 1793 => to_unsigned(127, 10), 1794 => to_unsigned(693, 10), 1795 => to_unsigned(593, 10), 1796 => to_unsigned(985, 10), 1797 => to_unsigned(18, 10), 1798 => to_unsigned(482, 10), 1799 => to_unsigned(840, 10), 1800 => to_unsigned(970, 10), 1801 => to_unsigned(640, 10), 1802 => to_unsigned(161, 10), 1803 => to_unsigned(93, 10), 1804 => to_unsigned(971, 10), 1805 => to_unsigned(866, 10), 1806 => to_unsigned(1022, 10), 1807 => to_unsigned(977, 10), 1808 => to_unsigned(331, 10), 1809 => to_unsigned(975, 10), 1810 => to_unsigned(485, 10), 1811 => to_unsigned(503, 10), 1812 => to_unsigned(337, 10), 1813 => to_unsigned(837, 10), 1814 => to_unsigned(267, 10), 1815 => to_unsigned(770, 10), 1816 => to_unsigned(889, 10), 1817 => to_unsigned(922, 10), 1818 => to_unsigned(936, 10), 1819 => to_unsigned(25, 10), 1820 => to_unsigned(587, 10), 1821 => to_unsigned(359, 10), 1822 => to_unsigned(121, 10), 1823 => to_unsigned(396, 10), 1824 => to_unsigned(726, 10), 1825 => to_unsigned(340, 10), 1826 => to_unsigned(416, 10), 1827 => to_unsigned(57, 10), 1828 => to_unsigned(566, 10), 1829 => to_unsigned(1, 10), 1830 => to_unsigned(565, 10), 1831 => to_unsigned(787, 10), 1832 => to_unsigned(590, 10), 1833 => to_unsigned(765, 10), 1834 => to_unsigned(43, 10), 1835 => to_unsigned(83, 10), 1836 => to_unsigned(201, 10), 1837 => to_unsigned(945, 10), 1838 => to_unsigned(932, 10), 1839 => to_unsigned(34, 10), 1840 => to_unsigned(390, 10), 1841 => to_unsigned(763, 10), 1842 => to_unsigned(890, 10), 1843 => to_unsigned(21, 10), 1844 => to_unsigned(933, 10), 1845 => to_unsigned(978, 10), 1846 => to_unsigned(848, 10), 1847 => to_unsigned(198, 10), 1848 => to_unsigned(463, 10), 1849 => to_unsigned(111, 10), 1850 => to_unsigned(934, 10), 1851 => to_unsigned(617, 10), 1852 => to_unsigned(77, 10), 1853 => to_unsigned(953, 10), 1854 => to_unsigned(788, 10), 1855 => to_unsigned(769, 10), 1856 => to_unsigned(432, 10), 1857 => to_unsigned(430, 10), 1858 => to_unsigned(309, 10), 1859 => to_unsigned(542, 10), 1860 => to_unsigned(289, 10), 1861 => to_unsigned(839, 10), 1862 => to_unsigned(179, 10), 1863 => to_unsigned(307, 10), 1864 => to_unsigned(302, 10), 1865 => to_unsigned(628, 10), 1866 => to_unsigned(350, 10), 1867 => to_unsigned(853, 10), 1868 => to_unsigned(558, 10), 1869 => to_unsigned(963, 10), 1870 => to_unsigned(232, 10), 1871 => to_unsigned(665, 10), 1872 => to_unsigned(1018, 10), 1873 => to_unsigned(753, 10), 1874 => to_unsigned(1000, 10), 1875 => to_unsigned(809, 10), 1876 => to_unsigned(342, 10), 1877 => to_unsigned(705, 10), 1878 => to_unsigned(611, 10), 1879 => to_unsigned(576, 10), 1880 => to_unsigned(35, 10), 1881 => to_unsigned(588, 10), 1882 => to_unsigned(278, 10), 1883 => to_unsigned(829, 10), 1884 => to_unsigned(445, 10), 1885 => to_unsigned(916, 10), 1886 => to_unsigned(1000, 10), 1887 => to_unsigned(103, 10), 1888 => to_unsigned(558, 10), 1889 => to_unsigned(560, 10), 1890 => to_unsigned(92, 10), 1891 => to_unsigned(77, 10), 1892 => to_unsigned(901, 10), 1893 => to_unsigned(18, 10), 1894 => to_unsigned(269, 10), 1895 => to_unsigned(326, 10), 1896 => to_unsigned(94, 10), 1897 => to_unsigned(325, 10), 1898 => to_unsigned(1004, 10), 1899 => to_unsigned(342, 10), 1900 => to_unsigned(929, 10), 1901 => to_unsigned(836, 10), 1902 => to_unsigned(782, 10), 1903 => to_unsigned(190, 10), 1904 => to_unsigned(686, 10), 1905 => to_unsigned(677, 10), 1906 => to_unsigned(460, 10), 1907 => to_unsigned(43, 10), 1908 => to_unsigned(454, 10), 1909 => to_unsigned(552, 10), 1910 => to_unsigned(411, 10), 1911 => to_unsigned(299, 10), 1912 => to_unsigned(899, 10), 1913 => to_unsigned(17, 10), 1914 => to_unsigned(47, 10), 1915 => to_unsigned(944, 10), 1916 => to_unsigned(204, 10), 1917 => to_unsigned(431, 10), 1918 => to_unsigned(799, 10), 1919 => to_unsigned(271, 10), 1920 => to_unsigned(465, 10), 1921 => to_unsigned(267, 10), 1922 => to_unsigned(809, 10), 1923 => to_unsigned(513, 10), 1924 => to_unsigned(790, 10), 1925 => to_unsigned(102, 10), 1926 => to_unsigned(55, 10), 1927 => to_unsigned(773, 10), 1928 => to_unsigned(875, 10), 1929 => to_unsigned(963, 10), 1930 => to_unsigned(273, 10), 1931 => to_unsigned(817, 10), 1932 => to_unsigned(368, 10), 1933 => to_unsigned(792, 10), 1934 => to_unsigned(187, 10), 1935 => to_unsigned(691, 10), 1936 => to_unsigned(593, 10), 1937 => to_unsigned(85, 10), 1938 => to_unsigned(314, 10), 1939 => to_unsigned(256, 10), 1940 => to_unsigned(594, 10), 1941 => to_unsigned(977, 10), 1942 => to_unsigned(540, 10), 1943 => to_unsigned(15, 10), 1944 => to_unsigned(612, 10), 1945 => to_unsigned(484, 10), 1946 => to_unsigned(300, 10), 1947 => to_unsigned(351, 10), 1948 => to_unsigned(705, 10), 1949 => to_unsigned(270, 10), 1950 => to_unsigned(32, 10), 1951 => to_unsigned(48, 10), 1952 => to_unsigned(386, 10), 1953 => to_unsigned(107, 10), 1954 => to_unsigned(916, 10), 1955 => to_unsigned(648, 10), 1956 => to_unsigned(913, 10), 1957 => to_unsigned(54, 10), 1958 => to_unsigned(83, 10), 1959 => to_unsigned(626, 10), 1960 => to_unsigned(674, 10), 1961 => to_unsigned(584, 10), 1962 => to_unsigned(599, 10), 1963 => to_unsigned(86, 10), 1964 => to_unsigned(89, 10), 1965 => to_unsigned(361, 10), 1966 => to_unsigned(831, 10), 1967 => to_unsigned(717, 10), 1968 => to_unsigned(376, 10), 1969 => to_unsigned(943, 10), 1970 => to_unsigned(270, 10), 1971 => to_unsigned(696, 10), 1972 => to_unsigned(680, 10), 1973 => to_unsigned(694, 10), 1974 => to_unsigned(592, 10), 1975 => to_unsigned(806, 10), 1976 => to_unsigned(25, 10), 1977 => to_unsigned(441, 10), 1978 => to_unsigned(216, 10), 1979 => to_unsigned(337, 10), 1980 => to_unsigned(63, 10), 1981 => to_unsigned(114, 10), 1982 => to_unsigned(165, 10), 1983 => to_unsigned(734, 10), 1984 => to_unsigned(961, 10), 1985 => to_unsigned(777, 10), 1986 => to_unsigned(621, 10), 1987 => to_unsigned(827, 10), 1988 => to_unsigned(750, 10), 1989 => to_unsigned(385, 10), 1990 => to_unsigned(280, 10), 1991 => to_unsigned(421, 10), 1992 => to_unsigned(888, 10), 1993 => to_unsigned(536, 10), 1994 => to_unsigned(60, 10), 1995 => to_unsigned(977, 10), 1996 => to_unsigned(231, 10), 1997 => to_unsigned(741, 10), 1998 => to_unsigned(454, 10), 1999 => to_unsigned(235, 10), 2000 => to_unsigned(462, 10), 2001 => to_unsigned(216, 10), 2002 => to_unsigned(488, 10), 2003 => to_unsigned(983, 10), 2004 => to_unsigned(549, 10), 2005 => to_unsigned(540, 10), 2006 => to_unsigned(130, 10), 2007 => to_unsigned(724, 10), 2008 => to_unsigned(440, 10), 2009 => to_unsigned(463, 10), 2010 => to_unsigned(797, 10), 2011 => to_unsigned(719, 10), 2012 => to_unsigned(8, 10), 2013 => to_unsigned(1001, 10), 2014 => to_unsigned(274, 10), 2015 => to_unsigned(863, 10), 2016 => to_unsigned(712, 10), 2017 => to_unsigned(699, 10), 2018 => to_unsigned(222, 10), 2019 => to_unsigned(687, 10), 2020 => to_unsigned(127, 10), 2021 => to_unsigned(997, 10), 2022 => to_unsigned(742, 10), 2023 => to_unsigned(592, 10), 2024 => to_unsigned(389, 10), 2025 => to_unsigned(172, 10), 2026 => to_unsigned(598, 10), 2027 => to_unsigned(501, 10), 2028 => to_unsigned(548, 10), 2029 => to_unsigned(814, 10), 2030 => to_unsigned(1014, 10), 2031 => to_unsigned(781, 10), 2032 => to_unsigned(113, 10), 2033 => to_unsigned(143, 10), 2034 => to_unsigned(368, 10), 2035 => to_unsigned(456, 10), 2036 => to_unsigned(31, 10), 2037 => to_unsigned(985, 10), 2038 => to_unsigned(45, 10), 2039 => to_unsigned(21, 10), 2040 => to_unsigned(592, 10), 2041 => to_unsigned(162, 10), 2042 => to_unsigned(649, 10), 2043 => to_unsigned(393, 10), 2044 => to_unsigned(349, 10), 2045 => to_unsigned(798, 10), 2046 => to_unsigned(266, 10), 2047 => to_unsigned(998, 10)),
            7 => (0 => to_unsigned(931, 10), 1 => to_unsigned(376, 10), 2 => to_unsigned(952, 10), 3 => to_unsigned(558, 10), 4 => to_unsigned(94, 10), 5 => to_unsigned(155, 10), 6 => to_unsigned(437, 10), 7 => to_unsigned(580, 10), 8 => to_unsigned(209, 10), 9 => to_unsigned(697, 10), 10 => to_unsigned(301, 10), 11 => to_unsigned(884, 10), 12 => to_unsigned(266, 10), 13 => to_unsigned(684, 10), 14 => to_unsigned(151, 10), 15 => to_unsigned(490, 10), 16 => to_unsigned(81, 10), 17 => to_unsigned(807, 10), 18 => to_unsigned(760, 10), 19 => to_unsigned(189, 10), 20 => to_unsigned(438, 10), 21 => to_unsigned(359, 10), 22 => to_unsigned(922, 10), 23 => to_unsigned(117, 10), 24 => to_unsigned(697, 10), 25 => to_unsigned(857, 10), 26 => to_unsigned(946, 10), 27 => to_unsigned(102, 10), 28 => to_unsigned(219, 10), 29 => to_unsigned(762, 10), 30 => to_unsigned(23, 10), 31 => to_unsigned(545, 10), 32 => to_unsigned(798, 10), 33 => to_unsigned(808, 10), 34 => to_unsigned(420, 10), 35 => to_unsigned(987, 10), 36 => to_unsigned(377, 10), 37 => to_unsigned(336, 10), 38 => to_unsigned(211, 10), 39 => to_unsigned(494, 10), 40 => to_unsigned(376, 10), 41 => to_unsigned(382, 10), 42 => to_unsigned(565, 10), 43 => to_unsigned(153, 10), 44 => to_unsigned(1023, 10), 45 => to_unsigned(392, 10), 46 => to_unsigned(29, 10), 47 => to_unsigned(825, 10), 48 => to_unsigned(335, 10), 49 => to_unsigned(623, 10), 50 => to_unsigned(64, 10), 51 => to_unsigned(760, 10), 52 => to_unsigned(691, 10), 53 => to_unsigned(444, 10), 54 => to_unsigned(245, 10), 55 => to_unsigned(55, 10), 56 => to_unsigned(139, 10), 57 => to_unsigned(498, 10), 58 => to_unsigned(342, 10), 59 => to_unsigned(226, 10), 60 => to_unsigned(473, 10), 61 => to_unsigned(936, 10), 62 => to_unsigned(371, 10), 63 => to_unsigned(224, 10), 64 => to_unsigned(950, 10), 65 => to_unsigned(733, 10), 66 => to_unsigned(196, 10), 67 => to_unsigned(437, 10), 68 => to_unsigned(167, 10), 69 => to_unsigned(56, 10), 70 => to_unsigned(110, 10), 71 => to_unsigned(329, 10), 72 => to_unsigned(323, 10), 73 => to_unsigned(202, 10), 74 => to_unsigned(895, 10), 75 => to_unsigned(150, 10), 76 => to_unsigned(284, 10), 77 => to_unsigned(344, 10), 78 => to_unsigned(1021, 10), 79 => to_unsigned(854, 10), 80 => to_unsigned(516, 10), 81 => to_unsigned(852, 10), 82 => to_unsigned(596, 10), 83 => to_unsigned(702, 10), 84 => to_unsigned(93, 10), 85 => to_unsigned(1004, 10), 86 => to_unsigned(1011, 10), 87 => to_unsigned(111, 10), 88 => to_unsigned(436, 10), 89 => to_unsigned(142, 10), 90 => to_unsigned(452, 10), 91 => to_unsigned(87, 10), 92 => to_unsigned(750, 10), 93 => to_unsigned(515, 10), 94 => to_unsigned(441, 10), 95 => to_unsigned(946, 10), 96 => to_unsigned(983, 10), 97 => to_unsigned(646, 10), 98 => to_unsigned(586, 10), 99 => to_unsigned(884, 10), 100 => to_unsigned(462, 10), 101 => to_unsigned(780, 10), 102 => to_unsigned(146, 10), 103 => to_unsigned(447, 10), 104 => to_unsigned(88, 10), 105 => to_unsigned(840, 10), 106 => to_unsigned(284, 10), 107 => to_unsigned(634, 10), 108 => to_unsigned(406, 10), 109 => to_unsigned(184, 10), 110 => to_unsigned(264, 10), 111 => to_unsigned(210, 10), 112 => to_unsigned(760, 10), 113 => to_unsigned(653, 10), 114 => to_unsigned(511, 10), 115 => to_unsigned(242, 10), 116 => to_unsigned(923, 10), 117 => to_unsigned(948, 10), 118 => to_unsigned(690, 10), 119 => to_unsigned(974, 10), 120 => to_unsigned(783, 10), 121 => to_unsigned(905, 10), 122 => to_unsigned(237, 10), 123 => to_unsigned(178, 10), 124 => to_unsigned(95, 10), 125 => to_unsigned(395, 10), 126 => to_unsigned(221, 10), 127 => to_unsigned(841, 10), 128 => to_unsigned(648, 10), 129 => to_unsigned(431, 10), 130 => to_unsigned(641, 10), 131 => to_unsigned(281, 10), 132 => to_unsigned(717, 10), 133 => to_unsigned(822, 10), 134 => to_unsigned(576, 10), 135 => to_unsigned(377, 10), 136 => to_unsigned(864, 10), 137 => to_unsigned(585, 10), 138 => to_unsigned(992, 10), 139 => to_unsigned(178, 10), 140 => to_unsigned(315, 10), 141 => to_unsigned(51, 10), 142 => to_unsigned(217, 10), 143 => to_unsigned(979, 10), 144 => to_unsigned(318, 10), 145 => to_unsigned(227, 10), 146 => to_unsigned(249, 10), 147 => to_unsigned(960, 10), 148 => to_unsigned(484, 10), 149 => to_unsigned(370, 10), 150 => to_unsigned(291, 10), 151 => to_unsigned(89, 10), 152 => to_unsigned(424, 10), 153 => to_unsigned(46, 10), 154 => to_unsigned(702, 10), 155 => to_unsigned(29, 10), 156 => to_unsigned(313, 10), 157 => to_unsigned(230, 10), 158 => to_unsigned(356, 10), 159 => to_unsigned(55, 10), 160 => to_unsigned(483, 10), 161 => to_unsigned(733, 10), 162 => to_unsigned(148, 10), 163 => to_unsigned(54, 10), 164 => to_unsigned(376, 10), 165 => to_unsigned(722, 10), 166 => to_unsigned(891, 10), 167 => to_unsigned(320, 10), 168 => to_unsigned(257, 10), 169 => to_unsigned(662, 10), 170 => to_unsigned(233, 10), 171 => to_unsigned(687, 10), 172 => to_unsigned(786, 10), 173 => to_unsigned(114, 10), 174 => to_unsigned(763, 10), 175 => to_unsigned(8, 10), 176 => to_unsigned(175, 10), 177 => to_unsigned(624, 10), 178 => to_unsigned(533, 10), 179 => to_unsigned(942, 10), 180 => to_unsigned(466, 10), 181 => to_unsigned(1021, 10), 182 => to_unsigned(204, 10), 183 => to_unsigned(399, 10), 184 => to_unsigned(733, 10), 185 => to_unsigned(762, 10), 186 => to_unsigned(719, 10), 187 => to_unsigned(434, 10), 188 => to_unsigned(135, 10), 189 => to_unsigned(151, 10), 190 => to_unsigned(351, 10), 191 => to_unsigned(494, 10), 192 => to_unsigned(21, 10), 193 => to_unsigned(103, 10), 194 => to_unsigned(142, 10), 195 => to_unsigned(317, 10), 196 => to_unsigned(921, 10), 197 => to_unsigned(850, 10), 198 => to_unsigned(836, 10), 199 => to_unsigned(495, 10), 200 => to_unsigned(735, 10), 201 => to_unsigned(609, 10), 202 => to_unsigned(191, 10), 203 => to_unsigned(326, 10), 204 => to_unsigned(289, 10), 205 => to_unsigned(406, 10), 206 => to_unsigned(764, 10), 207 => to_unsigned(876, 10), 208 => to_unsigned(201, 10), 209 => to_unsigned(791, 10), 210 => to_unsigned(855, 10), 211 => to_unsigned(95, 10), 212 => to_unsigned(999, 10), 213 => to_unsigned(495, 10), 214 => to_unsigned(14, 10), 215 => to_unsigned(425, 10), 216 => to_unsigned(393, 10), 217 => to_unsigned(228, 10), 218 => to_unsigned(24, 10), 219 => to_unsigned(883, 10), 220 => to_unsigned(835, 10), 221 => to_unsigned(1013, 10), 222 => to_unsigned(5, 10), 223 => to_unsigned(831, 10), 224 => to_unsigned(586, 10), 225 => to_unsigned(870, 10), 226 => to_unsigned(412, 10), 227 => to_unsigned(607, 10), 228 => to_unsigned(22, 10), 229 => to_unsigned(617, 10), 230 => to_unsigned(502, 10), 231 => to_unsigned(200, 10), 232 => to_unsigned(254, 10), 233 => to_unsigned(458, 10), 234 => to_unsigned(341, 10), 235 => to_unsigned(670, 10), 236 => to_unsigned(978, 10), 237 => to_unsigned(57, 10), 238 => to_unsigned(990, 10), 239 => to_unsigned(604, 10), 240 => to_unsigned(747, 10), 241 => to_unsigned(543, 10), 242 => to_unsigned(478, 10), 243 => to_unsigned(672, 10), 244 => to_unsigned(553, 10), 245 => to_unsigned(120, 10), 246 => to_unsigned(796, 10), 247 => to_unsigned(580, 10), 248 => to_unsigned(490, 10), 249 => to_unsigned(833, 10), 250 => to_unsigned(255, 10), 251 => to_unsigned(354, 10), 252 => to_unsigned(482, 10), 253 => to_unsigned(918, 10), 254 => to_unsigned(240, 10), 255 => to_unsigned(237, 10), 256 => to_unsigned(454, 10), 257 => to_unsigned(873, 10), 258 => to_unsigned(601, 10), 259 => to_unsigned(364, 10), 260 => to_unsigned(467, 10), 261 => to_unsigned(1022, 10), 262 => to_unsigned(905, 10), 263 => to_unsigned(994, 10), 264 => to_unsigned(86, 10), 265 => to_unsigned(870, 10), 266 => to_unsigned(681, 10), 267 => to_unsigned(315, 10), 268 => to_unsigned(440, 10), 269 => to_unsigned(181, 10), 270 => to_unsigned(156, 10), 271 => to_unsigned(919, 10), 272 => to_unsigned(260, 10), 273 => to_unsigned(381, 10), 274 => to_unsigned(87, 10), 275 => to_unsigned(103, 10), 276 => to_unsigned(529, 10), 277 => to_unsigned(62, 10), 278 => to_unsigned(136, 10), 279 => to_unsigned(713, 10), 280 => to_unsigned(756, 10), 281 => to_unsigned(504, 10), 282 => to_unsigned(705, 10), 283 => to_unsigned(892, 10), 284 => to_unsigned(479, 10), 285 => to_unsigned(399, 10), 286 => to_unsigned(465, 10), 287 => to_unsigned(325, 10), 288 => to_unsigned(647, 10), 289 => to_unsigned(109, 10), 290 => to_unsigned(706, 10), 291 => to_unsigned(155, 10), 292 => to_unsigned(866, 10), 293 => to_unsigned(198, 10), 294 => to_unsigned(664, 10), 295 => to_unsigned(1010, 10), 296 => to_unsigned(356, 10), 297 => to_unsigned(365, 10), 298 => to_unsigned(524, 10), 299 => to_unsigned(949, 10), 300 => to_unsigned(525, 10), 301 => to_unsigned(349, 10), 302 => to_unsigned(1005, 10), 303 => to_unsigned(413, 10), 304 => to_unsigned(977, 10), 305 => to_unsigned(330, 10), 306 => to_unsigned(680, 10), 307 => to_unsigned(283, 10), 308 => to_unsigned(30, 10), 309 => to_unsigned(610, 10), 310 => to_unsigned(152, 10), 311 => to_unsigned(450, 10), 312 => to_unsigned(826, 10), 313 => to_unsigned(393, 10), 314 => to_unsigned(575, 10), 315 => to_unsigned(997, 10), 316 => to_unsigned(262, 10), 317 => to_unsigned(364, 10), 318 => to_unsigned(773, 10), 319 => to_unsigned(939, 10), 320 => to_unsigned(371, 10), 321 => to_unsigned(102, 10), 322 => to_unsigned(774, 10), 323 => to_unsigned(631, 10), 324 => to_unsigned(314, 10), 325 => to_unsigned(545, 10), 326 => to_unsigned(266, 10), 327 => to_unsigned(398, 10), 328 => to_unsigned(242, 10), 329 => to_unsigned(600, 10), 330 => to_unsigned(905, 10), 331 => to_unsigned(278, 10), 332 => to_unsigned(936, 10), 333 => to_unsigned(642, 10), 334 => to_unsigned(243, 10), 335 => to_unsigned(722, 10), 336 => to_unsigned(291, 10), 337 => to_unsigned(936, 10), 338 => to_unsigned(1018, 10), 339 => to_unsigned(842, 10), 340 => to_unsigned(672, 10), 341 => to_unsigned(947, 10), 342 => to_unsigned(662, 10), 343 => to_unsigned(149, 10), 344 => to_unsigned(312, 10), 345 => to_unsigned(682, 10), 346 => to_unsigned(73, 10), 347 => to_unsigned(882, 10), 348 => to_unsigned(976, 10), 349 => to_unsigned(746, 10), 350 => to_unsigned(683, 10), 351 => to_unsigned(855, 10), 352 => to_unsigned(885, 10), 353 => to_unsigned(475, 10), 354 => to_unsigned(822, 10), 355 => to_unsigned(762, 10), 356 => to_unsigned(727, 10), 357 => to_unsigned(382, 10), 358 => to_unsigned(109, 10), 359 => to_unsigned(697, 10), 360 => to_unsigned(334, 10), 361 => to_unsigned(174, 10), 362 => to_unsigned(800, 10), 363 => to_unsigned(232, 10), 364 => to_unsigned(905, 10), 365 => to_unsigned(480, 10), 366 => to_unsigned(790, 10), 367 => to_unsigned(55, 10), 368 => to_unsigned(356, 10), 369 => to_unsigned(493, 10), 370 => to_unsigned(629, 10), 371 => to_unsigned(431, 10), 372 => to_unsigned(798, 10), 373 => to_unsigned(509, 10), 374 => to_unsigned(8, 10), 375 => to_unsigned(481, 10), 376 => to_unsigned(622, 10), 377 => to_unsigned(12, 10), 378 => to_unsigned(737, 10), 379 => to_unsigned(216, 10), 380 => to_unsigned(680, 10), 381 => to_unsigned(36, 10), 382 => to_unsigned(803, 10), 383 => to_unsigned(111, 10), 384 => to_unsigned(134, 10), 385 => to_unsigned(431, 10), 386 => to_unsigned(281, 10), 387 => to_unsigned(238, 10), 388 => to_unsigned(434, 10), 389 => to_unsigned(261, 10), 390 => to_unsigned(167, 10), 391 => to_unsigned(425, 10), 392 => to_unsigned(572, 10), 393 => to_unsigned(633, 10), 394 => to_unsigned(191, 10), 395 => to_unsigned(171, 10), 396 => to_unsigned(921, 10), 397 => to_unsigned(433, 10), 398 => to_unsigned(97, 10), 399 => to_unsigned(58, 10), 400 => to_unsigned(759, 10), 401 => to_unsigned(589, 10), 402 => to_unsigned(883, 10), 403 => to_unsigned(180, 10), 404 => to_unsigned(557, 10), 405 => to_unsigned(7, 10), 406 => to_unsigned(207, 10), 407 => to_unsigned(403, 10), 408 => to_unsigned(249, 10), 409 => to_unsigned(508, 10), 410 => to_unsigned(307, 10), 411 => to_unsigned(691, 10), 412 => to_unsigned(674, 10), 413 => to_unsigned(863, 10), 414 => to_unsigned(666, 10), 415 => to_unsigned(747, 10), 416 => to_unsigned(181, 10), 417 => to_unsigned(836, 10), 418 => to_unsigned(825, 10), 419 => to_unsigned(857, 10), 420 => to_unsigned(370, 10), 421 => to_unsigned(217, 10), 422 => to_unsigned(916, 10), 423 => to_unsigned(960, 10), 424 => to_unsigned(439, 10), 425 => to_unsigned(10, 10), 426 => to_unsigned(158, 10), 427 => to_unsigned(753, 10), 428 => to_unsigned(715, 10), 429 => to_unsigned(888, 10), 430 => to_unsigned(284, 10), 431 => to_unsigned(908, 10), 432 => to_unsigned(373, 10), 433 => to_unsigned(818, 10), 434 => to_unsigned(776, 10), 435 => to_unsigned(517, 10), 436 => to_unsigned(581, 10), 437 => to_unsigned(549, 10), 438 => to_unsigned(497, 10), 439 => to_unsigned(458, 10), 440 => to_unsigned(815, 10), 441 => to_unsigned(320, 10), 442 => to_unsigned(756, 10), 443 => to_unsigned(111, 10), 444 => to_unsigned(403, 10), 445 => to_unsigned(756, 10), 446 => to_unsigned(947, 10), 447 => to_unsigned(26, 10), 448 => to_unsigned(653, 10), 449 => to_unsigned(920, 10), 450 => to_unsigned(618, 10), 451 => to_unsigned(786, 10), 452 => to_unsigned(73, 10), 453 => to_unsigned(316, 10), 454 => to_unsigned(652, 10), 455 => to_unsigned(27, 10), 456 => to_unsigned(205, 10), 457 => to_unsigned(776, 10), 458 => to_unsigned(438, 10), 459 => to_unsigned(375, 10), 460 => to_unsigned(738, 10), 461 => to_unsigned(579, 10), 462 => to_unsigned(6, 10), 463 => to_unsigned(206, 10), 464 => to_unsigned(337, 10), 465 => to_unsigned(585, 10), 466 => to_unsigned(785, 10), 467 => to_unsigned(724, 10), 468 => to_unsigned(1015, 10), 469 => to_unsigned(873, 10), 470 => to_unsigned(455, 10), 471 => to_unsigned(14, 10), 472 => to_unsigned(853, 10), 473 => to_unsigned(224, 10), 474 => to_unsigned(994, 10), 475 => to_unsigned(305, 10), 476 => to_unsigned(882, 10), 477 => to_unsigned(131, 10), 478 => to_unsigned(228, 10), 479 => to_unsigned(605, 10), 480 => to_unsigned(377, 10), 481 => to_unsigned(790, 10), 482 => to_unsigned(527, 10), 483 => to_unsigned(232, 10), 484 => to_unsigned(865, 10), 485 => to_unsigned(101, 10), 486 => to_unsigned(593, 10), 487 => to_unsigned(78, 10), 488 => to_unsigned(387, 10), 489 => to_unsigned(480, 10), 490 => to_unsigned(313, 10), 491 => to_unsigned(400, 10), 492 => to_unsigned(229, 10), 493 => to_unsigned(196, 10), 494 => to_unsigned(376, 10), 495 => to_unsigned(691, 10), 496 => to_unsigned(880, 10), 497 => to_unsigned(479, 10), 498 => to_unsigned(24, 10), 499 => to_unsigned(637, 10), 500 => to_unsigned(268, 10), 501 => to_unsigned(535, 10), 502 => to_unsigned(949, 10), 503 => to_unsigned(397, 10), 504 => to_unsigned(300, 10), 505 => to_unsigned(918, 10), 506 => to_unsigned(695, 10), 507 => to_unsigned(599, 10), 508 => to_unsigned(983, 10), 509 => to_unsigned(854, 10), 510 => to_unsigned(338, 10), 511 => to_unsigned(280, 10), 512 => to_unsigned(1017, 10), 513 => to_unsigned(492, 10), 514 => to_unsigned(588, 10), 515 => to_unsigned(639, 10), 516 => to_unsigned(614, 10), 517 => to_unsigned(366, 10), 518 => to_unsigned(523, 10), 519 => to_unsigned(909, 10), 520 => to_unsigned(256, 10), 521 => to_unsigned(63, 10), 522 => to_unsigned(527, 10), 523 => to_unsigned(574, 10), 524 => to_unsigned(624, 10), 525 => to_unsigned(872, 10), 526 => to_unsigned(507, 10), 527 => to_unsigned(601, 10), 528 => to_unsigned(417, 10), 529 => to_unsigned(361, 10), 530 => to_unsigned(346, 10), 531 => to_unsigned(107, 10), 532 => to_unsigned(395, 10), 533 => to_unsigned(349, 10), 534 => to_unsigned(311, 10), 535 => to_unsigned(202, 10), 536 => to_unsigned(277, 10), 537 => to_unsigned(344, 10), 538 => to_unsigned(461, 10), 539 => to_unsigned(545, 10), 540 => to_unsigned(236, 10), 541 => to_unsigned(521, 10), 542 => to_unsigned(429, 10), 543 => to_unsigned(675, 10), 544 => to_unsigned(354, 10), 545 => to_unsigned(293, 10), 546 => to_unsigned(215, 10), 547 => to_unsigned(106, 10), 548 => to_unsigned(363, 10), 549 => to_unsigned(957, 10), 550 => to_unsigned(629, 10), 551 => to_unsigned(107, 10), 552 => to_unsigned(706, 10), 553 => to_unsigned(294, 10), 554 => to_unsigned(747, 10), 555 => to_unsigned(686, 10), 556 => to_unsigned(385, 10), 557 => to_unsigned(234, 10), 558 => to_unsigned(349, 10), 559 => to_unsigned(570, 10), 560 => to_unsigned(223, 10), 561 => to_unsigned(580, 10), 562 => to_unsigned(430, 10), 563 => to_unsigned(601, 10), 564 => to_unsigned(119, 10), 565 => to_unsigned(621, 10), 566 => to_unsigned(809, 10), 567 => to_unsigned(376, 10), 568 => to_unsigned(775, 10), 569 => to_unsigned(492, 10), 570 => to_unsigned(67, 10), 571 => to_unsigned(122, 10), 572 => to_unsigned(167, 10), 573 => to_unsigned(391, 10), 574 => to_unsigned(788, 10), 575 => to_unsigned(856, 10), 576 => to_unsigned(920, 10), 577 => to_unsigned(289, 10), 578 => to_unsigned(434, 10), 579 => to_unsigned(720, 10), 580 => to_unsigned(635, 10), 581 => to_unsigned(841, 10), 582 => to_unsigned(28, 10), 583 => to_unsigned(846, 10), 584 => to_unsigned(414, 10), 585 => to_unsigned(429, 10), 586 => to_unsigned(714, 10), 587 => to_unsigned(993, 10), 588 => to_unsigned(924, 10), 589 => to_unsigned(959, 10), 590 => to_unsigned(573, 10), 591 => to_unsigned(966, 10), 592 => to_unsigned(168, 10), 593 => to_unsigned(454, 10), 594 => to_unsigned(488, 10), 595 => to_unsigned(469, 10), 596 => to_unsigned(369, 10), 597 => to_unsigned(408, 10), 598 => to_unsigned(49, 10), 599 => to_unsigned(951, 10), 600 => to_unsigned(15, 10), 601 => to_unsigned(139, 10), 602 => to_unsigned(302, 10), 603 => to_unsigned(536, 10), 604 => to_unsigned(594, 10), 605 => to_unsigned(216, 10), 606 => to_unsigned(343, 10), 607 => to_unsigned(610, 10), 608 => to_unsigned(517, 10), 609 => to_unsigned(334, 10), 610 => to_unsigned(1015, 10), 611 => to_unsigned(31, 10), 612 => to_unsigned(111, 10), 613 => to_unsigned(953, 10), 614 => to_unsigned(295, 10), 615 => to_unsigned(383, 10), 616 => to_unsigned(498, 10), 617 => to_unsigned(888, 10), 618 => to_unsigned(742, 10), 619 => to_unsigned(438, 10), 620 => to_unsigned(244, 10), 621 => to_unsigned(593, 10), 622 => to_unsigned(830, 10), 623 => to_unsigned(354, 10), 624 => to_unsigned(424, 10), 625 => to_unsigned(384, 10), 626 => to_unsigned(787, 10), 627 => to_unsigned(614, 10), 628 => to_unsigned(667, 10), 629 => to_unsigned(604, 10), 630 => to_unsigned(133, 10), 631 => to_unsigned(921, 10), 632 => to_unsigned(707, 10), 633 => to_unsigned(262, 10), 634 => to_unsigned(532, 10), 635 => to_unsigned(522, 10), 636 => to_unsigned(769, 10), 637 => to_unsigned(39, 10), 638 => to_unsigned(377, 10), 639 => to_unsigned(533, 10), 640 => to_unsigned(717, 10), 641 => to_unsigned(677, 10), 642 => to_unsigned(267, 10), 643 => to_unsigned(694, 10), 644 => to_unsigned(281, 10), 645 => to_unsigned(1015, 10), 646 => to_unsigned(1014, 10), 647 => to_unsigned(757, 10), 648 => to_unsigned(580, 10), 649 => to_unsigned(745, 10), 650 => to_unsigned(128, 10), 651 => to_unsigned(734, 10), 652 => to_unsigned(244, 10), 653 => to_unsigned(357, 10), 654 => to_unsigned(732, 10), 655 => to_unsigned(9, 10), 656 => to_unsigned(127, 10), 657 => to_unsigned(209, 10), 658 => to_unsigned(702, 10), 659 => to_unsigned(783, 10), 660 => to_unsigned(309, 10), 661 => to_unsigned(307, 10), 662 => to_unsigned(885, 10), 663 => to_unsigned(423, 10), 664 => to_unsigned(592, 10), 665 => to_unsigned(235, 10), 666 => to_unsigned(1017, 10), 667 => to_unsigned(280, 10), 668 => to_unsigned(762, 10), 669 => to_unsigned(678, 10), 670 => to_unsigned(998, 10), 671 => to_unsigned(683, 10), 672 => to_unsigned(17, 10), 673 => to_unsigned(300, 10), 674 => to_unsigned(437, 10), 675 => to_unsigned(532, 10), 676 => to_unsigned(9, 10), 677 => to_unsigned(415, 10), 678 => to_unsigned(135, 10), 679 => to_unsigned(90, 10), 680 => to_unsigned(55, 10), 681 => to_unsigned(342, 10), 682 => to_unsigned(1018, 10), 683 => to_unsigned(1023, 10), 684 => to_unsigned(480, 10), 685 => to_unsigned(772, 10), 686 => to_unsigned(530, 10), 687 => to_unsigned(339, 10), 688 => to_unsigned(557, 10), 689 => to_unsigned(650, 10), 690 => to_unsigned(607, 10), 691 => to_unsigned(134, 10), 692 => to_unsigned(491, 10), 693 => to_unsigned(1020, 10), 694 => to_unsigned(115, 10), 695 => to_unsigned(361, 10), 696 => to_unsigned(774, 10), 697 => to_unsigned(741, 10), 698 => to_unsigned(363, 10), 699 => to_unsigned(357, 10), 700 => to_unsigned(431, 10), 701 => to_unsigned(729, 10), 702 => to_unsigned(914, 10), 703 => to_unsigned(271, 10), 704 => to_unsigned(753, 10), 705 => to_unsigned(220, 10), 706 => to_unsigned(239, 10), 707 => to_unsigned(773, 10), 708 => to_unsigned(647, 10), 709 => to_unsigned(396, 10), 710 => to_unsigned(187, 10), 711 => to_unsigned(996, 10), 712 => to_unsigned(688, 10), 713 => to_unsigned(275, 10), 714 => to_unsigned(103, 10), 715 => to_unsigned(928, 10), 716 => to_unsigned(309, 10), 717 => to_unsigned(580, 10), 718 => to_unsigned(509, 10), 719 => to_unsigned(690, 10), 720 => to_unsigned(554, 10), 721 => to_unsigned(317, 10), 722 => to_unsigned(309, 10), 723 => to_unsigned(967, 10), 724 => to_unsigned(692, 10), 725 => to_unsigned(642, 10), 726 => to_unsigned(746, 10), 727 => to_unsigned(791, 10), 728 => to_unsigned(613, 10), 729 => to_unsigned(140, 10), 730 => to_unsigned(108, 10), 731 => to_unsigned(288, 10), 732 => to_unsigned(617, 10), 733 => to_unsigned(352, 10), 734 => to_unsigned(963, 10), 735 => to_unsigned(21, 10), 736 => to_unsigned(667, 10), 737 => to_unsigned(346, 10), 738 => to_unsigned(829, 10), 739 => to_unsigned(771, 10), 740 => to_unsigned(757, 10), 741 => to_unsigned(118, 10), 742 => to_unsigned(298, 10), 743 => to_unsigned(485, 10), 744 => to_unsigned(462, 10), 745 => to_unsigned(476, 10), 746 => to_unsigned(469, 10), 747 => to_unsigned(821, 10), 748 => to_unsigned(353, 10), 749 => to_unsigned(918, 10), 750 => to_unsigned(556, 10), 751 => to_unsigned(916, 10), 752 => to_unsigned(903, 10), 753 => to_unsigned(284, 10), 754 => to_unsigned(202, 10), 755 => to_unsigned(714, 10), 756 => to_unsigned(81, 10), 757 => to_unsigned(12, 10), 758 => to_unsigned(481, 10), 759 => to_unsigned(926, 10), 760 => to_unsigned(558, 10), 761 => to_unsigned(981, 10), 762 => to_unsigned(242, 10), 763 => to_unsigned(718, 10), 764 => to_unsigned(806, 10), 765 => to_unsigned(1020, 10), 766 => to_unsigned(833, 10), 767 => to_unsigned(445, 10), 768 => to_unsigned(886, 10), 769 => to_unsigned(451, 10), 770 => to_unsigned(294, 10), 771 => to_unsigned(31, 10), 772 => to_unsigned(1020, 10), 773 => to_unsigned(859, 10), 774 => to_unsigned(955, 10), 775 => to_unsigned(150, 10), 776 => to_unsigned(656, 10), 777 => to_unsigned(116, 10), 778 => to_unsigned(245, 10), 779 => to_unsigned(297, 10), 780 => to_unsigned(718, 10), 781 => to_unsigned(369, 10), 782 => to_unsigned(353, 10), 783 => to_unsigned(547, 10), 784 => to_unsigned(972, 10), 785 => to_unsigned(632, 10), 786 => to_unsigned(1010, 10), 787 => to_unsigned(160, 10), 788 => to_unsigned(837, 10), 789 => to_unsigned(421, 10), 790 => to_unsigned(657, 10), 791 => to_unsigned(968, 10), 792 => to_unsigned(126, 10), 793 => to_unsigned(693, 10), 794 => to_unsigned(83, 10), 795 => to_unsigned(825, 10), 796 => to_unsigned(381, 10), 797 => to_unsigned(520, 10), 798 => to_unsigned(653, 10), 799 => to_unsigned(309, 10), 800 => to_unsigned(520, 10), 801 => to_unsigned(354, 10), 802 => to_unsigned(685, 10), 803 => to_unsigned(453, 10), 804 => to_unsigned(401, 10), 805 => to_unsigned(511, 10), 806 => to_unsigned(914, 10), 807 => to_unsigned(65, 10), 808 => to_unsigned(262, 10), 809 => to_unsigned(218, 10), 810 => to_unsigned(376, 10), 811 => to_unsigned(267, 10), 812 => to_unsigned(762, 10), 813 => to_unsigned(169, 10), 814 => to_unsigned(252, 10), 815 => to_unsigned(716, 10), 816 => to_unsigned(994, 10), 817 => to_unsigned(392, 10), 818 => to_unsigned(93, 10), 819 => to_unsigned(253, 10), 820 => to_unsigned(90, 10), 821 => to_unsigned(318, 10), 822 => to_unsigned(787, 10), 823 => to_unsigned(263, 10), 824 => to_unsigned(1017, 10), 825 => to_unsigned(188, 10), 826 => to_unsigned(721, 10), 827 => to_unsigned(591, 10), 828 => to_unsigned(326, 10), 829 => to_unsigned(353, 10), 830 => to_unsigned(290, 10), 831 => to_unsigned(552, 10), 832 => to_unsigned(769, 10), 833 => to_unsigned(78, 10), 834 => to_unsigned(664, 10), 835 => to_unsigned(99, 10), 836 => to_unsigned(453, 10), 837 => to_unsigned(987, 10), 838 => to_unsigned(575, 10), 839 => to_unsigned(541, 10), 840 => to_unsigned(749, 10), 841 => to_unsigned(320, 10), 842 => to_unsigned(583, 10), 843 => to_unsigned(442, 10), 844 => to_unsigned(303, 10), 845 => to_unsigned(66, 10), 846 => to_unsigned(554, 10), 847 => to_unsigned(84, 10), 848 => to_unsigned(350, 10), 849 => to_unsigned(259, 10), 850 => to_unsigned(998, 10), 851 => to_unsigned(79, 10), 852 => to_unsigned(83, 10), 853 => to_unsigned(589, 10), 854 => to_unsigned(929, 10), 855 => to_unsigned(744, 10), 856 => to_unsigned(28, 10), 857 => to_unsigned(957, 10), 858 => to_unsigned(662, 10), 859 => to_unsigned(452, 10), 860 => to_unsigned(982, 10), 861 => to_unsigned(641, 10), 862 => to_unsigned(432, 10), 863 => to_unsigned(238, 10), 864 => to_unsigned(418, 10), 865 => to_unsigned(705, 10), 866 => to_unsigned(850, 10), 867 => to_unsigned(994, 10), 868 => to_unsigned(559, 10), 869 => to_unsigned(501, 10), 870 => to_unsigned(101, 10), 871 => to_unsigned(530, 10), 872 => to_unsigned(674, 10), 873 => to_unsigned(373, 10), 874 => to_unsigned(819, 10), 875 => to_unsigned(37, 10), 876 => to_unsigned(325, 10), 877 => to_unsigned(817, 10), 878 => to_unsigned(453, 10), 879 => to_unsigned(196, 10), 880 => to_unsigned(432, 10), 881 => to_unsigned(555, 10), 882 => to_unsigned(769, 10), 883 => to_unsigned(778, 10), 884 => to_unsigned(787, 10), 885 => to_unsigned(584, 10), 886 => to_unsigned(794, 10), 887 => to_unsigned(817, 10), 888 => to_unsigned(363, 10), 889 => to_unsigned(866, 10), 890 => to_unsigned(195, 10), 891 => to_unsigned(906, 10), 892 => to_unsigned(375, 10), 893 => to_unsigned(898, 10), 894 => to_unsigned(18, 10), 895 => to_unsigned(799, 10), 896 => to_unsigned(547, 10), 897 => to_unsigned(476, 10), 898 => to_unsigned(560, 10), 899 => to_unsigned(813, 10), 900 => to_unsigned(358, 10), 901 => to_unsigned(5, 10), 902 => to_unsigned(69, 10), 903 => to_unsigned(315, 10), 904 => to_unsigned(478, 10), 905 => to_unsigned(241, 10), 906 => to_unsigned(294, 10), 907 => to_unsigned(1005, 10), 908 => to_unsigned(991, 10), 909 => to_unsigned(328, 10), 910 => to_unsigned(944, 10), 911 => to_unsigned(710, 10), 912 => to_unsigned(718, 10), 913 => to_unsigned(386, 10), 914 => to_unsigned(277, 10), 915 => to_unsigned(193, 10), 916 => to_unsigned(147, 10), 917 => to_unsigned(602, 10), 918 => to_unsigned(151, 10), 919 => to_unsigned(877, 10), 920 => to_unsigned(887, 10), 921 => to_unsigned(327, 10), 922 => to_unsigned(537, 10), 923 => to_unsigned(153, 10), 924 => to_unsigned(904, 10), 925 => to_unsigned(825, 10), 926 => to_unsigned(204, 10), 927 => to_unsigned(345, 10), 928 => to_unsigned(223, 10), 929 => to_unsigned(262, 10), 930 => to_unsigned(244, 10), 931 => to_unsigned(98, 10), 932 => to_unsigned(935, 10), 933 => to_unsigned(203, 10), 934 => to_unsigned(411, 10), 935 => to_unsigned(172, 10), 936 => to_unsigned(368, 10), 937 => to_unsigned(55, 10), 938 => to_unsigned(627, 10), 939 => to_unsigned(153, 10), 940 => to_unsigned(803, 10), 941 => to_unsigned(943, 10), 942 => to_unsigned(242, 10), 943 => to_unsigned(25, 10), 944 => to_unsigned(751, 10), 945 => to_unsigned(938, 10), 946 => to_unsigned(439, 10), 947 => to_unsigned(949, 10), 948 => to_unsigned(187, 10), 949 => to_unsigned(296, 10), 950 => to_unsigned(49, 10), 951 => to_unsigned(77, 10), 952 => to_unsigned(602, 10), 953 => to_unsigned(412, 10), 954 => to_unsigned(450, 10), 955 => to_unsigned(580, 10), 956 => to_unsigned(332, 10), 957 => to_unsigned(720, 10), 958 => to_unsigned(300, 10), 959 => to_unsigned(591, 10), 960 => to_unsigned(737, 10), 961 => to_unsigned(99, 10), 962 => to_unsigned(767, 10), 963 => to_unsigned(590, 10), 964 => to_unsigned(658, 10), 965 => to_unsigned(277, 10), 966 => to_unsigned(161, 10), 967 => to_unsigned(412, 10), 968 => to_unsigned(9, 10), 969 => to_unsigned(273, 10), 970 => to_unsigned(776, 10), 971 => to_unsigned(622, 10), 972 => to_unsigned(340, 10), 973 => to_unsigned(537, 10), 974 => to_unsigned(295, 10), 975 => to_unsigned(855, 10), 976 => to_unsigned(773, 10), 977 => to_unsigned(634, 10), 978 => to_unsigned(56, 10), 979 => to_unsigned(838, 10), 980 => to_unsigned(801, 10), 981 => to_unsigned(682, 10), 982 => to_unsigned(738, 10), 983 => to_unsigned(1020, 10), 984 => to_unsigned(1009, 10), 985 => to_unsigned(102, 10), 986 => to_unsigned(284, 10), 987 => to_unsigned(138, 10), 988 => to_unsigned(169, 10), 989 => to_unsigned(877, 10), 990 => to_unsigned(996, 10), 991 => to_unsigned(604, 10), 992 => to_unsigned(774, 10), 993 => to_unsigned(307, 10), 994 => to_unsigned(13, 10), 995 => to_unsigned(398, 10), 996 => to_unsigned(69, 10), 997 => to_unsigned(944, 10), 998 => to_unsigned(850, 10), 999 => to_unsigned(546, 10), 1000 => to_unsigned(300, 10), 1001 => to_unsigned(122, 10), 1002 => to_unsigned(282, 10), 1003 => to_unsigned(561, 10), 1004 => to_unsigned(131, 10), 1005 => to_unsigned(417, 10), 1006 => to_unsigned(94, 10), 1007 => to_unsigned(929, 10), 1008 => to_unsigned(986, 10), 1009 => to_unsigned(434, 10), 1010 => to_unsigned(678, 10), 1011 => to_unsigned(186, 10), 1012 => to_unsigned(1001, 10), 1013 => to_unsigned(333, 10), 1014 => to_unsigned(637, 10), 1015 => to_unsigned(535, 10), 1016 => to_unsigned(73, 10), 1017 => to_unsigned(483, 10), 1018 => to_unsigned(828, 10), 1019 => to_unsigned(301, 10), 1020 => to_unsigned(685, 10), 1021 => to_unsigned(913, 10), 1022 => to_unsigned(714, 10), 1023 => to_unsigned(89, 10), 1024 => to_unsigned(368, 10), 1025 => to_unsigned(582, 10), 1026 => to_unsigned(889, 10), 1027 => to_unsigned(249, 10), 1028 => to_unsigned(366, 10), 1029 => to_unsigned(640, 10), 1030 => to_unsigned(1003, 10), 1031 => to_unsigned(303, 10), 1032 => to_unsigned(737, 10), 1033 => to_unsigned(472, 10), 1034 => to_unsigned(997, 10), 1035 => to_unsigned(863, 10), 1036 => to_unsigned(879, 10), 1037 => to_unsigned(296, 10), 1038 => to_unsigned(101, 10), 1039 => to_unsigned(560, 10), 1040 => to_unsigned(451, 10), 1041 => to_unsigned(752, 10), 1042 => to_unsigned(295, 10), 1043 => to_unsigned(68, 10), 1044 => to_unsigned(39, 10), 1045 => to_unsigned(774, 10), 1046 => to_unsigned(50, 10), 1047 => to_unsigned(100, 10), 1048 => to_unsigned(943, 10), 1049 => to_unsigned(857, 10), 1050 => to_unsigned(523, 10), 1051 => to_unsigned(135, 10), 1052 => to_unsigned(29, 10), 1053 => to_unsigned(951, 10), 1054 => to_unsigned(942, 10), 1055 => to_unsigned(13, 10), 1056 => to_unsigned(195, 10), 1057 => to_unsigned(103, 10), 1058 => to_unsigned(19, 10), 1059 => to_unsigned(657, 10), 1060 => to_unsigned(936, 10), 1061 => to_unsigned(137, 10), 1062 => to_unsigned(712, 10), 1063 => to_unsigned(720, 10), 1064 => to_unsigned(844, 10), 1065 => to_unsigned(984, 10), 1066 => to_unsigned(73, 10), 1067 => to_unsigned(872, 10), 1068 => to_unsigned(901, 10), 1069 => to_unsigned(253, 10), 1070 => to_unsigned(889, 10), 1071 => to_unsigned(319, 10), 1072 => to_unsigned(499, 10), 1073 => to_unsigned(548, 10), 1074 => to_unsigned(46, 10), 1075 => to_unsigned(472, 10), 1076 => to_unsigned(631, 10), 1077 => to_unsigned(659, 10), 1078 => to_unsigned(319, 10), 1079 => to_unsigned(83, 10), 1080 => to_unsigned(247, 10), 1081 => to_unsigned(441, 10), 1082 => to_unsigned(519, 10), 1083 => to_unsigned(483, 10), 1084 => to_unsigned(295, 10), 1085 => to_unsigned(451, 10), 1086 => to_unsigned(592, 10), 1087 => to_unsigned(741, 10), 1088 => to_unsigned(394, 10), 1089 => to_unsigned(208, 10), 1090 => to_unsigned(474, 10), 1091 => to_unsigned(806, 10), 1092 => to_unsigned(843, 10), 1093 => to_unsigned(82, 10), 1094 => to_unsigned(739, 10), 1095 => to_unsigned(216, 10), 1096 => to_unsigned(177, 10), 1097 => to_unsigned(370, 10), 1098 => to_unsigned(596, 10), 1099 => to_unsigned(463, 10), 1100 => to_unsigned(265, 10), 1101 => to_unsigned(646, 10), 1102 => to_unsigned(898, 10), 1103 => to_unsigned(983, 10), 1104 => to_unsigned(573, 10), 1105 => to_unsigned(435, 10), 1106 => to_unsigned(839, 10), 1107 => to_unsigned(451, 10), 1108 => to_unsigned(371, 10), 1109 => to_unsigned(211, 10), 1110 => to_unsigned(365, 10), 1111 => to_unsigned(551, 10), 1112 => to_unsigned(910, 10), 1113 => to_unsigned(133, 10), 1114 => to_unsigned(531, 10), 1115 => to_unsigned(366, 10), 1116 => to_unsigned(375, 10), 1117 => to_unsigned(744, 10), 1118 => to_unsigned(194, 10), 1119 => to_unsigned(753, 10), 1120 => to_unsigned(682, 10), 1121 => to_unsigned(1002, 10), 1122 => to_unsigned(973, 10), 1123 => to_unsigned(408, 10), 1124 => to_unsigned(544, 10), 1125 => to_unsigned(614, 10), 1126 => to_unsigned(325, 10), 1127 => to_unsigned(811, 10), 1128 => to_unsigned(951, 10), 1129 => to_unsigned(27, 10), 1130 => to_unsigned(618, 10), 1131 => to_unsigned(0, 10), 1132 => to_unsigned(273, 10), 1133 => to_unsigned(122, 10), 1134 => to_unsigned(872, 10), 1135 => to_unsigned(358, 10), 1136 => to_unsigned(591, 10), 1137 => to_unsigned(410, 10), 1138 => to_unsigned(590, 10), 1139 => to_unsigned(408, 10), 1140 => to_unsigned(706, 10), 1141 => to_unsigned(89, 10), 1142 => to_unsigned(776, 10), 1143 => to_unsigned(950, 10), 1144 => to_unsigned(190, 10), 1145 => to_unsigned(460, 10), 1146 => to_unsigned(603, 10), 1147 => to_unsigned(528, 10), 1148 => to_unsigned(882, 10), 1149 => to_unsigned(531, 10), 1150 => to_unsigned(1002, 10), 1151 => to_unsigned(54, 10), 1152 => to_unsigned(184, 10), 1153 => to_unsigned(890, 10), 1154 => to_unsigned(632, 10), 1155 => to_unsigned(880, 10), 1156 => to_unsigned(379, 10), 1157 => to_unsigned(232, 10), 1158 => to_unsigned(190, 10), 1159 => to_unsigned(137, 10), 1160 => to_unsigned(140, 10), 1161 => to_unsigned(949, 10), 1162 => to_unsigned(974, 10), 1163 => to_unsigned(959, 10), 1164 => to_unsigned(849, 10), 1165 => to_unsigned(240, 10), 1166 => to_unsigned(772, 10), 1167 => to_unsigned(407, 10), 1168 => to_unsigned(1010, 10), 1169 => to_unsigned(359, 10), 1170 => to_unsigned(58, 10), 1171 => to_unsigned(417, 10), 1172 => to_unsigned(773, 10), 1173 => to_unsigned(91, 10), 1174 => to_unsigned(525, 10), 1175 => to_unsigned(316, 10), 1176 => to_unsigned(981, 10), 1177 => to_unsigned(684, 10), 1178 => to_unsigned(547, 10), 1179 => to_unsigned(78, 10), 1180 => to_unsigned(18, 10), 1181 => to_unsigned(941, 10), 1182 => to_unsigned(56, 10), 1183 => to_unsigned(887, 10), 1184 => to_unsigned(55, 10), 1185 => to_unsigned(335, 10), 1186 => to_unsigned(445, 10), 1187 => to_unsigned(746, 10), 1188 => to_unsigned(943, 10), 1189 => to_unsigned(62, 10), 1190 => to_unsigned(528, 10), 1191 => to_unsigned(362, 10), 1192 => to_unsigned(804, 10), 1193 => to_unsigned(220, 10), 1194 => to_unsigned(694, 10), 1195 => to_unsigned(320, 10), 1196 => to_unsigned(874, 10), 1197 => to_unsigned(606, 10), 1198 => to_unsigned(40, 10), 1199 => to_unsigned(616, 10), 1200 => to_unsigned(429, 10), 1201 => to_unsigned(906, 10), 1202 => to_unsigned(760, 10), 1203 => to_unsigned(664, 10), 1204 => to_unsigned(146, 10), 1205 => to_unsigned(1014, 10), 1206 => to_unsigned(289, 10), 1207 => to_unsigned(297, 10), 1208 => to_unsigned(774, 10), 1209 => to_unsigned(995, 10), 1210 => to_unsigned(697, 10), 1211 => to_unsigned(511, 10), 1212 => to_unsigned(749, 10), 1213 => to_unsigned(450, 10), 1214 => to_unsigned(374, 10), 1215 => to_unsigned(623, 10), 1216 => to_unsigned(336, 10), 1217 => to_unsigned(670, 10), 1218 => to_unsigned(253, 10), 1219 => to_unsigned(626, 10), 1220 => to_unsigned(572, 10), 1221 => to_unsigned(110, 10), 1222 => to_unsigned(754, 10), 1223 => to_unsigned(319, 10), 1224 => to_unsigned(337, 10), 1225 => to_unsigned(287, 10), 1226 => to_unsigned(699, 10), 1227 => to_unsigned(504, 10), 1228 => to_unsigned(661, 10), 1229 => to_unsigned(736, 10), 1230 => to_unsigned(445, 10), 1231 => to_unsigned(87, 10), 1232 => to_unsigned(497, 10), 1233 => to_unsigned(189, 10), 1234 => to_unsigned(635, 10), 1235 => to_unsigned(924, 10), 1236 => to_unsigned(731, 10), 1237 => to_unsigned(779, 10), 1238 => to_unsigned(841, 10), 1239 => to_unsigned(899, 10), 1240 => to_unsigned(720, 10), 1241 => to_unsigned(947, 10), 1242 => to_unsigned(841, 10), 1243 => to_unsigned(915, 10), 1244 => to_unsigned(67, 10), 1245 => to_unsigned(800, 10), 1246 => to_unsigned(368, 10), 1247 => to_unsigned(73, 10), 1248 => to_unsigned(106, 10), 1249 => to_unsigned(744, 10), 1250 => to_unsigned(782, 10), 1251 => to_unsigned(57, 10), 1252 => to_unsigned(229, 10), 1253 => to_unsigned(303, 10), 1254 => to_unsigned(827, 10), 1255 => to_unsigned(216, 10), 1256 => to_unsigned(660, 10), 1257 => to_unsigned(353, 10), 1258 => to_unsigned(852, 10), 1259 => to_unsigned(728, 10), 1260 => to_unsigned(998, 10), 1261 => to_unsigned(519, 10), 1262 => to_unsigned(460, 10), 1263 => to_unsigned(510, 10), 1264 => to_unsigned(138, 10), 1265 => to_unsigned(456, 10), 1266 => to_unsigned(499, 10), 1267 => to_unsigned(513, 10), 1268 => to_unsigned(988, 10), 1269 => to_unsigned(754, 10), 1270 => to_unsigned(92, 10), 1271 => to_unsigned(38, 10), 1272 => to_unsigned(464, 10), 1273 => to_unsigned(156, 10), 1274 => to_unsigned(878, 10), 1275 => to_unsigned(69, 10), 1276 => to_unsigned(801, 10), 1277 => to_unsigned(324, 10), 1278 => to_unsigned(550, 10), 1279 => to_unsigned(636, 10), 1280 => to_unsigned(875, 10), 1281 => to_unsigned(558, 10), 1282 => to_unsigned(778, 10), 1283 => to_unsigned(255, 10), 1284 => to_unsigned(415, 10), 1285 => to_unsigned(660, 10), 1286 => to_unsigned(747, 10), 1287 => to_unsigned(476, 10), 1288 => to_unsigned(775, 10), 1289 => to_unsigned(796, 10), 1290 => to_unsigned(790, 10), 1291 => to_unsigned(906, 10), 1292 => to_unsigned(133, 10), 1293 => to_unsigned(756, 10), 1294 => to_unsigned(893, 10), 1295 => to_unsigned(446, 10), 1296 => to_unsigned(78, 10), 1297 => to_unsigned(322, 10), 1298 => to_unsigned(735, 10), 1299 => to_unsigned(852, 10), 1300 => to_unsigned(6, 10), 1301 => to_unsigned(74, 10), 1302 => to_unsigned(300, 10), 1303 => to_unsigned(114, 10), 1304 => to_unsigned(888, 10), 1305 => to_unsigned(900, 10), 1306 => to_unsigned(835, 10), 1307 => to_unsigned(748, 10), 1308 => to_unsigned(252, 10), 1309 => to_unsigned(623, 10), 1310 => to_unsigned(195, 10), 1311 => to_unsigned(92, 10), 1312 => to_unsigned(336, 10), 1313 => to_unsigned(335, 10), 1314 => to_unsigned(635, 10), 1315 => to_unsigned(915, 10), 1316 => to_unsigned(583, 10), 1317 => to_unsigned(586, 10), 1318 => to_unsigned(826, 10), 1319 => to_unsigned(451, 10), 1320 => to_unsigned(123, 10), 1321 => to_unsigned(36, 10), 1322 => to_unsigned(272, 10), 1323 => to_unsigned(890, 10), 1324 => to_unsigned(753, 10), 1325 => to_unsigned(972, 10), 1326 => to_unsigned(541, 10), 1327 => to_unsigned(364, 10), 1328 => to_unsigned(677, 10), 1329 => to_unsigned(176, 10), 1330 => to_unsigned(478, 10), 1331 => to_unsigned(862, 10), 1332 => to_unsigned(362, 10), 1333 => to_unsigned(457, 10), 1334 => to_unsigned(462, 10), 1335 => to_unsigned(783, 10), 1336 => to_unsigned(199, 10), 1337 => to_unsigned(870, 10), 1338 => to_unsigned(214, 10), 1339 => to_unsigned(426, 10), 1340 => to_unsigned(786, 10), 1341 => to_unsigned(23, 10), 1342 => to_unsigned(208, 10), 1343 => to_unsigned(948, 10), 1344 => to_unsigned(702, 10), 1345 => to_unsigned(824, 10), 1346 => to_unsigned(262, 10), 1347 => to_unsigned(682, 10), 1348 => to_unsigned(689, 10), 1349 => to_unsigned(108, 10), 1350 => to_unsigned(696, 10), 1351 => to_unsigned(701, 10), 1352 => to_unsigned(187, 10), 1353 => to_unsigned(633, 10), 1354 => to_unsigned(598, 10), 1355 => to_unsigned(414, 10), 1356 => to_unsigned(798, 10), 1357 => to_unsigned(171, 10), 1358 => to_unsigned(742, 10), 1359 => to_unsigned(778, 10), 1360 => to_unsigned(625, 10), 1361 => to_unsigned(510, 10), 1362 => to_unsigned(309, 10), 1363 => to_unsigned(961, 10), 1364 => to_unsigned(359, 10), 1365 => to_unsigned(85, 10), 1366 => to_unsigned(566, 10), 1367 => to_unsigned(685, 10), 1368 => to_unsigned(604, 10), 1369 => to_unsigned(455, 10), 1370 => to_unsigned(234, 10), 1371 => to_unsigned(853, 10), 1372 => to_unsigned(32, 10), 1373 => to_unsigned(78, 10), 1374 => to_unsigned(745, 10), 1375 => to_unsigned(728, 10), 1376 => to_unsigned(178, 10), 1377 => to_unsigned(10, 10), 1378 => to_unsigned(427, 10), 1379 => to_unsigned(8, 10), 1380 => to_unsigned(696, 10), 1381 => to_unsigned(140, 10), 1382 => to_unsigned(498, 10), 1383 => to_unsigned(186, 10), 1384 => to_unsigned(538, 10), 1385 => to_unsigned(5, 10), 1386 => to_unsigned(1010, 10), 1387 => to_unsigned(508, 10), 1388 => to_unsigned(819, 10), 1389 => to_unsigned(962, 10), 1390 => to_unsigned(665, 10), 1391 => to_unsigned(91, 10), 1392 => to_unsigned(548, 10), 1393 => to_unsigned(875, 10), 1394 => to_unsigned(627, 10), 1395 => to_unsigned(55, 10), 1396 => to_unsigned(116, 10), 1397 => to_unsigned(185, 10), 1398 => to_unsigned(245, 10), 1399 => to_unsigned(437, 10), 1400 => to_unsigned(162, 10), 1401 => to_unsigned(749, 10), 1402 => to_unsigned(111, 10), 1403 => to_unsigned(893, 10), 1404 => to_unsigned(30, 10), 1405 => to_unsigned(633, 10), 1406 => to_unsigned(511, 10), 1407 => to_unsigned(746, 10), 1408 => to_unsigned(76, 10), 1409 => to_unsigned(192, 10), 1410 => to_unsigned(1012, 10), 1411 => to_unsigned(915, 10), 1412 => to_unsigned(578, 10), 1413 => to_unsigned(844, 10), 1414 => to_unsigned(542, 10), 1415 => to_unsigned(23, 10), 1416 => to_unsigned(705, 10), 1417 => to_unsigned(838, 10), 1418 => to_unsigned(13, 10), 1419 => to_unsigned(408, 10), 1420 => to_unsigned(785, 10), 1421 => to_unsigned(309, 10), 1422 => to_unsigned(49, 10), 1423 => to_unsigned(807, 10), 1424 => to_unsigned(947, 10), 1425 => to_unsigned(914, 10), 1426 => to_unsigned(626, 10), 1427 => to_unsigned(540, 10), 1428 => to_unsigned(77, 10), 1429 => to_unsigned(987, 10), 1430 => to_unsigned(502, 10), 1431 => to_unsigned(172, 10), 1432 => to_unsigned(778, 10), 1433 => to_unsigned(355, 10), 1434 => to_unsigned(834, 10), 1435 => to_unsigned(319, 10), 1436 => to_unsigned(203, 10), 1437 => to_unsigned(728, 10), 1438 => to_unsigned(296, 10), 1439 => to_unsigned(242, 10), 1440 => to_unsigned(381, 10), 1441 => to_unsigned(147, 10), 1442 => to_unsigned(375, 10), 1443 => to_unsigned(148, 10), 1444 => to_unsigned(96, 10), 1445 => to_unsigned(687, 10), 1446 => to_unsigned(124, 10), 1447 => to_unsigned(223, 10), 1448 => to_unsigned(128, 10), 1449 => to_unsigned(302, 10), 1450 => to_unsigned(102, 10), 1451 => to_unsigned(970, 10), 1452 => to_unsigned(268, 10), 1453 => to_unsigned(207, 10), 1454 => to_unsigned(831, 10), 1455 => to_unsigned(494, 10), 1456 => to_unsigned(109, 10), 1457 => to_unsigned(749, 10), 1458 => to_unsigned(974, 10), 1459 => to_unsigned(454, 10), 1460 => to_unsigned(275, 10), 1461 => to_unsigned(110, 10), 1462 => to_unsigned(576, 10), 1463 => to_unsigned(587, 10), 1464 => to_unsigned(25, 10), 1465 => to_unsigned(783, 10), 1466 => to_unsigned(676, 10), 1467 => to_unsigned(720, 10), 1468 => to_unsigned(621, 10), 1469 => to_unsigned(363, 10), 1470 => to_unsigned(986, 10), 1471 => to_unsigned(937, 10), 1472 => to_unsigned(894, 10), 1473 => to_unsigned(33, 10), 1474 => to_unsigned(590, 10), 1475 => to_unsigned(262, 10), 1476 => to_unsigned(739, 10), 1477 => to_unsigned(164, 10), 1478 => to_unsigned(726, 10), 1479 => to_unsigned(666, 10), 1480 => to_unsigned(27, 10), 1481 => to_unsigned(59, 10), 1482 => to_unsigned(843, 10), 1483 => to_unsigned(415, 10), 1484 => to_unsigned(259, 10), 1485 => to_unsigned(227, 10), 1486 => to_unsigned(781, 10), 1487 => to_unsigned(479, 10), 1488 => to_unsigned(526, 10), 1489 => to_unsigned(831, 10), 1490 => to_unsigned(118, 10), 1491 => to_unsigned(555, 10), 1492 => to_unsigned(658, 10), 1493 => to_unsigned(394, 10), 1494 => to_unsigned(379, 10), 1495 => to_unsigned(826, 10), 1496 => to_unsigned(550, 10), 1497 => to_unsigned(447, 10), 1498 => to_unsigned(320, 10), 1499 => to_unsigned(32, 10), 1500 => to_unsigned(993, 10), 1501 => to_unsigned(1000, 10), 1502 => to_unsigned(949, 10), 1503 => to_unsigned(705, 10), 1504 => to_unsigned(751, 10), 1505 => to_unsigned(78, 10), 1506 => to_unsigned(701, 10), 1507 => to_unsigned(991, 10), 1508 => to_unsigned(242, 10), 1509 => to_unsigned(835, 10), 1510 => to_unsigned(149, 10), 1511 => to_unsigned(131, 10), 1512 => to_unsigned(728, 10), 1513 => to_unsigned(266, 10), 1514 => to_unsigned(836, 10), 1515 => to_unsigned(199, 10), 1516 => to_unsigned(270, 10), 1517 => to_unsigned(955, 10), 1518 => to_unsigned(930, 10), 1519 => to_unsigned(619, 10), 1520 => to_unsigned(71, 10), 1521 => to_unsigned(558, 10), 1522 => to_unsigned(232, 10), 1523 => to_unsigned(356, 10), 1524 => to_unsigned(147, 10), 1525 => to_unsigned(266, 10), 1526 => to_unsigned(473, 10), 1527 => to_unsigned(741, 10), 1528 => to_unsigned(707, 10), 1529 => to_unsigned(535, 10), 1530 => to_unsigned(849, 10), 1531 => to_unsigned(350, 10), 1532 => to_unsigned(278, 10), 1533 => to_unsigned(250, 10), 1534 => to_unsigned(110, 10), 1535 => to_unsigned(3, 10), 1536 => to_unsigned(892, 10), 1537 => to_unsigned(808, 10), 1538 => to_unsigned(8, 10), 1539 => to_unsigned(746, 10), 1540 => to_unsigned(149, 10), 1541 => to_unsigned(956, 10), 1542 => to_unsigned(686, 10), 1543 => to_unsigned(582, 10), 1544 => to_unsigned(334, 10), 1545 => to_unsigned(276, 10), 1546 => to_unsigned(230, 10), 1547 => to_unsigned(944, 10), 1548 => to_unsigned(753, 10), 1549 => to_unsigned(210, 10), 1550 => to_unsigned(76, 10), 1551 => to_unsigned(445, 10), 1552 => to_unsigned(659, 10), 1553 => to_unsigned(226, 10), 1554 => to_unsigned(855, 10), 1555 => to_unsigned(440, 10), 1556 => to_unsigned(230, 10), 1557 => to_unsigned(907, 10), 1558 => to_unsigned(50, 10), 1559 => to_unsigned(626, 10), 1560 => to_unsigned(233, 10), 1561 => to_unsigned(815, 10), 1562 => to_unsigned(11, 10), 1563 => to_unsigned(1006, 10), 1564 => to_unsigned(741, 10), 1565 => to_unsigned(304, 10), 1566 => to_unsigned(434, 10), 1567 => to_unsigned(849, 10), 1568 => to_unsigned(1000, 10), 1569 => to_unsigned(171, 10), 1570 => to_unsigned(280, 10), 1571 => to_unsigned(269, 10), 1572 => to_unsigned(115, 10), 1573 => to_unsigned(824, 10), 1574 => to_unsigned(655, 10), 1575 => to_unsigned(687, 10), 1576 => to_unsigned(147, 10), 1577 => to_unsigned(882, 10), 1578 => to_unsigned(294, 10), 1579 => to_unsigned(379, 10), 1580 => to_unsigned(447, 10), 1581 => to_unsigned(48, 10), 1582 => to_unsigned(340, 10), 1583 => to_unsigned(918, 10), 1584 => to_unsigned(40, 10), 1585 => to_unsigned(293, 10), 1586 => to_unsigned(40, 10), 1587 => to_unsigned(720, 10), 1588 => to_unsigned(684, 10), 1589 => to_unsigned(182, 10), 1590 => to_unsigned(94, 10), 1591 => to_unsigned(392, 10), 1592 => to_unsigned(375, 10), 1593 => to_unsigned(446, 10), 1594 => to_unsigned(208, 10), 1595 => to_unsigned(1002, 10), 1596 => to_unsigned(174, 10), 1597 => to_unsigned(797, 10), 1598 => to_unsigned(841, 10), 1599 => to_unsigned(260, 10), 1600 => to_unsigned(644, 10), 1601 => to_unsigned(32, 10), 1602 => to_unsigned(263, 10), 1603 => to_unsigned(140, 10), 1604 => to_unsigned(110, 10), 1605 => to_unsigned(726, 10), 1606 => to_unsigned(390, 10), 1607 => to_unsigned(20, 10), 1608 => to_unsigned(1003, 10), 1609 => to_unsigned(925, 10), 1610 => to_unsigned(209, 10), 1611 => to_unsigned(324, 10), 1612 => to_unsigned(365, 10), 1613 => to_unsigned(381, 10), 1614 => to_unsigned(937, 10), 1615 => to_unsigned(756, 10), 1616 => to_unsigned(895, 10), 1617 => to_unsigned(162, 10), 1618 => to_unsigned(977, 10), 1619 => to_unsigned(387, 10), 1620 => to_unsigned(318, 10), 1621 => to_unsigned(844, 10), 1622 => to_unsigned(943, 10), 1623 => to_unsigned(479, 10), 1624 => to_unsigned(904, 10), 1625 => to_unsigned(302, 10), 1626 => to_unsigned(668, 10), 1627 => to_unsigned(620, 10), 1628 => to_unsigned(13, 10), 1629 => to_unsigned(500, 10), 1630 => to_unsigned(481, 10), 1631 => to_unsigned(348, 10), 1632 => to_unsigned(665, 10), 1633 => to_unsigned(973, 10), 1634 => to_unsigned(859, 10), 1635 => to_unsigned(29, 10), 1636 => to_unsigned(7, 10), 1637 => to_unsigned(474, 10), 1638 => to_unsigned(2, 10), 1639 => to_unsigned(458, 10), 1640 => to_unsigned(388, 10), 1641 => to_unsigned(957, 10), 1642 => to_unsigned(377, 10), 1643 => to_unsigned(730, 10), 1644 => to_unsigned(435, 10), 1645 => to_unsigned(706, 10), 1646 => to_unsigned(540, 10), 1647 => to_unsigned(440, 10), 1648 => to_unsigned(714, 10), 1649 => to_unsigned(340, 10), 1650 => to_unsigned(708, 10), 1651 => to_unsigned(184, 10), 1652 => to_unsigned(506, 10), 1653 => to_unsigned(526, 10), 1654 => to_unsigned(966, 10), 1655 => to_unsigned(349, 10), 1656 => to_unsigned(87, 10), 1657 => to_unsigned(66, 10), 1658 => to_unsigned(182, 10), 1659 => to_unsigned(798, 10), 1660 => to_unsigned(323, 10), 1661 => to_unsigned(605, 10), 1662 => to_unsigned(20, 10), 1663 => to_unsigned(182, 10), 1664 => to_unsigned(335, 10), 1665 => to_unsigned(922, 10), 1666 => to_unsigned(446, 10), 1667 => to_unsigned(1018, 10), 1668 => to_unsigned(57, 10), 1669 => to_unsigned(248, 10), 1670 => to_unsigned(347, 10), 1671 => to_unsigned(472, 10), 1672 => to_unsigned(1001, 10), 1673 => to_unsigned(709, 10), 1674 => to_unsigned(973, 10), 1675 => to_unsigned(653, 10), 1676 => to_unsigned(193, 10), 1677 => to_unsigned(249, 10), 1678 => to_unsigned(742, 10), 1679 => to_unsigned(13, 10), 1680 => to_unsigned(58, 10), 1681 => to_unsigned(680, 10), 1682 => to_unsigned(968, 10), 1683 => to_unsigned(484, 10), 1684 => to_unsigned(1018, 10), 1685 => to_unsigned(123, 10), 1686 => to_unsigned(391, 10), 1687 => to_unsigned(151, 10), 1688 => to_unsigned(331, 10), 1689 => to_unsigned(580, 10), 1690 => to_unsigned(689, 10), 1691 => to_unsigned(578, 10), 1692 => to_unsigned(728, 10), 1693 => to_unsigned(700, 10), 1694 => to_unsigned(445, 10), 1695 => to_unsigned(479, 10), 1696 => to_unsigned(816, 10), 1697 => to_unsigned(814, 10), 1698 => to_unsigned(1005, 10), 1699 => to_unsigned(632, 10), 1700 => to_unsigned(576, 10), 1701 => to_unsigned(733, 10), 1702 => to_unsigned(617, 10), 1703 => to_unsigned(989, 10), 1704 => to_unsigned(843, 10), 1705 => to_unsigned(25, 10), 1706 => to_unsigned(719, 10), 1707 => to_unsigned(471, 10), 1708 => to_unsigned(777, 10), 1709 => to_unsigned(195, 10), 1710 => to_unsigned(427, 10), 1711 => to_unsigned(327, 10), 1712 => to_unsigned(124, 10), 1713 => to_unsigned(990, 10), 1714 => to_unsigned(1009, 10), 1715 => to_unsigned(266, 10), 1716 => to_unsigned(656, 10), 1717 => to_unsigned(194, 10), 1718 => to_unsigned(218, 10), 1719 => to_unsigned(802, 10), 1720 => to_unsigned(307, 10), 1721 => to_unsigned(52, 10), 1722 => to_unsigned(989, 10), 1723 => to_unsigned(829, 10), 1724 => to_unsigned(809, 10), 1725 => to_unsigned(267, 10), 1726 => to_unsigned(158, 10), 1727 => to_unsigned(180, 10), 1728 => to_unsigned(692, 10), 1729 => to_unsigned(68, 10), 1730 => to_unsigned(799, 10), 1731 => to_unsigned(1023, 10), 1732 => to_unsigned(932, 10), 1733 => to_unsigned(406, 10), 1734 => to_unsigned(870, 10), 1735 => to_unsigned(693, 10), 1736 => to_unsigned(799, 10), 1737 => to_unsigned(792, 10), 1738 => to_unsigned(351, 10), 1739 => to_unsigned(168, 10), 1740 => to_unsigned(6, 10), 1741 => to_unsigned(891, 10), 1742 => to_unsigned(833, 10), 1743 => to_unsigned(753, 10), 1744 => to_unsigned(389, 10), 1745 => to_unsigned(691, 10), 1746 => to_unsigned(433, 10), 1747 => to_unsigned(515, 10), 1748 => to_unsigned(247, 10), 1749 => to_unsigned(537, 10), 1750 => to_unsigned(5, 10), 1751 => to_unsigned(738, 10), 1752 => to_unsigned(382, 10), 1753 => to_unsigned(800, 10), 1754 => to_unsigned(750, 10), 1755 => to_unsigned(779, 10), 1756 => to_unsigned(844, 10), 1757 => to_unsigned(215, 10), 1758 => to_unsigned(965, 10), 1759 => to_unsigned(646, 10), 1760 => to_unsigned(847, 10), 1761 => to_unsigned(185, 10), 1762 => to_unsigned(315, 10), 1763 => to_unsigned(498, 10), 1764 => to_unsigned(967, 10), 1765 => to_unsigned(682, 10), 1766 => to_unsigned(647, 10), 1767 => to_unsigned(56, 10), 1768 => to_unsigned(262, 10), 1769 => to_unsigned(413, 10), 1770 => to_unsigned(174, 10), 1771 => to_unsigned(267, 10), 1772 => to_unsigned(611, 10), 1773 => to_unsigned(257, 10), 1774 => to_unsigned(44, 10), 1775 => to_unsigned(190, 10), 1776 => to_unsigned(274, 10), 1777 => to_unsigned(687, 10), 1778 => to_unsigned(1022, 10), 1779 => to_unsigned(998, 10), 1780 => to_unsigned(780, 10), 1781 => to_unsigned(866, 10), 1782 => to_unsigned(566, 10), 1783 => to_unsigned(441, 10), 1784 => to_unsigned(448, 10), 1785 => to_unsigned(283, 10), 1786 => to_unsigned(826, 10), 1787 => to_unsigned(391, 10), 1788 => to_unsigned(682, 10), 1789 => to_unsigned(995, 10), 1790 => to_unsigned(976, 10), 1791 => to_unsigned(114, 10), 1792 => to_unsigned(583, 10), 1793 => to_unsigned(431, 10), 1794 => to_unsigned(287, 10), 1795 => to_unsigned(660, 10), 1796 => to_unsigned(361, 10), 1797 => to_unsigned(304, 10), 1798 => to_unsigned(260, 10), 1799 => to_unsigned(514, 10), 1800 => to_unsigned(224, 10), 1801 => to_unsigned(875, 10), 1802 => to_unsigned(669, 10), 1803 => to_unsigned(984, 10), 1804 => to_unsigned(485, 10), 1805 => to_unsigned(394, 10), 1806 => to_unsigned(921, 10), 1807 => to_unsigned(508, 10), 1808 => to_unsigned(131, 10), 1809 => to_unsigned(64, 10), 1810 => to_unsigned(969, 10), 1811 => to_unsigned(57, 10), 1812 => to_unsigned(580, 10), 1813 => to_unsigned(504, 10), 1814 => to_unsigned(472, 10), 1815 => to_unsigned(900, 10), 1816 => to_unsigned(353, 10), 1817 => to_unsigned(480, 10), 1818 => to_unsigned(11, 10), 1819 => to_unsigned(285, 10), 1820 => to_unsigned(226, 10), 1821 => to_unsigned(703, 10), 1822 => to_unsigned(48, 10), 1823 => to_unsigned(611, 10), 1824 => to_unsigned(545, 10), 1825 => to_unsigned(508, 10), 1826 => to_unsigned(379, 10), 1827 => to_unsigned(539, 10), 1828 => to_unsigned(544, 10), 1829 => to_unsigned(908, 10), 1830 => to_unsigned(524, 10), 1831 => to_unsigned(771, 10), 1832 => to_unsigned(995, 10), 1833 => to_unsigned(1017, 10), 1834 => to_unsigned(118, 10), 1835 => to_unsigned(693, 10), 1836 => to_unsigned(901, 10), 1837 => to_unsigned(903, 10), 1838 => to_unsigned(96, 10), 1839 => to_unsigned(228, 10), 1840 => to_unsigned(598, 10), 1841 => to_unsigned(978, 10), 1842 => to_unsigned(91, 10), 1843 => to_unsigned(159, 10), 1844 => to_unsigned(717, 10), 1845 => to_unsigned(582, 10), 1846 => to_unsigned(922, 10), 1847 => to_unsigned(519, 10), 1848 => to_unsigned(221, 10), 1849 => to_unsigned(99, 10), 1850 => to_unsigned(285, 10), 1851 => to_unsigned(253, 10), 1852 => to_unsigned(278, 10), 1853 => to_unsigned(684, 10), 1854 => to_unsigned(304, 10), 1855 => to_unsigned(738, 10), 1856 => to_unsigned(225, 10), 1857 => to_unsigned(868, 10), 1858 => to_unsigned(942, 10), 1859 => to_unsigned(303, 10), 1860 => to_unsigned(474, 10), 1861 => to_unsigned(631, 10), 1862 => to_unsigned(975, 10), 1863 => to_unsigned(563, 10), 1864 => to_unsigned(213, 10), 1865 => to_unsigned(648, 10), 1866 => to_unsigned(115, 10), 1867 => to_unsigned(40, 10), 1868 => to_unsigned(979, 10), 1869 => to_unsigned(162, 10), 1870 => to_unsigned(633, 10), 1871 => to_unsigned(422, 10), 1872 => to_unsigned(283, 10), 1873 => to_unsigned(626, 10), 1874 => to_unsigned(846, 10), 1875 => to_unsigned(549, 10), 1876 => to_unsigned(74, 10), 1877 => to_unsigned(355, 10), 1878 => to_unsigned(417, 10), 1879 => to_unsigned(486, 10), 1880 => to_unsigned(597, 10), 1881 => to_unsigned(767, 10), 1882 => to_unsigned(824, 10), 1883 => to_unsigned(334, 10), 1884 => to_unsigned(122, 10), 1885 => to_unsigned(362, 10), 1886 => to_unsigned(759, 10), 1887 => to_unsigned(654, 10), 1888 => to_unsigned(818, 10), 1889 => to_unsigned(630, 10), 1890 => to_unsigned(226, 10), 1891 => to_unsigned(23, 10), 1892 => to_unsigned(731, 10), 1893 => to_unsigned(615, 10), 1894 => to_unsigned(144, 10), 1895 => to_unsigned(831, 10), 1896 => to_unsigned(739, 10), 1897 => to_unsigned(209, 10), 1898 => to_unsigned(93, 10), 1899 => to_unsigned(680, 10), 1900 => to_unsigned(773, 10), 1901 => to_unsigned(439, 10), 1902 => to_unsigned(669, 10), 1903 => to_unsigned(892, 10), 1904 => to_unsigned(225, 10), 1905 => to_unsigned(45, 10), 1906 => to_unsigned(527, 10), 1907 => to_unsigned(101, 10), 1908 => to_unsigned(758, 10), 1909 => to_unsigned(955, 10), 1910 => to_unsigned(789, 10), 1911 => to_unsigned(263, 10), 1912 => to_unsigned(234, 10), 1913 => to_unsigned(341, 10), 1914 => to_unsigned(19, 10), 1915 => to_unsigned(595, 10), 1916 => to_unsigned(67, 10), 1917 => to_unsigned(369, 10), 1918 => to_unsigned(204, 10), 1919 => to_unsigned(79, 10), 1920 => to_unsigned(198, 10), 1921 => to_unsigned(518, 10), 1922 => to_unsigned(718, 10), 1923 => to_unsigned(450, 10), 1924 => to_unsigned(917, 10), 1925 => to_unsigned(506, 10), 1926 => to_unsigned(195, 10), 1927 => to_unsigned(947, 10), 1928 => to_unsigned(731, 10), 1929 => to_unsigned(606, 10), 1930 => to_unsigned(31, 10), 1931 => to_unsigned(627, 10), 1932 => to_unsigned(481, 10), 1933 => to_unsigned(615, 10), 1934 => to_unsigned(361, 10), 1935 => to_unsigned(829, 10), 1936 => to_unsigned(375, 10), 1937 => to_unsigned(437, 10), 1938 => to_unsigned(672, 10), 1939 => to_unsigned(656, 10), 1940 => to_unsigned(949, 10), 1941 => to_unsigned(327, 10), 1942 => to_unsigned(857, 10), 1943 => to_unsigned(435, 10), 1944 => to_unsigned(882, 10), 1945 => to_unsigned(889, 10), 1946 => to_unsigned(265, 10), 1947 => to_unsigned(904, 10), 1948 => to_unsigned(167, 10), 1949 => to_unsigned(1004, 10), 1950 => to_unsigned(82, 10), 1951 => to_unsigned(522, 10), 1952 => to_unsigned(909, 10), 1953 => to_unsigned(671, 10), 1954 => to_unsigned(556, 10), 1955 => to_unsigned(352, 10), 1956 => to_unsigned(607, 10), 1957 => to_unsigned(454, 10), 1958 => to_unsigned(322, 10), 1959 => to_unsigned(680, 10), 1960 => to_unsigned(445, 10), 1961 => to_unsigned(1016, 10), 1962 => to_unsigned(238, 10), 1963 => to_unsigned(731, 10), 1964 => to_unsigned(469, 10), 1965 => to_unsigned(756, 10), 1966 => to_unsigned(940, 10), 1967 => to_unsigned(603, 10), 1968 => to_unsigned(992, 10), 1969 => to_unsigned(767, 10), 1970 => to_unsigned(552, 10), 1971 => to_unsigned(138, 10), 1972 => to_unsigned(180, 10), 1973 => to_unsigned(709, 10), 1974 => to_unsigned(394, 10), 1975 => to_unsigned(90, 10), 1976 => to_unsigned(1014, 10), 1977 => to_unsigned(886, 10), 1978 => to_unsigned(917, 10), 1979 => to_unsigned(676, 10), 1980 => to_unsigned(690, 10), 1981 => to_unsigned(751, 10), 1982 => to_unsigned(276, 10), 1983 => to_unsigned(440, 10), 1984 => to_unsigned(383, 10), 1985 => to_unsigned(101, 10), 1986 => to_unsigned(696, 10), 1987 => to_unsigned(441, 10), 1988 => to_unsigned(658, 10), 1989 => to_unsigned(402, 10), 1990 => to_unsigned(540, 10), 1991 => to_unsigned(898, 10), 1992 => to_unsigned(561, 10), 1993 => to_unsigned(303, 10), 1994 => to_unsigned(179, 10), 1995 => to_unsigned(483, 10), 1996 => to_unsigned(758, 10), 1997 => to_unsigned(720, 10), 1998 => to_unsigned(113, 10), 1999 => to_unsigned(462, 10), 2000 => to_unsigned(398, 10), 2001 => to_unsigned(776, 10), 2002 => to_unsigned(958, 10), 2003 => to_unsigned(773, 10), 2004 => to_unsigned(324, 10), 2005 => to_unsigned(555, 10), 2006 => to_unsigned(421, 10), 2007 => to_unsigned(453, 10), 2008 => to_unsigned(814, 10), 2009 => to_unsigned(196, 10), 2010 => to_unsigned(41, 10), 2011 => to_unsigned(910, 10), 2012 => to_unsigned(528, 10), 2013 => to_unsigned(216, 10), 2014 => to_unsigned(181, 10), 2015 => to_unsigned(794, 10), 2016 => to_unsigned(57, 10), 2017 => to_unsigned(777, 10), 2018 => to_unsigned(560, 10), 2019 => to_unsigned(84, 10), 2020 => to_unsigned(90, 10), 2021 => to_unsigned(0, 10), 2022 => to_unsigned(205, 10), 2023 => to_unsigned(131, 10), 2024 => to_unsigned(322, 10), 2025 => to_unsigned(10, 10), 2026 => to_unsigned(1005, 10), 2027 => to_unsigned(720, 10), 2028 => to_unsigned(699, 10), 2029 => to_unsigned(514, 10), 2030 => to_unsigned(966, 10), 2031 => to_unsigned(444, 10), 2032 => to_unsigned(1008, 10), 2033 => to_unsigned(316, 10), 2034 => to_unsigned(863, 10), 2035 => to_unsigned(156, 10), 2036 => to_unsigned(501, 10), 2037 => to_unsigned(184, 10), 2038 => to_unsigned(852, 10), 2039 => to_unsigned(262, 10), 2040 => to_unsigned(17, 10), 2041 => to_unsigned(1019, 10), 2042 => to_unsigned(947, 10), 2043 => to_unsigned(788, 10), 2044 => to_unsigned(347, 10), 2045 => to_unsigned(658, 10), 2046 => to_unsigned(498, 10), 2047 => to_unsigned(197, 10)),
            8 => (0 => to_unsigned(723, 10), 1 => to_unsigned(561, 10), 2 => to_unsigned(513, 10), 3 => to_unsigned(143, 10), 4 => to_unsigned(336, 10), 5 => to_unsigned(397, 10), 6 => to_unsigned(840, 10), 7 => to_unsigned(810, 10), 8 => to_unsigned(613, 10), 9 => to_unsigned(755, 10), 10 => to_unsigned(260, 10), 11 => to_unsigned(542, 10), 12 => to_unsigned(934, 10), 13 => to_unsigned(632, 10), 14 => to_unsigned(966, 10), 15 => to_unsigned(883, 10), 16 => to_unsigned(945, 10), 17 => to_unsigned(427, 10), 18 => to_unsigned(857, 10), 19 => to_unsigned(638, 10), 20 => to_unsigned(928, 10), 21 => to_unsigned(223, 10), 22 => to_unsigned(298, 10), 23 => to_unsigned(317, 10), 24 => to_unsigned(117, 10), 25 => to_unsigned(321, 10), 26 => to_unsigned(987, 10), 27 => to_unsigned(448, 10), 28 => to_unsigned(444, 10), 29 => to_unsigned(768, 10), 30 => to_unsigned(911, 10), 31 => to_unsigned(640, 10), 32 => to_unsigned(226, 10), 33 => to_unsigned(999, 10), 34 => to_unsigned(282, 10), 35 => to_unsigned(225, 10), 36 => to_unsigned(753, 10), 37 => to_unsigned(129, 10), 38 => to_unsigned(572, 10), 39 => to_unsigned(223, 10), 40 => to_unsigned(410, 10), 41 => to_unsigned(637, 10), 42 => to_unsigned(419, 10), 43 => to_unsigned(170, 10), 44 => to_unsigned(91, 10), 45 => to_unsigned(724, 10), 46 => to_unsigned(956, 10), 47 => to_unsigned(275, 10), 48 => to_unsigned(723, 10), 49 => to_unsigned(393, 10), 50 => to_unsigned(124, 10), 51 => to_unsigned(965, 10), 52 => to_unsigned(815, 10), 53 => to_unsigned(958, 10), 54 => to_unsigned(386, 10), 55 => to_unsigned(991, 10), 56 => to_unsigned(907, 10), 57 => to_unsigned(881, 10), 58 => to_unsigned(273, 10), 59 => to_unsigned(196, 10), 60 => to_unsigned(463, 10), 61 => to_unsigned(953, 10), 62 => to_unsigned(385, 10), 63 => to_unsigned(384, 10), 64 => to_unsigned(515, 10), 65 => to_unsigned(56, 10), 66 => to_unsigned(322, 10), 67 => to_unsigned(198, 10), 68 => to_unsigned(704, 10), 69 => to_unsigned(322, 10), 70 => to_unsigned(974, 10), 71 => to_unsigned(118, 10), 72 => to_unsigned(546, 10), 73 => to_unsigned(1004, 10), 74 => to_unsigned(351, 10), 75 => to_unsigned(888, 10), 76 => to_unsigned(828, 10), 77 => to_unsigned(127, 10), 78 => to_unsigned(30, 10), 79 => to_unsigned(477, 10), 80 => to_unsigned(894, 10), 81 => to_unsigned(273, 10), 82 => to_unsigned(324, 10), 83 => to_unsigned(192, 10), 84 => to_unsigned(252, 10), 85 => to_unsigned(707, 10), 86 => to_unsigned(951, 10), 87 => to_unsigned(699, 10), 88 => to_unsigned(101, 10), 89 => to_unsigned(215, 10), 90 => to_unsigned(259, 10), 91 => to_unsigned(871, 10), 92 => to_unsigned(262, 10), 93 => to_unsigned(201, 10), 94 => to_unsigned(272, 10), 95 => to_unsigned(632, 10), 96 => to_unsigned(787, 10), 97 => to_unsigned(83, 10), 98 => to_unsigned(788, 10), 99 => to_unsigned(233, 10), 100 => to_unsigned(833, 10), 101 => to_unsigned(286, 10), 102 => to_unsigned(948, 10), 103 => to_unsigned(351, 10), 104 => to_unsigned(679, 10), 105 => to_unsigned(923, 10), 106 => to_unsigned(416, 10), 107 => to_unsigned(597, 10), 108 => to_unsigned(109, 10), 109 => to_unsigned(548, 10), 110 => to_unsigned(641, 10), 111 => to_unsigned(999, 10), 112 => to_unsigned(515, 10), 113 => to_unsigned(682, 10), 114 => to_unsigned(532, 10), 115 => to_unsigned(107, 10), 116 => to_unsigned(85, 10), 117 => to_unsigned(208, 10), 118 => to_unsigned(762, 10), 119 => to_unsigned(906, 10), 120 => to_unsigned(64, 10), 121 => to_unsigned(989, 10), 122 => to_unsigned(648, 10), 123 => to_unsigned(104, 10), 124 => to_unsigned(973, 10), 125 => to_unsigned(948, 10), 126 => to_unsigned(260, 10), 127 => to_unsigned(515, 10), 128 => to_unsigned(322, 10), 129 => to_unsigned(258, 10), 130 => to_unsigned(261, 10), 131 => to_unsigned(818, 10), 132 => to_unsigned(693, 10), 133 => to_unsigned(553, 10), 134 => to_unsigned(649, 10), 135 => to_unsigned(880, 10), 136 => to_unsigned(266, 10), 137 => to_unsigned(451, 10), 138 => to_unsigned(283, 10), 139 => to_unsigned(615, 10), 140 => to_unsigned(987, 10), 141 => to_unsigned(407, 10), 142 => to_unsigned(673, 10), 143 => to_unsigned(511, 10), 144 => to_unsigned(1017, 10), 145 => to_unsigned(84, 10), 146 => to_unsigned(519, 10), 147 => to_unsigned(218, 10), 148 => to_unsigned(890, 10), 149 => to_unsigned(598, 10), 150 => to_unsigned(7, 10), 151 => to_unsigned(623, 10), 152 => to_unsigned(226, 10), 153 => to_unsigned(814, 10), 154 => to_unsigned(751, 10), 155 => to_unsigned(110, 10), 156 => to_unsigned(780, 10), 157 => to_unsigned(787, 10), 158 => to_unsigned(887, 10), 159 => to_unsigned(339, 10), 160 => to_unsigned(492, 10), 161 => to_unsigned(364, 10), 162 => to_unsigned(22, 10), 163 => to_unsigned(450, 10), 164 => to_unsigned(334, 10), 165 => to_unsigned(836, 10), 166 => to_unsigned(206, 10), 167 => to_unsigned(478, 10), 168 => to_unsigned(222, 10), 169 => to_unsigned(277, 10), 170 => to_unsigned(373, 10), 171 => to_unsigned(1018, 10), 172 => to_unsigned(720, 10), 173 => to_unsigned(658, 10), 174 => to_unsigned(352, 10), 175 => to_unsigned(369, 10), 176 => to_unsigned(593, 10), 177 => to_unsigned(970, 10), 178 => to_unsigned(265, 10), 179 => to_unsigned(442, 10), 180 => to_unsigned(606, 10), 181 => to_unsigned(260, 10), 182 => to_unsigned(684, 10), 183 => to_unsigned(161, 10), 184 => to_unsigned(993, 10), 185 => to_unsigned(655, 10), 186 => to_unsigned(254, 10), 187 => to_unsigned(706, 10), 188 => to_unsigned(445, 10), 189 => to_unsigned(680, 10), 190 => to_unsigned(656, 10), 191 => to_unsigned(77, 10), 192 => to_unsigned(149, 10), 193 => to_unsigned(893, 10), 194 => to_unsigned(331, 10), 195 => to_unsigned(505, 10), 196 => to_unsigned(593, 10), 197 => to_unsigned(1010, 10), 198 => to_unsigned(623, 10), 199 => to_unsigned(569, 10), 200 => to_unsigned(998, 10), 201 => to_unsigned(549, 10), 202 => to_unsigned(714, 10), 203 => to_unsigned(361, 10), 204 => to_unsigned(770, 10), 205 => to_unsigned(120, 10), 206 => to_unsigned(727, 10), 207 => to_unsigned(198, 10), 208 => to_unsigned(532, 10), 209 => to_unsigned(20, 10), 210 => to_unsigned(189, 10), 211 => to_unsigned(358, 10), 212 => to_unsigned(901, 10), 213 => to_unsigned(49, 10), 214 => to_unsigned(325, 10), 215 => to_unsigned(373, 10), 216 => to_unsigned(848, 10), 217 => to_unsigned(972, 10), 218 => to_unsigned(918, 10), 219 => to_unsigned(756, 10), 220 => to_unsigned(690, 10), 221 => to_unsigned(207, 10), 222 => to_unsigned(295, 10), 223 => to_unsigned(964, 10), 224 => to_unsigned(935, 10), 225 => to_unsigned(273, 10), 226 => to_unsigned(432, 10), 227 => to_unsigned(351, 10), 228 => to_unsigned(26, 10), 229 => to_unsigned(29, 10), 230 => to_unsigned(651, 10), 231 => to_unsigned(383, 10), 232 => to_unsigned(742, 10), 233 => to_unsigned(321, 10), 234 => to_unsigned(378, 10), 235 => to_unsigned(1010, 10), 236 => to_unsigned(925, 10), 237 => to_unsigned(814, 10), 238 => to_unsigned(253, 10), 239 => to_unsigned(747, 10), 240 => to_unsigned(48, 10), 241 => to_unsigned(119, 10), 242 => to_unsigned(230, 10), 243 => to_unsigned(563, 10), 244 => to_unsigned(895, 10), 245 => to_unsigned(3, 10), 246 => to_unsigned(849, 10), 247 => to_unsigned(318, 10), 248 => to_unsigned(465, 10), 249 => to_unsigned(4, 10), 250 => to_unsigned(978, 10), 251 => to_unsigned(81, 10), 252 => to_unsigned(738, 10), 253 => to_unsigned(707, 10), 254 => to_unsigned(925, 10), 255 => to_unsigned(561, 10), 256 => to_unsigned(113, 10), 257 => to_unsigned(659, 10), 258 => to_unsigned(814, 10), 259 => to_unsigned(338, 10), 260 => to_unsigned(807, 10), 261 => to_unsigned(330, 10), 262 => to_unsigned(637, 10), 263 => to_unsigned(221, 10), 264 => to_unsigned(712, 10), 265 => to_unsigned(638, 10), 266 => to_unsigned(424, 10), 267 => to_unsigned(984, 10), 268 => to_unsigned(98, 10), 269 => to_unsigned(366, 10), 270 => to_unsigned(187, 10), 271 => to_unsigned(213, 10), 272 => to_unsigned(750, 10), 273 => to_unsigned(5, 10), 274 => to_unsigned(68, 10), 275 => to_unsigned(548, 10), 276 => to_unsigned(636, 10), 277 => to_unsigned(551, 10), 278 => to_unsigned(118, 10), 279 => to_unsigned(597, 10), 280 => to_unsigned(761, 10), 281 => to_unsigned(676, 10), 282 => to_unsigned(174, 10), 283 => to_unsigned(716, 10), 284 => to_unsigned(717, 10), 285 => to_unsigned(195, 10), 286 => to_unsigned(173, 10), 287 => to_unsigned(552, 10), 288 => to_unsigned(931, 10), 289 => to_unsigned(617, 10), 290 => to_unsigned(487, 10), 291 => to_unsigned(696, 10), 292 => to_unsigned(1010, 10), 293 => to_unsigned(286, 10), 294 => to_unsigned(426, 10), 295 => to_unsigned(849, 10), 296 => to_unsigned(347, 10), 297 => to_unsigned(323, 10), 298 => to_unsigned(282, 10), 299 => to_unsigned(907, 10), 300 => to_unsigned(42, 10), 301 => to_unsigned(715, 10), 302 => to_unsigned(121, 10), 303 => to_unsigned(147, 10), 304 => to_unsigned(883, 10), 305 => to_unsigned(341, 10), 306 => to_unsigned(899, 10), 307 => to_unsigned(100, 10), 308 => to_unsigned(52, 10), 309 => to_unsigned(382, 10), 310 => to_unsigned(917, 10), 311 => to_unsigned(378, 10), 312 => to_unsigned(745, 10), 313 => to_unsigned(241, 10), 314 => to_unsigned(236, 10), 315 => to_unsigned(743, 10), 316 => to_unsigned(474, 10), 317 => to_unsigned(621, 10), 318 => to_unsigned(733, 10), 319 => to_unsigned(849, 10), 320 => to_unsigned(525, 10), 321 => to_unsigned(190, 10), 322 => to_unsigned(321, 10), 323 => to_unsigned(630, 10), 324 => to_unsigned(789, 10), 325 => to_unsigned(587, 10), 326 => to_unsigned(340, 10), 327 => to_unsigned(201, 10), 328 => to_unsigned(892, 10), 329 => to_unsigned(779, 10), 330 => to_unsigned(647, 10), 331 => to_unsigned(668, 10), 332 => to_unsigned(655, 10), 333 => to_unsigned(357, 10), 334 => to_unsigned(859, 10), 335 => to_unsigned(149, 10), 336 => to_unsigned(281, 10), 337 => to_unsigned(728, 10), 338 => to_unsigned(486, 10), 339 => to_unsigned(201, 10), 340 => to_unsigned(73, 10), 341 => to_unsigned(251, 10), 342 => to_unsigned(929, 10), 343 => to_unsigned(460, 10), 344 => to_unsigned(129, 10), 345 => to_unsigned(860, 10), 346 => to_unsigned(120, 10), 347 => to_unsigned(743, 10), 348 => to_unsigned(1005, 10), 349 => to_unsigned(292, 10), 350 => to_unsigned(220, 10), 351 => to_unsigned(931, 10), 352 => to_unsigned(43, 10), 353 => to_unsigned(195, 10), 354 => to_unsigned(412, 10), 355 => to_unsigned(9, 10), 356 => to_unsigned(163, 10), 357 => to_unsigned(518, 10), 358 => to_unsigned(399, 10), 359 => to_unsigned(886, 10), 360 => to_unsigned(471, 10), 361 => to_unsigned(465, 10), 362 => to_unsigned(742, 10), 363 => to_unsigned(985, 10), 364 => to_unsigned(390, 10), 365 => to_unsigned(593, 10), 366 => to_unsigned(999, 10), 367 => to_unsigned(85, 10), 368 => to_unsigned(637, 10), 369 => to_unsigned(203, 10), 370 => to_unsigned(409, 10), 371 => to_unsigned(808, 10), 372 => to_unsigned(263, 10), 373 => to_unsigned(1004, 10), 374 => to_unsigned(27, 10), 375 => to_unsigned(493, 10), 376 => to_unsigned(906, 10), 377 => to_unsigned(297, 10), 378 => to_unsigned(460, 10), 379 => to_unsigned(831, 10), 380 => to_unsigned(858, 10), 381 => to_unsigned(714, 10), 382 => to_unsigned(740, 10), 383 => to_unsigned(805, 10), 384 => to_unsigned(608, 10), 385 => to_unsigned(5, 10), 386 => to_unsigned(764, 10), 387 => to_unsigned(953, 10), 388 => to_unsigned(313, 10), 389 => to_unsigned(713, 10), 390 => to_unsigned(346, 10), 391 => to_unsigned(43, 10), 392 => to_unsigned(294, 10), 393 => to_unsigned(600, 10), 394 => to_unsigned(644, 10), 395 => to_unsigned(586, 10), 396 => to_unsigned(478, 10), 397 => to_unsigned(217, 10), 398 => to_unsigned(636, 10), 399 => to_unsigned(309, 10), 400 => to_unsigned(175, 10), 401 => to_unsigned(928, 10), 402 => to_unsigned(27, 10), 403 => to_unsigned(89, 10), 404 => to_unsigned(27, 10), 405 => to_unsigned(642, 10), 406 => to_unsigned(318, 10), 407 => to_unsigned(445, 10), 408 => to_unsigned(398, 10), 409 => to_unsigned(875, 10), 410 => to_unsigned(961, 10), 411 => to_unsigned(513, 10), 412 => to_unsigned(776, 10), 413 => to_unsigned(890, 10), 414 => to_unsigned(359, 10), 415 => to_unsigned(568, 10), 416 => to_unsigned(310, 10), 417 => to_unsigned(923, 10), 418 => to_unsigned(60, 10), 419 => to_unsigned(825, 10), 420 => to_unsigned(392, 10), 421 => to_unsigned(21, 10), 422 => to_unsigned(129, 10), 423 => to_unsigned(61, 10), 424 => to_unsigned(516, 10), 425 => to_unsigned(273, 10), 426 => to_unsigned(131, 10), 427 => to_unsigned(286, 10), 428 => to_unsigned(172, 10), 429 => to_unsigned(306, 10), 430 => to_unsigned(87, 10), 431 => to_unsigned(592, 10), 432 => to_unsigned(127, 10), 433 => to_unsigned(345, 10), 434 => to_unsigned(603, 10), 435 => to_unsigned(15, 10), 436 => to_unsigned(536, 10), 437 => to_unsigned(769, 10), 438 => to_unsigned(1011, 10), 439 => to_unsigned(692, 10), 440 => to_unsigned(266, 10), 441 => to_unsigned(329, 10), 442 => to_unsigned(941, 10), 443 => to_unsigned(841, 10), 444 => to_unsigned(641, 10), 445 => to_unsigned(586, 10), 446 => to_unsigned(553, 10), 447 => to_unsigned(106, 10), 448 => to_unsigned(541, 10), 449 => to_unsigned(978, 10), 450 => to_unsigned(588, 10), 451 => to_unsigned(509, 10), 452 => to_unsigned(192, 10), 453 => to_unsigned(443, 10), 454 => to_unsigned(861, 10), 455 => to_unsigned(66, 10), 456 => to_unsigned(581, 10), 457 => to_unsigned(528, 10), 458 => to_unsigned(14, 10), 459 => to_unsigned(10, 10), 460 => to_unsigned(132, 10), 461 => to_unsigned(508, 10), 462 => to_unsigned(446, 10), 463 => to_unsigned(6, 10), 464 => to_unsigned(620, 10), 465 => to_unsigned(151, 10), 466 => to_unsigned(85, 10), 467 => to_unsigned(772, 10), 468 => to_unsigned(55, 10), 469 => to_unsigned(104, 10), 470 => to_unsigned(769, 10), 471 => to_unsigned(463, 10), 472 => to_unsigned(717, 10), 473 => to_unsigned(683, 10), 474 => to_unsigned(1010, 10), 475 => to_unsigned(553, 10), 476 => to_unsigned(432, 10), 477 => to_unsigned(350, 10), 478 => to_unsigned(104, 10), 479 => to_unsigned(483, 10), 480 => to_unsigned(589, 10), 481 => to_unsigned(347, 10), 482 => to_unsigned(39, 10), 483 => to_unsigned(972, 10), 484 => to_unsigned(425, 10), 485 => to_unsigned(774, 10), 486 => to_unsigned(808, 10), 487 => to_unsigned(17, 10), 488 => to_unsigned(933, 10), 489 => to_unsigned(130, 10), 490 => to_unsigned(956, 10), 491 => to_unsigned(377, 10), 492 => to_unsigned(106, 10), 493 => to_unsigned(707, 10), 494 => to_unsigned(252, 10), 495 => to_unsigned(428, 10), 496 => to_unsigned(637, 10), 497 => to_unsigned(554, 10), 498 => to_unsigned(972, 10), 499 => to_unsigned(216, 10), 500 => to_unsigned(636, 10), 501 => to_unsigned(505, 10), 502 => to_unsigned(878, 10), 503 => to_unsigned(845, 10), 504 => to_unsigned(515, 10), 505 => to_unsigned(937, 10), 506 => to_unsigned(82, 10), 507 => to_unsigned(500, 10), 508 => to_unsigned(341, 10), 509 => to_unsigned(231, 10), 510 => to_unsigned(613, 10), 511 => to_unsigned(187, 10), 512 => to_unsigned(475, 10), 513 => to_unsigned(909, 10), 514 => to_unsigned(279, 10), 515 => to_unsigned(372, 10), 516 => to_unsigned(846, 10), 517 => to_unsigned(81, 10), 518 => to_unsigned(600, 10), 519 => to_unsigned(866, 10), 520 => to_unsigned(14, 10), 521 => to_unsigned(644, 10), 522 => to_unsigned(120, 10), 523 => to_unsigned(542, 10), 524 => to_unsigned(92, 10), 525 => to_unsigned(181, 10), 526 => to_unsigned(738, 10), 527 => to_unsigned(849, 10), 528 => to_unsigned(289, 10), 529 => to_unsigned(970, 10), 530 => to_unsigned(34, 10), 531 => to_unsigned(958, 10), 532 => to_unsigned(697, 10), 533 => to_unsigned(661, 10), 534 => to_unsigned(593, 10), 535 => to_unsigned(964, 10), 536 => to_unsigned(526, 10), 537 => to_unsigned(864, 10), 538 => to_unsigned(996, 10), 539 => to_unsigned(747, 10), 540 => to_unsigned(24, 10), 541 => to_unsigned(352, 10), 542 => to_unsigned(970, 10), 543 => to_unsigned(958, 10), 544 => to_unsigned(255, 10), 545 => to_unsigned(766, 10), 546 => to_unsigned(772, 10), 547 => to_unsigned(366, 10), 548 => to_unsigned(256, 10), 549 => to_unsigned(80, 10), 550 => to_unsigned(290, 10), 551 => to_unsigned(337, 10), 552 => to_unsigned(99, 10), 553 => to_unsigned(121, 10), 554 => to_unsigned(584, 10), 555 => to_unsigned(93, 10), 556 => to_unsigned(909, 10), 557 => to_unsigned(539, 10), 558 => to_unsigned(585, 10), 559 => to_unsigned(945, 10), 560 => to_unsigned(693, 10), 561 => to_unsigned(165, 10), 562 => to_unsigned(181, 10), 563 => to_unsigned(1022, 10), 564 => to_unsigned(485, 10), 565 => to_unsigned(52, 10), 566 => to_unsigned(661, 10), 567 => to_unsigned(149, 10), 568 => to_unsigned(684, 10), 569 => to_unsigned(374, 10), 570 => to_unsigned(811, 10), 571 => to_unsigned(675, 10), 572 => to_unsigned(872, 10), 573 => to_unsigned(28, 10), 574 => to_unsigned(493, 10), 575 => to_unsigned(970, 10), 576 => to_unsigned(88, 10), 577 => to_unsigned(410, 10), 578 => to_unsigned(132, 10), 579 => to_unsigned(65, 10), 580 => to_unsigned(281, 10), 581 => to_unsigned(24, 10), 582 => to_unsigned(443, 10), 583 => to_unsigned(430, 10), 584 => to_unsigned(676, 10), 585 => to_unsigned(486, 10), 586 => to_unsigned(850, 10), 587 => to_unsigned(298, 10), 588 => to_unsigned(15, 10), 589 => to_unsigned(40, 10), 590 => to_unsigned(871, 10), 591 => to_unsigned(0, 10), 592 => to_unsigned(140, 10), 593 => to_unsigned(769, 10), 594 => to_unsigned(560, 10), 595 => to_unsigned(188, 10), 596 => to_unsigned(417, 10), 597 => to_unsigned(1022, 10), 598 => to_unsigned(203, 10), 599 => to_unsigned(125, 10), 600 => to_unsigned(935, 10), 601 => to_unsigned(587, 10), 602 => to_unsigned(235, 10), 603 => to_unsigned(706, 10), 604 => to_unsigned(411, 10), 605 => to_unsigned(724, 10), 606 => to_unsigned(384, 10), 607 => to_unsigned(665, 10), 608 => to_unsigned(292, 10), 609 => to_unsigned(993, 10), 610 => to_unsigned(256, 10), 611 => to_unsigned(226, 10), 612 => to_unsigned(336, 10), 613 => to_unsigned(856, 10), 614 => to_unsigned(696, 10), 615 => to_unsigned(535, 10), 616 => to_unsigned(853, 10), 617 => to_unsigned(409, 10), 618 => to_unsigned(173, 10), 619 => to_unsigned(144, 10), 620 => to_unsigned(988, 10), 621 => to_unsigned(59, 10), 622 => to_unsigned(915, 10), 623 => to_unsigned(581, 10), 624 => to_unsigned(524, 10), 625 => to_unsigned(770, 10), 626 => to_unsigned(683, 10), 627 => to_unsigned(561, 10), 628 => to_unsigned(610, 10), 629 => to_unsigned(63, 10), 630 => to_unsigned(248, 10), 631 => to_unsigned(982, 10), 632 => to_unsigned(674, 10), 633 => to_unsigned(389, 10), 634 => to_unsigned(287, 10), 635 => to_unsigned(567, 10), 636 => to_unsigned(936, 10), 637 => to_unsigned(83, 10), 638 => to_unsigned(806, 10), 639 => to_unsigned(504, 10), 640 => to_unsigned(698, 10), 641 => to_unsigned(824, 10), 642 => to_unsigned(932, 10), 643 => to_unsigned(575, 10), 644 => to_unsigned(87, 10), 645 => to_unsigned(472, 10), 646 => to_unsigned(1012, 10), 647 => to_unsigned(1022, 10), 648 => to_unsigned(935, 10), 649 => to_unsigned(585, 10), 650 => to_unsigned(1004, 10), 651 => to_unsigned(574, 10), 652 => to_unsigned(150, 10), 653 => to_unsigned(850, 10), 654 => to_unsigned(815, 10), 655 => to_unsigned(817, 10), 656 => to_unsigned(314, 10), 657 => to_unsigned(865, 10), 658 => to_unsigned(119, 10), 659 => to_unsigned(750, 10), 660 => to_unsigned(849, 10), 661 => to_unsigned(348, 10), 662 => to_unsigned(61, 10), 663 => to_unsigned(397, 10), 664 => to_unsigned(717, 10), 665 => to_unsigned(665, 10), 666 => to_unsigned(34, 10), 667 => to_unsigned(525, 10), 668 => to_unsigned(218, 10), 669 => to_unsigned(545, 10), 670 => to_unsigned(894, 10), 671 => to_unsigned(849, 10), 672 => to_unsigned(696, 10), 673 => to_unsigned(1016, 10), 674 => to_unsigned(241, 10), 675 => to_unsigned(473, 10), 676 => to_unsigned(373, 10), 677 => to_unsigned(1003, 10), 678 => to_unsigned(181, 10), 679 => to_unsigned(752, 10), 680 => to_unsigned(943, 10), 681 => to_unsigned(1005, 10), 682 => to_unsigned(564, 10), 683 => to_unsigned(362, 10), 684 => to_unsigned(100, 10), 685 => to_unsigned(477, 10), 686 => to_unsigned(838, 10), 687 => to_unsigned(488, 10), 688 => to_unsigned(720, 10), 689 => to_unsigned(157, 10), 690 => to_unsigned(451, 10), 691 => to_unsigned(654, 10), 692 => to_unsigned(403, 10), 693 => to_unsigned(988, 10), 694 => to_unsigned(366, 10), 695 => to_unsigned(895, 10), 696 => to_unsigned(291, 10), 697 => to_unsigned(931, 10), 698 => to_unsigned(225, 10), 699 => to_unsigned(447, 10), 700 => to_unsigned(1021, 10), 701 => to_unsigned(9, 10), 702 => to_unsigned(933, 10), 703 => to_unsigned(93, 10), 704 => to_unsigned(1011, 10), 705 => to_unsigned(834, 10), 706 => to_unsigned(1010, 10), 707 => to_unsigned(78, 10), 708 => to_unsigned(135, 10), 709 => to_unsigned(769, 10), 710 => to_unsigned(746, 10), 711 => to_unsigned(237, 10), 712 => to_unsigned(202, 10), 713 => to_unsigned(425, 10), 714 => to_unsigned(142, 10), 715 => to_unsigned(898, 10), 716 => to_unsigned(340, 10), 717 => to_unsigned(92, 10), 718 => to_unsigned(176, 10), 719 => to_unsigned(741, 10), 720 => to_unsigned(874, 10), 721 => to_unsigned(838, 10), 722 => to_unsigned(748, 10), 723 => to_unsigned(972, 10), 724 => to_unsigned(628, 10), 725 => to_unsigned(966, 10), 726 => to_unsigned(623, 10), 727 => to_unsigned(843, 10), 728 => to_unsigned(278, 10), 729 => to_unsigned(22, 10), 730 => to_unsigned(22, 10), 731 => to_unsigned(625, 10), 732 => to_unsigned(354, 10), 733 => to_unsigned(655, 10), 734 => to_unsigned(253, 10), 735 => to_unsigned(668, 10), 736 => to_unsigned(664, 10), 737 => to_unsigned(822, 10), 738 => to_unsigned(435, 10), 739 => to_unsigned(843, 10), 740 => to_unsigned(429, 10), 741 => to_unsigned(809, 10), 742 => to_unsigned(1021, 10), 743 => to_unsigned(970, 10), 744 => to_unsigned(775, 10), 745 => to_unsigned(1008, 10), 746 => to_unsigned(549, 10), 747 => to_unsigned(466, 10), 748 => to_unsigned(469, 10), 749 => to_unsigned(348, 10), 750 => to_unsigned(263, 10), 751 => to_unsigned(693, 10), 752 => to_unsigned(416, 10), 753 => to_unsigned(381, 10), 754 => to_unsigned(640, 10), 755 => to_unsigned(418, 10), 756 => to_unsigned(370, 10), 757 => to_unsigned(747, 10), 758 => to_unsigned(357, 10), 759 => to_unsigned(732, 10), 760 => to_unsigned(638, 10), 761 => to_unsigned(157, 10), 762 => to_unsigned(966, 10), 763 => to_unsigned(580, 10), 764 => to_unsigned(9, 10), 765 => to_unsigned(135, 10), 766 => to_unsigned(338, 10), 767 => to_unsigned(364, 10), 768 => to_unsigned(606, 10), 769 => to_unsigned(845, 10), 770 => to_unsigned(621, 10), 771 => to_unsigned(767, 10), 772 => to_unsigned(473, 10), 773 => to_unsigned(359, 10), 774 => to_unsigned(34, 10), 775 => to_unsigned(111, 10), 776 => to_unsigned(617, 10), 777 => to_unsigned(173, 10), 778 => to_unsigned(404, 10), 779 => to_unsigned(747, 10), 780 => to_unsigned(728, 10), 781 => to_unsigned(143, 10), 782 => to_unsigned(847, 10), 783 => to_unsigned(853, 10), 784 => to_unsigned(427, 10), 785 => to_unsigned(55, 10), 786 => to_unsigned(966, 10), 787 => to_unsigned(414, 10), 788 => to_unsigned(662, 10), 789 => to_unsigned(928, 10), 790 => to_unsigned(881, 10), 791 => to_unsigned(146, 10), 792 => to_unsigned(522, 10), 793 => to_unsigned(477, 10), 794 => to_unsigned(767, 10), 795 => to_unsigned(346, 10), 796 => to_unsigned(971, 10), 797 => to_unsigned(538, 10), 798 => to_unsigned(925, 10), 799 => to_unsigned(464, 10), 800 => to_unsigned(840, 10), 801 => to_unsigned(8, 10), 802 => to_unsigned(674, 10), 803 => to_unsigned(860, 10), 804 => to_unsigned(678, 10), 805 => to_unsigned(127, 10), 806 => to_unsigned(360, 10), 807 => to_unsigned(896, 10), 808 => to_unsigned(356, 10), 809 => to_unsigned(509, 10), 810 => to_unsigned(538, 10), 811 => to_unsigned(142, 10), 812 => to_unsigned(378, 10), 813 => to_unsigned(827, 10), 814 => to_unsigned(482, 10), 815 => to_unsigned(672, 10), 816 => to_unsigned(51, 10), 817 => to_unsigned(231, 10), 818 => to_unsigned(612, 10), 819 => to_unsigned(724, 10), 820 => to_unsigned(697, 10), 821 => to_unsigned(510, 10), 822 => to_unsigned(3, 10), 823 => to_unsigned(636, 10), 824 => to_unsigned(287, 10), 825 => to_unsigned(654, 10), 826 => to_unsigned(257, 10), 827 => to_unsigned(991, 10), 828 => to_unsigned(544, 10), 829 => to_unsigned(380, 10), 830 => to_unsigned(758, 10), 831 => to_unsigned(625, 10), 832 => to_unsigned(993, 10), 833 => to_unsigned(139, 10), 834 => to_unsigned(970, 10), 835 => to_unsigned(504, 10), 836 => to_unsigned(498, 10), 837 => to_unsigned(305, 10), 838 => to_unsigned(396, 10), 839 => to_unsigned(834, 10), 840 => to_unsigned(773, 10), 841 => to_unsigned(143, 10), 842 => to_unsigned(535, 10), 843 => to_unsigned(381, 10), 844 => to_unsigned(306, 10), 845 => to_unsigned(924, 10), 846 => to_unsigned(270, 10), 847 => to_unsigned(234, 10), 848 => to_unsigned(437, 10), 849 => to_unsigned(319, 10), 850 => to_unsigned(660, 10), 851 => to_unsigned(104, 10), 852 => to_unsigned(254, 10), 853 => to_unsigned(389, 10), 854 => to_unsigned(51, 10), 855 => to_unsigned(532, 10), 856 => to_unsigned(484, 10), 857 => to_unsigned(222, 10), 858 => to_unsigned(828, 10), 859 => to_unsigned(51, 10), 860 => to_unsigned(833, 10), 861 => to_unsigned(421, 10), 862 => to_unsigned(726, 10), 863 => to_unsigned(184, 10), 864 => to_unsigned(918, 10), 865 => to_unsigned(293, 10), 866 => to_unsigned(975, 10), 867 => to_unsigned(276, 10), 868 => to_unsigned(762, 10), 869 => to_unsigned(951, 10), 870 => to_unsigned(304, 10), 871 => to_unsigned(943, 10), 872 => to_unsigned(748, 10), 873 => to_unsigned(297, 10), 874 => to_unsigned(74, 10), 875 => to_unsigned(228, 10), 876 => to_unsigned(739, 10), 877 => to_unsigned(170, 10), 878 => to_unsigned(14, 10), 879 => to_unsigned(286, 10), 880 => to_unsigned(175, 10), 881 => to_unsigned(987, 10), 882 => to_unsigned(192, 10), 883 => to_unsigned(866, 10), 884 => to_unsigned(5, 10), 885 => to_unsigned(826, 10), 886 => to_unsigned(691, 10), 887 => to_unsigned(718, 10), 888 => to_unsigned(736, 10), 889 => to_unsigned(256, 10), 890 => to_unsigned(67, 10), 891 => to_unsigned(76, 10), 892 => to_unsigned(601, 10), 893 => to_unsigned(159, 10), 894 => to_unsigned(259, 10), 895 => to_unsigned(747, 10), 896 => to_unsigned(327, 10), 897 => to_unsigned(860, 10), 898 => to_unsigned(1007, 10), 899 => to_unsigned(436, 10), 900 => to_unsigned(141, 10), 901 => to_unsigned(687, 10), 902 => to_unsigned(13, 10), 903 => to_unsigned(954, 10), 904 => to_unsigned(446, 10), 905 => to_unsigned(487, 10), 906 => to_unsigned(142, 10), 907 => to_unsigned(730, 10), 908 => to_unsigned(936, 10), 909 => to_unsigned(188, 10), 910 => to_unsigned(150, 10), 911 => to_unsigned(494, 10), 912 => to_unsigned(960, 10), 913 => to_unsigned(110, 10), 914 => to_unsigned(155, 10), 915 => to_unsigned(752, 10), 916 => to_unsigned(899, 10), 917 => to_unsigned(987, 10), 918 => to_unsigned(831, 10), 919 => to_unsigned(540, 10), 920 => to_unsigned(16, 10), 921 => to_unsigned(412, 10), 922 => to_unsigned(53, 10), 923 => to_unsigned(627, 10), 924 => to_unsigned(661, 10), 925 => to_unsigned(602, 10), 926 => to_unsigned(105, 10), 927 => to_unsigned(953, 10), 928 => to_unsigned(452, 10), 929 => to_unsigned(171, 10), 930 => to_unsigned(191, 10), 931 => to_unsigned(844, 10), 932 => to_unsigned(436, 10), 933 => to_unsigned(62, 10), 934 => to_unsigned(983, 10), 935 => to_unsigned(85, 10), 936 => to_unsigned(162, 10), 937 => to_unsigned(646, 10), 938 => to_unsigned(340, 10), 939 => to_unsigned(438, 10), 940 => to_unsigned(568, 10), 941 => to_unsigned(805, 10), 942 => to_unsigned(271, 10), 943 => to_unsigned(382, 10), 944 => to_unsigned(782, 10), 945 => to_unsigned(957, 10), 946 => to_unsigned(354, 10), 947 => to_unsigned(281, 10), 948 => to_unsigned(908, 10), 949 => to_unsigned(452, 10), 950 => to_unsigned(105, 10), 951 => to_unsigned(442, 10), 952 => to_unsigned(653, 10), 953 => to_unsigned(698, 10), 954 => to_unsigned(683, 10), 955 => to_unsigned(672, 10), 956 => to_unsigned(82, 10), 957 => to_unsigned(334, 10), 958 => to_unsigned(806, 10), 959 => to_unsigned(893, 10), 960 => to_unsigned(830, 10), 961 => to_unsigned(484, 10), 962 => to_unsigned(680, 10), 963 => to_unsigned(986, 10), 964 => to_unsigned(734, 10), 965 => to_unsigned(807, 10), 966 => to_unsigned(955, 10), 967 => to_unsigned(0, 10), 968 => to_unsigned(161, 10), 969 => to_unsigned(180, 10), 970 => to_unsigned(728, 10), 971 => to_unsigned(720, 10), 972 => to_unsigned(264, 10), 973 => to_unsigned(96, 10), 974 => to_unsigned(705, 10), 975 => to_unsigned(272, 10), 976 => to_unsigned(407, 10), 977 => to_unsigned(861, 10), 978 => to_unsigned(263, 10), 979 => to_unsigned(605, 10), 980 => to_unsigned(165, 10), 981 => to_unsigned(641, 10), 982 => to_unsigned(688, 10), 983 => to_unsigned(312, 10), 984 => to_unsigned(681, 10), 985 => to_unsigned(622, 10), 986 => to_unsigned(871, 10), 987 => to_unsigned(16, 10), 988 => to_unsigned(810, 10), 989 => to_unsigned(697, 10), 990 => to_unsigned(637, 10), 991 => to_unsigned(676, 10), 992 => to_unsigned(794, 10), 993 => to_unsigned(288, 10), 994 => to_unsigned(1008, 10), 995 => to_unsigned(20, 10), 996 => to_unsigned(682, 10), 997 => to_unsigned(701, 10), 998 => to_unsigned(137, 10), 999 => to_unsigned(786, 10), 1000 => to_unsigned(932, 10), 1001 => to_unsigned(849, 10), 1002 => to_unsigned(118, 10), 1003 => to_unsigned(889, 10), 1004 => to_unsigned(19, 10), 1005 => to_unsigned(456, 10), 1006 => to_unsigned(190, 10), 1007 => to_unsigned(281, 10), 1008 => to_unsigned(409, 10), 1009 => to_unsigned(651, 10), 1010 => to_unsigned(803, 10), 1011 => to_unsigned(945, 10), 1012 => to_unsigned(868, 10), 1013 => to_unsigned(981, 10), 1014 => to_unsigned(381, 10), 1015 => to_unsigned(399, 10), 1016 => to_unsigned(179, 10), 1017 => to_unsigned(986, 10), 1018 => to_unsigned(284, 10), 1019 => to_unsigned(738, 10), 1020 => to_unsigned(914, 10), 1021 => to_unsigned(606, 10), 1022 => to_unsigned(92, 10), 1023 => to_unsigned(1001, 10), 1024 => to_unsigned(408, 10), 1025 => to_unsigned(837, 10), 1026 => to_unsigned(87, 10), 1027 => to_unsigned(346, 10), 1028 => to_unsigned(276, 10), 1029 => to_unsigned(967, 10), 1030 => to_unsigned(578, 10), 1031 => to_unsigned(16, 10), 1032 => to_unsigned(755, 10), 1033 => to_unsigned(347, 10), 1034 => to_unsigned(565, 10), 1035 => to_unsigned(413, 10), 1036 => to_unsigned(199, 10), 1037 => to_unsigned(739, 10), 1038 => to_unsigned(165, 10), 1039 => to_unsigned(38, 10), 1040 => to_unsigned(650, 10), 1041 => to_unsigned(546, 10), 1042 => to_unsigned(340, 10), 1043 => to_unsigned(782, 10), 1044 => to_unsigned(542, 10), 1045 => to_unsigned(54, 10), 1046 => to_unsigned(601, 10), 1047 => to_unsigned(166, 10), 1048 => to_unsigned(736, 10), 1049 => to_unsigned(443, 10), 1050 => to_unsigned(865, 10), 1051 => to_unsigned(440, 10), 1052 => to_unsigned(275, 10), 1053 => to_unsigned(851, 10), 1054 => to_unsigned(413, 10), 1055 => to_unsigned(229, 10), 1056 => to_unsigned(894, 10), 1057 => to_unsigned(897, 10), 1058 => to_unsigned(254, 10), 1059 => to_unsigned(565, 10), 1060 => to_unsigned(200, 10), 1061 => to_unsigned(644, 10), 1062 => to_unsigned(165, 10), 1063 => to_unsigned(435, 10), 1064 => to_unsigned(870, 10), 1065 => to_unsigned(601, 10), 1066 => to_unsigned(473, 10), 1067 => to_unsigned(758, 10), 1068 => to_unsigned(37, 10), 1069 => to_unsigned(316, 10), 1070 => to_unsigned(742, 10), 1071 => to_unsigned(628, 10), 1072 => to_unsigned(279, 10), 1073 => to_unsigned(633, 10), 1074 => to_unsigned(1022, 10), 1075 => to_unsigned(369, 10), 1076 => to_unsigned(439, 10), 1077 => to_unsigned(333, 10), 1078 => to_unsigned(370, 10), 1079 => to_unsigned(160, 10), 1080 => to_unsigned(532, 10), 1081 => to_unsigned(892, 10), 1082 => to_unsigned(284, 10), 1083 => to_unsigned(625, 10), 1084 => to_unsigned(421, 10), 1085 => to_unsigned(966, 10), 1086 => to_unsigned(755, 10), 1087 => to_unsigned(576, 10), 1088 => to_unsigned(485, 10), 1089 => to_unsigned(849, 10), 1090 => to_unsigned(510, 10), 1091 => to_unsigned(592, 10), 1092 => to_unsigned(725, 10), 1093 => to_unsigned(329, 10), 1094 => to_unsigned(116, 10), 1095 => to_unsigned(619, 10), 1096 => to_unsigned(322, 10), 1097 => to_unsigned(641, 10), 1098 => to_unsigned(129, 10), 1099 => to_unsigned(871, 10), 1100 => to_unsigned(726, 10), 1101 => to_unsigned(404, 10), 1102 => to_unsigned(126, 10), 1103 => to_unsigned(330, 10), 1104 => to_unsigned(1004, 10), 1105 => to_unsigned(905, 10), 1106 => to_unsigned(644, 10), 1107 => to_unsigned(557, 10), 1108 => to_unsigned(311, 10), 1109 => to_unsigned(599, 10), 1110 => to_unsigned(63, 10), 1111 => to_unsigned(624, 10), 1112 => to_unsigned(328, 10), 1113 => to_unsigned(887, 10), 1114 => to_unsigned(912, 10), 1115 => to_unsigned(290, 10), 1116 => to_unsigned(813, 10), 1117 => to_unsigned(926, 10), 1118 => to_unsigned(904, 10), 1119 => to_unsigned(163, 10), 1120 => to_unsigned(186, 10), 1121 => to_unsigned(700, 10), 1122 => to_unsigned(988, 10), 1123 => to_unsigned(182, 10), 1124 => to_unsigned(535, 10), 1125 => to_unsigned(901, 10), 1126 => to_unsigned(867, 10), 1127 => to_unsigned(632, 10), 1128 => to_unsigned(92, 10), 1129 => to_unsigned(972, 10), 1130 => to_unsigned(548, 10), 1131 => to_unsigned(90, 10), 1132 => to_unsigned(660, 10), 1133 => to_unsigned(483, 10), 1134 => to_unsigned(215, 10), 1135 => to_unsigned(253, 10), 1136 => to_unsigned(834, 10), 1137 => to_unsigned(714, 10), 1138 => to_unsigned(900, 10), 1139 => to_unsigned(125, 10), 1140 => to_unsigned(241, 10), 1141 => to_unsigned(483, 10), 1142 => to_unsigned(291, 10), 1143 => to_unsigned(563, 10), 1144 => to_unsigned(274, 10), 1145 => to_unsigned(274, 10), 1146 => to_unsigned(794, 10), 1147 => to_unsigned(255, 10), 1148 => to_unsigned(570, 10), 1149 => to_unsigned(490, 10), 1150 => to_unsigned(801, 10), 1151 => to_unsigned(167, 10), 1152 => to_unsigned(851, 10), 1153 => to_unsigned(851, 10), 1154 => to_unsigned(516, 10), 1155 => to_unsigned(910, 10), 1156 => to_unsigned(203, 10), 1157 => to_unsigned(613, 10), 1158 => to_unsigned(85, 10), 1159 => to_unsigned(5, 10), 1160 => to_unsigned(1001, 10), 1161 => to_unsigned(654, 10), 1162 => to_unsigned(966, 10), 1163 => to_unsigned(78, 10), 1164 => to_unsigned(390, 10), 1165 => to_unsigned(586, 10), 1166 => to_unsigned(145, 10), 1167 => to_unsigned(109, 10), 1168 => to_unsigned(215, 10), 1169 => to_unsigned(194, 10), 1170 => to_unsigned(726, 10), 1171 => to_unsigned(828, 10), 1172 => to_unsigned(146, 10), 1173 => to_unsigned(208, 10), 1174 => to_unsigned(119, 10), 1175 => to_unsigned(48, 10), 1176 => to_unsigned(322, 10), 1177 => to_unsigned(840, 10), 1178 => to_unsigned(213, 10), 1179 => to_unsigned(611, 10), 1180 => to_unsigned(907, 10), 1181 => to_unsigned(809, 10), 1182 => to_unsigned(591, 10), 1183 => to_unsigned(179, 10), 1184 => to_unsigned(916, 10), 1185 => to_unsigned(116, 10), 1186 => to_unsigned(86, 10), 1187 => to_unsigned(997, 10), 1188 => to_unsigned(345, 10), 1189 => to_unsigned(839, 10), 1190 => to_unsigned(728, 10), 1191 => to_unsigned(876, 10), 1192 => to_unsigned(299, 10), 1193 => to_unsigned(527, 10), 1194 => to_unsigned(239, 10), 1195 => to_unsigned(331, 10), 1196 => to_unsigned(535, 10), 1197 => to_unsigned(682, 10), 1198 => to_unsigned(89, 10), 1199 => to_unsigned(96, 10), 1200 => to_unsigned(885, 10), 1201 => to_unsigned(983, 10), 1202 => to_unsigned(231, 10), 1203 => to_unsigned(494, 10), 1204 => to_unsigned(146, 10), 1205 => to_unsigned(493, 10), 1206 => to_unsigned(429, 10), 1207 => to_unsigned(419, 10), 1208 => to_unsigned(929, 10), 1209 => to_unsigned(305, 10), 1210 => to_unsigned(812, 10), 1211 => to_unsigned(203, 10), 1212 => to_unsigned(445, 10), 1213 => to_unsigned(555, 10), 1214 => to_unsigned(290, 10), 1215 => to_unsigned(539, 10), 1216 => to_unsigned(910, 10), 1217 => to_unsigned(899, 10), 1218 => to_unsigned(840, 10), 1219 => to_unsigned(961, 10), 1220 => to_unsigned(264, 10), 1221 => to_unsigned(847, 10), 1222 => to_unsigned(77, 10), 1223 => to_unsigned(566, 10), 1224 => to_unsigned(1019, 10), 1225 => to_unsigned(301, 10), 1226 => to_unsigned(962, 10), 1227 => to_unsigned(52, 10), 1228 => to_unsigned(968, 10), 1229 => to_unsigned(637, 10), 1230 => to_unsigned(1015, 10), 1231 => to_unsigned(744, 10), 1232 => to_unsigned(698, 10), 1233 => to_unsigned(211, 10), 1234 => to_unsigned(396, 10), 1235 => to_unsigned(632, 10), 1236 => to_unsigned(402, 10), 1237 => to_unsigned(254, 10), 1238 => to_unsigned(304, 10), 1239 => to_unsigned(859, 10), 1240 => to_unsigned(475, 10), 1241 => to_unsigned(21, 10), 1242 => to_unsigned(144, 10), 1243 => to_unsigned(678, 10), 1244 => to_unsigned(196, 10), 1245 => to_unsigned(863, 10), 1246 => to_unsigned(791, 10), 1247 => to_unsigned(685, 10), 1248 => to_unsigned(227, 10), 1249 => to_unsigned(911, 10), 1250 => to_unsigned(529, 10), 1251 => to_unsigned(108, 10), 1252 => to_unsigned(459, 10), 1253 => to_unsigned(892, 10), 1254 => to_unsigned(801, 10), 1255 => to_unsigned(405, 10), 1256 => to_unsigned(24, 10), 1257 => to_unsigned(334, 10), 1258 => to_unsigned(465, 10), 1259 => to_unsigned(228, 10), 1260 => to_unsigned(669, 10), 1261 => to_unsigned(927, 10), 1262 => to_unsigned(493, 10), 1263 => to_unsigned(618, 10), 1264 => to_unsigned(965, 10), 1265 => to_unsigned(485, 10), 1266 => to_unsigned(898, 10), 1267 => to_unsigned(820, 10), 1268 => to_unsigned(285, 10), 1269 => to_unsigned(630, 10), 1270 => to_unsigned(799, 10), 1271 => to_unsigned(482, 10), 1272 => to_unsigned(67, 10), 1273 => to_unsigned(630, 10), 1274 => to_unsigned(652, 10), 1275 => to_unsigned(227, 10), 1276 => to_unsigned(660, 10), 1277 => to_unsigned(550, 10), 1278 => to_unsigned(817, 10), 1279 => to_unsigned(374, 10), 1280 => to_unsigned(812, 10), 1281 => to_unsigned(796, 10), 1282 => to_unsigned(648, 10), 1283 => to_unsigned(210, 10), 1284 => to_unsigned(138, 10), 1285 => to_unsigned(81, 10), 1286 => to_unsigned(929, 10), 1287 => to_unsigned(745, 10), 1288 => to_unsigned(344, 10), 1289 => to_unsigned(57, 10), 1290 => to_unsigned(566, 10), 1291 => to_unsigned(140, 10), 1292 => to_unsigned(205, 10), 1293 => to_unsigned(2, 10), 1294 => to_unsigned(91, 10), 1295 => to_unsigned(28, 10), 1296 => to_unsigned(788, 10), 1297 => to_unsigned(192, 10), 1298 => to_unsigned(552, 10), 1299 => to_unsigned(744, 10), 1300 => to_unsigned(234, 10), 1301 => to_unsigned(21, 10), 1302 => to_unsigned(373, 10), 1303 => to_unsigned(535, 10), 1304 => to_unsigned(81, 10), 1305 => to_unsigned(669, 10), 1306 => to_unsigned(738, 10), 1307 => to_unsigned(378, 10), 1308 => to_unsigned(490, 10), 1309 => to_unsigned(426, 10), 1310 => to_unsigned(155, 10), 1311 => to_unsigned(678, 10), 1312 => to_unsigned(246, 10), 1313 => to_unsigned(887, 10), 1314 => to_unsigned(521, 10), 1315 => to_unsigned(826, 10), 1316 => to_unsigned(765, 10), 1317 => to_unsigned(498, 10), 1318 => to_unsigned(290, 10), 1319 => to_unsigned(762, 10), 1320 => to_unsigned(55, 10), 1321 => to_unsigned(933, 10), 1322 => to_unsigned(687, 10), 1323 => to_unsigned(729, 10), 1324 => to_unsigned(661, 10), 1325 => to_unsigned(1006, 10), 1326 => to_unsigned(941, 10), 1327 => to_unsigned(31, 10), 1328 => to_unsigned(523, 10), 1329 => to_unsigned(653, 10), 1330 => to_unsigned(692, 10), 1331 => to_unsigned(527, 10), 1332 => to_unsigned(20, 10), 1333 => to_unsigned(905, 10), 1334 => to_unsigned(872, 10), 1335 => to_unsigned(144, 10), 1336 => to_unsigned(550, 10), 1337 => to_unsigned(936, 10), 1338 => to_unsigned(46, 10), 1339 => to_unsigned(507, 10), 1340 => to_unsigned(83, 10), 1341 => to_unsigned(376, 10), 1342 => to_unsigned(912, 10), 1343 => to_unsigned(69, 10), 1344 => to_unsigned(786, 10), 1345 => to_unsigned(90, 10), 1346 => to_unsigned(231, 10), 1347 => to_unsigned(608, 10), 1348 => to_unsigned(555, 10), 1349 => to_unsigned(1003, 10), 1350 => to_unsigned(680, 10), 1351 => to_unsigned(569, 10), 1352 => to_unsigned(586, 10), 1353 => to_unsigned(735, 10), 1354 => to_unsigned(838, 10), 1355 => to_unsigned(294, 10), 1356 => to_unsigned(665, 10), 1357 => to_unsigned(635, 10), 1358 => to_unsigned(73, 10), 1359 => to_unsigned(828, 10), 1360 => to_unsigned(100, 10), 1361 => to_unsigned(71, 10), 1362 => to_unsigned(659, 10), 1363 => to_unsigned(773, 10), 1364 => to_unsigned(774, 10), 1365 => to_unsigned(155, 10), 1366 => to_unsigned(409, 10), 1367 => to_unsigned(752, 10), 1368 => to_unsigned(339, 10), 1369 => to_unsigned(167, 10), 1370 => to_unsigned(506, 10), 1371 => to_unsigned(917, 10), 1372 => to_unsigned(760, 10), 1373 => to_unsigned(486, 10), 1374 => to_unsigned(332, 10), 1375 => to_unsigned(408, 10), 1376 => to_unsigned(223, 10), 1377 => to_unsigned(241, 10), 1378 => to_unsigned(91, 10), 1379 => to_unsigned(122, 10), 1380 => to_unsigned(62, 10), 1381 => to_unsigned(561, 10), 1382 => to_unsigned(819, 10), 1383 => to_unsigned(77, 10), 1384 => to_unsigned(781, 10), 1385 => to_unsigned(576, 10), 1386 => to_unsigned(844, 10), 1387 => to_unsigned(659, 10), 1388 => to_unsigned(695, 10), 1389 => to_unsigned(75, 10), 1390 => to_unsigned(316, 10), 1391 => to_unsigned(201, 10), 1392 => to_unsigned(91, 10), 1393 => to_unsigned(1000, 10), 1394 => to_unsigned(498, 10), 1395 => to_unsigned(935, 10), 1396 => to_unsigned(55, 10), 1397 => to_unsigned(867, 10), 1398 => to_unsigned(423, 10), 1399 => to_unsigned(826, 10), 1400 => to_unsigned(943, 10), 1401 => to_unsigned(1015, 10), 1402 => to_unsigned(172, 10), 1403 => to_unsigned(635, 10), 1404 => to_unsigned(15, 10), 1405 => to_unsigned(87, 10), 1406 => to_unsigned(863, 10), 1407 => to_unsigned(683, 10), 1408 => to_unsigned(466, 10), 1409 => to_unsigned(566, 10), 1410 => to_unsigned(268, 10), 1411 => to_unsigned(240, 10), 1412 => to_unsigned(767, 10), 1413 => to_unsigned(3, 10), 1414 => to_unsigned(872, 10), 1415 => to_unsigned(593, 10), 1416 => to_unsigned(779, 10), 1417 => to_unsigned(358, 10), 1418 => to_unsigned(511, 10), 1419 => to_unsigned(866, 10), 1420 => to_unsigned(316, 10), 1421 => to_unsigned(288, 10), 1422 => to_unsigned(385, 10), 1423 => to_unsigned(63, 10), 1424 => to_unsigned(811, 10), 1425 => to_unsigned(23, 10), 1426 => to_unsigned(513, 10), 1427 => to_unsigned(830, 10), 1428 => to_unsigned(248, 10), 1429 => to_unsigned(567, 10), 1430 => to_unsigned(306, 10), 1431 => to_unsigned(418, 10), 1432 => to_unsigned(35, 10), 1433 => to_unsigned(832, 10), 1434 => to_unsigned(795, 10), 1435 => to_unsigned(220, 10), 1436 => to_unsigned(654, 10), 1437 => to_unsigned(94, 10), 1438 => to_unsigned(649, 10), 1439 => to_unsigned(907, 10), 1440 => to_unsigned(985, 10), 1441 => to_unsigned(87, 10), 1442 => to_unsigned(884, 10), 1443 => to_unsigned(347, 10), 1444 => to_unsigned(286, 10), 1445 => to_unsigned(639, 10), 1446 => to_unsigned(607, 10), 1447 => to_unsigned(845, 10), 1448 => to_unsigned(968, 10), 1449 => to_unsigned(658, 10), 1450 => to_unsigned(656, 10), 1451 => to_unsigned(68, 10), 1452 => to_unsigned(398, 10), 1453 => to_unsigned(1015, 10), 1454 => to_unsigned(651, 10), 1455 => to_unsigned(983, 10), 1456 => to_unsigned(257, 10), 1457 => to_unsigned(1004, 10), 1458 => to_unsigned(571, 10), 1459 => to_unsigned(466, 10), 1460 => to_unsigned(839, 10), 1461 => to_unsigned(922, 10), 1462 => to_unsigned(373, 10), 1463 => to_unsigned(716, 10), 1464 => to_unsigned(809, 10), 1465 => to_unsigned(297, 10), 1466 => to_unsigned(688, 10), 1467 => to_unsigned(210, 10), 1468 => to_unsigned(580, 10), 1469 => to_unsigned(835, 10), 1470 => to_unsigned(873, 10), 1471 => to_unsigned(386, 10), 1472 => to_unsigned(534, 10), 1473 => to_unsigned(509, 10), 1474 => to_unsigned(10, 10), 1475 => to_unsigned(684, 10), 1476 => to_unsigned(104, 10), 1477 => to_unsigned(134, 10), 1478 => to_unsigned(117, 10), 1479 => to_unsigned(101, 10), 1480 => to_unsigned(677, 10), 1481 => to_unsigned(655, 10), 1482 => to_unsigned(849, 10), 1483 => to_unsigned(102, 10), 1484 => to_unsigned(999, 10), 1485 => to_unsigned(577, 10), 1486 => to_unsigned(999, 10), 1487 => to_unsigned(261, 10), 1488 => to_unsigned(326, 10), 1489 => to_unsigned(590, 10), 1490 => to_unsigned(154, 10), 1491 => to_unsigned(904, 10), 1492 => to_unsigned(456, 10), 1493 => to_unsigned(77, 10), 1494 => to_unsigned(792, 10), 1495 => to_unsigned(863, 10), 1496 => to_unsigned(304, 10), 1497 => to_unsigned(853, 10), 1498 => to_unsigned(117, 10), 1499 => to_unsigned(107, 10), 1500 => to_unsigned(576, 10), 1501 => to_unsigned(78, 10), 1502 => to_unsigned(732, 10), 1503 => to_unsigned(288, 10), 1504 => to_unsigned(254, 10), 1505 => to_unsigned(315, 10), 1506 => to_unsigned(449, 10), 1507 => to_unsigned(503, 10), 1508 => to_unsigned(758, 10), 1509 => to_unsigned(671, 10), 1510 => to_unsigned(597, 10), 1511 => to_unsigned(714, 10), 1512 => to_unsigned(831, 10), 1513 => to_unsigned(408, 10), 1514 => to_unsigned(655, 10), 1515 => to_unsigned(64, 10), 1516 => to_unsigned(633, 10), 1517 => to_unsigned(407, 10), 1518 => to_unsigned(314, 10), 1519 => to_unsigned(327, 10), 1520 => to_unsigned(358, 10), 1521 => to_unsigned(347, 10), 1522 => to_unsigned(83, 10), 1523 => to_unsigned(680, 10), 1524 => to_unsigned(681, 10), 1525 => to_unsigned(763, 10), 1526 => to_unsigned(466, 10), 1527 => to_unsigned(824, 10), 1528 => to_unsigned(1021, 10), 1529 => to_unsigned(406, 10), 1530 => to_unsigned(43, 10), 1531 => to_unsigned(444, 10), 1532 => to_unsigned(782, 10), 1533 => to_unsigned(165, 10), 1534 => to_unsigned(720, 10), 1535 => to_unsigned(96, 10), 1536 => to_unsigned(231, 10), 1537 => to_unsigned(680, 10), 1538 => to_unsigned(417, 10), 1539 => to_unsigned(800, 10), 1540 => to_unsigned(443, 10), 1541 => to_unsigned(863, 10), 1542 => to_unsigned(1004, 10), 1543 => to_unsigned(95, 10), 1544 => to_unsigned(221, 10), 1545 => to_unsigned(284, 10), 1546 => to_unsigned(687, 10), 1547 => to_unsigned(713, 10), 1548 => to_unsigned(702, 10), 1549 => to_unsigned(243, 10), 1550 => to_unsigned(25, 10), 1551 => to_unsigned(87, 10), 1552 => to_unsigned(673, 10), 1553 => to_unsigned(496, 10), 1554 => to_unsigned(162, 10), 1555 => to_unsigned(165, 10), 1556 => to_unsigned(985, 10), 1557 => to_unsigned(401, 10), 1558 => to_unsigned(247, 10), 1559 => to_unsigned(620, 10), 1560 => to_unsigned(114, 10), 1561 => to_unsigned(231, 10), 1562 => to_unsigned(922, 10), 1563 => to_unsigned(332, 10), 1564 => to_unsigned(973, 10), 1565 => to_unsigned(230, 10), 1566 => to_unsigned(348, 10), 1567 => to_unsigned(361, 10), 1568 => to_unsigned(306, 10), 1569 => to_unsigned(945, 10), 1570 => to_unsigned(664, 10), 1571 => to_unsigned(963, 10), 1572 => to_unsigned(664, 10), 1573 => to_unsigned(285, 10), 1574 => to_unsigned(452, 10), 1575 => to_unsigned(969, 10), 1576 => to_unsigned(324, 10), 1577 => to_unsigned(816, 10), 1578 => to_unsigned(360, 10), 1579 => to_unsigned(293, 10), 1580 => to_unsigned(762, 10), 1581 => to_unsigned(706, 10), 1582 => to_unsigned(86, 10), 1583 => to_unsigned(55, 10), 1584 => to_unsigned(200, 10), 1585 => to_unsigned(45, 10), 1586 => to_unsigned(320, 10), 1587 => to_unsigned(59, 10), 1588 => to_unsigned(453, 10), 1589 => to_unsigned(268, 10), 1590 => to_unsigned(955, 10), 1591 => to_unsigned(530, 10), 1592 => to_unsigned(842, 10), 1593 => to_unsigned(795, 10), 1594 => to_unsigned(386, 10), 1595 => to_unsigned(627, 10), 1596 => to_unsigned(270, 10), 1597 => to_unsigned(879, 10), 1598 => to_unsigned(369, 10), 1599 => to_unsigned(992, 10), 1600 => to_unsigned(390, 10), 1601 => to_unsigned(572, 10), 1602 => to_unsigned(1020, 10), 1603 => to_unsigned(132, 10), 1604 => to_unsigned(194, 10), 1605 => to_unsigned(706, 10), 1606 => to_unsigned(557, 10), 1607 => to_unsigned(217, 10), 1608 => to_unsigned(73, 10), 1609 => to_unsigned(506, 10), 1610 => to_unsigned(991, 10), 1611 => to_unsigned(638, 10), 1612 => to_unsigned(792, 10), 1613 => to_unsigned(335, 10), 1614 => to_unsigned(530, 10), 1615 => to_unsigned(270, 10), 1616 => to_unsigned(75, 10), 1617 => to_unsigned(170, 10), 1618 => to_unsigned(751, 10), 1619 => to_unsigned(416, 10), 1620 => to_unsigned(77, 10), 1621 => to_unsigned(910, 10), 1622 => to_unsigned(490, 10), 1623 => to_unsigned(18, 10), 1624 => to_unsigned(286, 10), 1625 => to_unsigned(842, 10), 1626 => to_unsigned(951, 10), 1627 => to_unsigned(633, 10), 1628 => to_unsigned(738, 10), 1629 => to_unsigned(685, 10), 1630 => to_unsigned(227, 10), 1631 => to_unsigned(811, 10), 1632 => to_unsigned(878, 10), 1633 => to_unsigned(85, 10), 1634 => to_unsigned(596, 10), 1635 => to_unsigned(534, 10), 1636 => to_unsigned(463, 10), 1637 => to_unsigned(417, 10), 1638 => to_unsigned(184, 10), 1639 => to_unsigned(987, 10), 1640 => to_unsigned(865, 10), 1641 => to_unsigned(992, 10), 1642 => to_unsigned(859, 10), 1643 => to_unsigned(608, 10), 1644 => to_unsigned(497, 10), 1645 => to_unsigned(476, 10), 1646 => to_unsigned(381, 10), 1647 => to_unsigned(773, 10), 1648 => to_unsigned(532, 10), 1649 => to_unsigned(381, 10), 1650 => to_unsigned(649, 10), 1651 => to_unsigned(613, 10), 1652 => to_unsigned(550, 10), 1653 => to_unsigned(785, 10), 1654 => to_unsigned(262, 10), 1655 => to_unsigned(452, 10), 1656 => to_unsigned(202, 10), 1657 => to_unsigned(94, 10), 1658 => to_unsigned(2, 10), 1659 => to_unsigned(878, 10), 1660 => to_unsigned(402, 10), 1661 => to_unsigned(56, 10), 1662 => to_unsigned(810, 10), 1663 => to_unsigned(543, 10), 1664 => to_unsigned(285, 10), 1665 => to_unsigned(564, 10), 1666 => to_unsigned(50, 10), 1667 => to_unsigned(955, 10), 1668 => to_unsigned(348, 10), 1669 => to_unsigned(356, 10), 1670 => to_unsigned(818, 10), 1671 => to_unsigned(341, 10), 1672 => to_unsigned(60, 10), 1673 => to_unsigned(675, 10), 1674 => to_unsigned(336, 10), 1675 => to_unsigned(745, 10), 1676 => to_unsigned(273, 10), 1677 => to_unsigned(795, 10), 1678 => to_unsigned(723, 10), 1679 => to_unsigned(77, 10), 1680 => to_unsigned(673, 10), 1681 => to_unsigned(729, 10), 1682 => to_unsigned(653, 10), 1683 => to_unsigned(892, 10), 1684 => to_unsigned(5, 10), 1685 => to_unsigned(681, 10), 1686 => to_unsigned(565, 10), 1687 => to_unsigned(600, 10), 1688 => to_unsigned(108, 10), 1689 => to_unsigned(258, 10), 1690 => to_unsigned(713, 10), 1691 => to_unsigned(975, 10), 1692 => to_unsigned(831, 10), 1693 => to_unsigned(771, 10), 1694 => to_unsigned(61, 10), 1695 => to_unsigned(192, 10), 1696 => to_unsigned(44, 10), 1697 => to_unsigned(848, 10), 1698 => to_unsigned(610, 10), 1699 => to_unsigned(670, 10), 1700 => to_unsigned(340, 10), 1701 => to_unsigned(614, 10), 1702 => to_unsigned(177, 10), 1703 => to_unsigned(218, 10), 1704 => to_unsigned(606, 10), 1705 => to_unsigned(598, 10), 1706 => to_unsigned(206, 10), 1707 => to_unsigned(951, 10), 1708 => to_unsigned(547, 10), 1709 => to_unsigned(576, 10), 1710 => to_unsigned(896, 10), 1711 => to_unsigned(973, 10), 1712 => to_unsigned(1014, 10), 1713 => to_unsigned(192, 10), 1714 => to_unsigned(750, 10), 1715 => to_unsigned(60, 10), 1716 => to_unsigned(840, 10), 1717 => to_unsigned(718, 10), 1718 => to_unsigned(776, 10), 1719 => to_unsigned(753, 10), 1720 => to_unsigned(873, 10), 1721 => to_unsigned(1017, 10), 1722 => to_unsigned(897, 10), 1723 => to_unsigned(449, 10), 1724 => to_unsigned(386, 10), 1725 => to_unsigned(271, 10), 1726 => to_unsigned(149, 10), 1727 => to_unsigned(942, 10), 1728 => to_unsigned(258, 10), 1729 => to_unsigned(848, 10), 1730 => to_unsigned(993, 10), 1731 => to_unsigned(720, 10), 1732 => to_unsigned(154, 10), 1733 => to_unsigned(71, 10), 1734 => to_unsigned(752, 10), 1735 => to_unsigned(909, 10), 1736 => to_unsigned(739, 10), 1737 => to_unsigned(132, 10), 1738 => to_unsigned(426, 10), 1739 => to_unsigned(710, 10), 1740 => to_unsigned(682, 10), 1741 => to_unsigned(763, 10), 1742 => to_unsigned(716, 10), 1743 => to_unsigned(353, 10), 1744 => to_unsigned(204, 10), 1745 => to_unsigned(62, 10), 1746 => to_unsigned(371, 10), 1747 => to_unsigned(684, 10), 1748 => to_unsigned(227, 10), 1749 => to_unsigned(461, 10), 1750 => to_unsigned(726, 10), 1751 => to_unsigned(55, 10), 1752 => to_unsigned(535, 10), 1753 => to_unsigned(587, 10), 1754 => to_unsigned(609, 10), 1755 => to_unsigned(937, 10), 1756 => to_unsigned(764, 10), 1757 => to_unsigned(782, 10), 1758 => to_unsigned(281, 10), 1759 => to_unsigned(746, 10), 1760 => to_unsigned(14, 10), 1761 => to_unsigned(108, 10), 1762 => to_unsigned(632, 10), 1763 => to_unsigned(671, 10), 1764 => to_unsigned(604, 10), 1765 => to_unsigned(750, 10), 1766 => to_unsigned(462, 10), 1767 => to_unsigned(114, 10), 1768 => to_unsigned(136, 10), 1769 => to_unsigned(790, 10), 1770 => to_unsigned(124, 10), 1771 => to_unsigned(110, 10), 1772 => to_unsigned(899, 10), 1773 => to_unsigned(515, 10), 1774 => to_unsigned(45, 10), 1775 => to_unsigned(120, 10), 1776 => to_unsigned(213, 10), 1777 => to_unsigned(767, 10), 1778 => to_unsigned(471, 10), 1779 => to_unsigned(679, 10), 1780 => to_unsigned(360, 10), 1781 => to_unsigned(129, 10), 1782 => to_unsigned(964, 10), 1783 => to_unsigned(298, 10), 1784 => to_unsigned(400, 10), 1785 => to_unsigned(784, 10), 1786 => to_unsigned(238, 10), 1787 => to_unsigned(929, 10), 1788 => to_unsigned(212, 10), 1789 => to_unsigned(601, 10), 1790 => to_unsigned(384, 10), 1791 => to_unsigned(451, 10), 1792 => to_unsigned(256, 10), 1793 => to_unsigned(773, 10), 1794 => to_unsigned(713, 10), 1795 => to_unsigned(445, 10), 1796 => to_unsigned(117, 10), 1797 => to_unsigned(962, 10), 1798 => to_unsigned(84, 10), 1799 => to_unsigned(87, 10), 1800 => to_unsigned(749, 10), 1801 => to_unsigned(561, 10), 1802 => to_unsigned(138, 10), 1803 => to_unsigned(155, 10), 1804 => to_unsigned(826, 10), 1805 => to_unsigned(42, 10), 1806 => to_unsigned(556, 10), 1807 => to_unsigned(253, 10), 1808 => to_unsigned(253, 10), 1809 => to_unsigned(550, 10), 1810 => to_unsigned(652, 10), 1811 => to_unsigned(138, 10), 1812 => to_unsigned(97, 10), 1813 => to_unsigned(288, 10), 1814 => to_unsigned(399, 10), 1815 => to_unsigned(304, 10), 1816 => to_unsigned(47, 10), 1817 => to_unsigned(985, 10), 1818 => to_unsigned(158, 10), 1819 => to_unsigned(534, 10), 1820 => to_unsigned(691, 10), 1821 => to_unsigned(305, 10), 1822 => to_unsigned(936, 10), 1823 => to_unsigned(908, 10), 1824 => to_unsigned(460, 10), 1825 => to_unsigned(180, 10), 1826 => to_unsigned(119, 10), 1827 => to_unsigned(524, 10), 1828 => to_unsigned(540, 10), 1829 => to_unsigned(749, 10), 1830 => to_unsigned(82, 10), 1831 => to_unsigned(691, 10), 1832 => to_unsigned(220, 10), 1833 => to_unsigned(171, 10), 1834 => to_unsigned(811, 10), 1835 => to_unsigned(42, 10), 1836 => to_unsigned(123, 10), 1837 => to_unsigned(454, 10), 1838 => to_unsigned(822, 10), 1839 => to_unsigned(985, 10), 1840 => to_unsigned(536, 10), 1841 => to_unsigned(772, 10), 1842 => to_unsigned(862, 10), 1843 => to_unsigned(572, 10), 1844 => to_unsigned(972, 10), 1845 => to_unsigned(782, 10), 1846 => to_unsigned(182, 10), 1847 => to_unsigned(562, 10), 1848 => to_unsigned(655, 10), 1849 => to_unsigned(103, 10), 1850 => to_unsigned(688, 10), 1851 => to_unsigned(140, 10), 1852 => to_unsigned(920, 10), 1853 => to_unsigned(479, 10), 1854 => to_unsigned(465, 10), 1855 => to_unsigned(582, 10), 1856 => to_unsigned(391, 10), 1857 => to_unsigned(905, 10), 1858 => to_unsigned(332, 10), 1859 => to_unsigned(564, 10), 1860 => to_unsigned(785, 10), 1861 => to_unsigned(421, 10), 1862 => to_unsigned(951, 10), 1863 => to_unsigned(729, 10), 1864 => to_unsigned(72, 10), 1865 => to_unsigned(894, 10), 1866 => to_unsigned(533, 10), 1867 => to_unsigned(273, 10), 1868 => to_unsigned(68, 10), 1869 => to_unsigned(925, 10), 1870 => to_unsigned(421, 10), 1871 => to_unsigned(153, 10), 1872 => to_unsigned(200, 10), 1873 => to_unsigned(999, 10), 1874 => to_unsigned(11, 10), 1875 => to_unsigned(599, 10), 1876 => to_unsigned(91, 10), 1877 => to_unsigned(912, 10), 1878 => to_unsigned(968, 10), 1879 => to_unsigned(20, 10), 1880 => to_unsigned(289, 10), 1881 => to_unsigned(537, 10), 1882 => to_unsigned(334, 10), 1883 => to_unsigned(137, 10), 1884 => to_unsigned(921, 10), 1885 => to_unsigned(708, 10), 1886 => to_unsigned(358, 10), 1887 => to_unsigned(97, 10), 1888 => to_unsigned(244, 10), 1889 => to_unsigned(256, 10), 1890 => to_unsigned(296, 10), 1891 => to_unsigned(717, 10), 1892 => to_unsigned(718, 10), 1893 => to_unsigned(715, 10), 1894 => to_unsigned(5, 10), 1895 => to_unsigned(24, 10), 1896 => to_unsigned(251, 10), 1897 => to_unsigned(781, 10), 1898 => to_unsigned(378, 10), 1899 => to_unsigned(746, 10), 1900 => to_unsigned(706, 10), 1901 => to_unsigned(898, 10), 1902 => to_unsigned(905, 10), 1903 => to_unsigned(992, 10), 1904 => to_unsigned(705, 10), 1905 => to_unsigned(237, 10), 1906 => to_unsigned(750, 10), 1907 => to_unsigned(1020, 10), 1908 => to_unsigned(39, 10), 1909 => to_unsigned(65, 10), 1910 => to_unsigned(850, 10), 1911 => to_unsigned(1015, 10), 1912 => to_unsigned(922, 10), 1913 => to_unsigned(681, 10), 1914 => to_unsigned(79, 10), 1915 => to_unsigned(647, 10), 1916 => to_unsigned(771, 10), 1917 => to_unsigned(879, 10), 1918 => to_unsigned(121, 10), 1919 => to_unsigned(936, 10), 1920 => to_unsigned(164, 10), 1921 => to_unsigned(813, 10), 1922 => to_unsigned(32, 10), 1923 => to_unsigned(590, 10), 1924 => to_unsigned(813, 10), 1925 => to_unsigned(302, 10), 1926 => to_unsigned(165, 10), 1927 => to_unsigned(1012, 10), 1928 => to_unsigned(996, 10), 1929 => to_unsigned(414, 10), 1930 => to_unsigned(651, 10), 1931 => to_unsigned(340, 10), 1932 => to_unsigned(374, 10), 1933 => to_unsigned(937, 10), 1934 => to_unsigned(740, 10), 1935 => to_unsigned(759, 10), 1936 => to_unsigned(920, 10), 1937 => to_unsigned(1008, 10), 1938 => to_unsigned(298, 10), 1939 => to_unsigned(808, 10), 1940 => to_unsigned(11, 10), 1941 => to_unsigned(545, 10), 1942 => to_unsigned(808, 10), 1943 => to_unsigned(685, 10), 1944 => to_unsigned(819, 10), 1945 => to_unsigned(502, 10), 1946 => to_unsigned(20, 10), 1947 => to_unsigned(916, 10), 1948 => to_unsigned(994, 10), 1949 => to_unsigned(332, 10), 1950 => to_unsigned(657, 10), 1951 => to_unsigned(7, 10), 1952 => to_unsigned(69, 10), 1953 => to_unsigned(840, 10), 1954 => to_unsigned(687, 10), 1955 => to_unsigned(803, 10), 1956 => to_unsigned(434, 10), 1957 => to_unsigned(887, 10), 1958 => to_unsigned(892, 10), 1959 => to_unsigned(957, 10), 1960 => to_unsigned(622, 10), 1961 => to_unsigned(683, 10), 1962 => to_unsigned(548, 10), 1963 => to_unsigned(926, 10), 1964 => to_unsigned(384, 10), 1965 => to_unsigned(154, 10), 1966 => to_unsigned(370, 10), 1967 => to_unsigned(863, 10), 1968 => to_unsigned(5, 10), 1969 => to_unsigned(940, 10), 1970 => to_unsigned(675, 10), 1971 => to_unsigned(117, 10), 1972 => to_unsigned(838, 10), 1973 => to_unsigned(722, 10), 1974 => to_unsigned(664, 10), 1975 => to_unsigned(532, 10), 1976 => to_unsigned(459, 10), 1977 => to_unsigned(490, 10), 1978 => to_unsigned(1003, 10), 1979 => to_unsigned(788, 10), 1980 => to_unsigned(812, 10), 1981 => to_unsigned(276, 10), 1982 => to_unsigned(605, 10), 1983 => to_unsigned(117, 10), 1984 => to_unsigned(696, 10), 1985 => to_unsigned(974, 10), 1986 => to_unsigned(64, 10), 1987 => to_unsigned(687, 10), 1988 => to_unsigned(586, 10), 1989 => to_unsigned(382, 10), 1990 => to_unsigned(629, 10), 1991 => to_unsigned(246, 10), 1992 => to_unsigned(434, 10), 1993 => to_unsigned(283, 10), 1994 => to_unsigned(726, 10), 1995 => to_unsigned(297, 10), 1996 => to_unsigned(178, 10), 1997 => to_unsigned(775, 10), 1998 => to_unsigned(200, 10), 1999 => to_unsigned(749, 10), 2000 => to_unsigned(32, 10), 2001 => to_unsigned(545, 10), 2002 => to_unsigned(825, 10), 2003 => to_unsigned(214, 10), 2004 => to_unsigned(25, 10), 2005 => to_unsigned(600, 10), 2006 => to_unsigned(126, 10), 2007 => to_unsigned(595, 10), 2008 => to_unsigned(536, 10), 2009 => to_unsigned(127, 10), 2010 => to_unsigned(363, 10), 2011 => to_unsigned(954, 10), 2012 => to_unsigned(31, 10), 2013 => to_unsigned(832, 10), 2014 => to_unsigned(190, 10), 2015 => to_unsigned(617, 10), 2016 => to_unsigned(323, 10), 2017 => to_unsigned(881, 10), 2018 => to_unsigned(421, 10), 2019 => to_unsigned(509, 10), 2020 => to_unsigned(425, 10), 2021 => to_unsigned(630, 10), 2022 => to_unsigned(688, 10), 2023 => to_unsigned(108, 10), 2024 => to_unsigned(265, 10), 2025 => to_unsigned(957, 10), 2026 => to_unsigned(639, 10), 2027 => to_unsigned(53, 10), 2028 => to_unsigned(852, 10), 2029 => to_unsigned(685, 10), 2030 => to_unsigned(792, 10), 2031 => to_unsigned(294, 10), 2032 => to_unsigned(247, 10), 2033 => to_unsigned(547, 10), 2034 => to_unsigned(380, 10), 2035 => to_unsigned(581, 10), 2036 => to_unsigned(934, 10), 2037 => to_unsigned(227, 10), 2038 => to_unsigned(868, 10), 2039 => to_unsigned(581, 10), 2040 => to_unsigned(281, 10), 2041 => to_unsigned(356, 10), 2042 => to_unsigned(376, 10), 2043 => to_unsigned(15, 10), 2044 => to_unsigned(257, 10), 2045 => to_unsigned(254, 10), 2046 => to_unsigned(182, 10), 2047 => to_unsigned(801, 10)),
            9 => (0 => to_unsigned(711, 10), 1 => to_unsigned(558, 10), 2 => to_unsigned(477, 10), 3 => to_unsigned(90, 10), 4 => to_unsigned(184, 10), 5 => to_unsigned(90, 10), 6 => to_unsigned(395, 10), 7 => to_unsigned(677, 10), 8 => to_unsigned(451, 10), 9 => to_unsigned(153, 10), 10 => to_unsigned(224, 10), 11 => to_unsigned(644, 10), 12 => to_unsigned(64, 10), 13 => to_unsigned(536, 10), 14 => to_unsigned(518, 10), 15 => to_unsigned(132, 10), 16 => to_unsigned(416, 10), 17 => to_unsigned(619, 10), 18 => to_unsigned(344, 10), 19 => to_unsigned(507, 10), 20 => to_unsigned(627, 10), 21 => to_unsigned(852, 10), 22 => to_unsigned(689, 10), 23 => to_unsigned(827, 10), 24 => to_unsigned(906, 10), 25 => to_unsigned(340, 10), 26 => to_unsigned(609, 10), 27 => to_unsigned(579, 10), 28 => to_unsigned(654, 10), 29 => to_unsigned(106, 10), 30 => to_unsigned(964, 10), 31 => to_unsigned(592, 10), 32 => to_unsigned(3, 10), 33 => to_unsigned(758, 10), 34 => to_unsigned(581, 10), 35 => to_unsigned(440, 10), 36 => to_unsigned(4, 10), 37 => to_unsigned(627, 10), 38 => to_unsigned(470, 10), 39 => to_unsigned(540, 10), 40 => to_unsigned(1, 10), 41 => to_unsigned(904, 10), 42 => to_unsigned(230, 10), 43 => to_unsigned(616, 10), 44 => to_unsigned(458, 10), 45 => to_unsigned(228, 10), 46 => to_unsigned(847, 10), 47 => to_unsigned(831, 10), 48 => to_unsigned(188, 10), 49 => to_unsigned(905, 10), 50 => to_unsigned(582, 10), 51 => to_unsigned(599, 10), 52 => to_unsigned(890, 10), 53 => to_unsigned(756, 10), 54 => to_unsigned(92, 10), 55 => to_unsigned(107, 10), 56 => to_unsigned(19, 10), 57 => to_unsigned(404, 10), 58 => to_unsigned(343, 10), 59 => to_unsigned(1002, 10), 60 => to_unsigned(1000, 10), 61 => to_unsigned(296, 10), 62 => to_unsigned(461, 10), 63 => to_unsigned(947, 10), 64 => to_unsigned(378, 10), 65 => to_unsigned(947, 10), 66 => to_unsigned(996, 10), 67 => to_unsigned(987, 10), 68 => to_unsigned(103, 10), 69 => to_unsigned(358, 10), 70 => to_unsigned(984, 10), 71 => to_unsigned(498, 10), 72 => to_unsigned(246, 10), 73 => to_unsigned(1008, 10), 74 => to_unsigned(363, 10), 75 => to_unsigned(602, 10), 76 => to_unsigned(238, 10), 77 => to_unsigned(789, 10), 78 => to_unsigned(78, 10), 79 => to_unsigned(755, 10), 80 => to_unsigned(119, 10), 81 => to_unsigned(505, 10), 82 => to_unsigned(652, 10), 83 => to_unsigned(204, 10), 84 => to_unsigned(156, 10), 85 => to_unsigned(46, 10), 86 => to_unsigned(674, 10), 87 => to_unsigned(715, 10), 88 => to_unsigned(362, 10), 89 => to_unsigned(784, 10), 90 => to_unsigned(297, 10), 91 => to_unsigned(973, 10), 92 => to_unsigned(551, 10), 93 => to_unsigned(85, 10), 94 => to_unsigned(239, 10), 95 => to_unsigned(904, 10), 96 => to_unsigned(569, 10), 97 => to_unsigned(141, 10), 98 => to_unsigned(285, 10), 99 => to_unsigned(676, 10), 100 => to_unsigned(478, 10), 101 => to_unsigned(1015, 10), 102 => to_unsigned(429, 10), 103 => to_unsigned(25, 10), 104 => to_unsigned(782, 10), 105 => to_unsigned(359, 10), 106 => to_unsigned(6, 10), 107 => to_unsigned(484, 10), 108 => to_unsigned(607, 10), 109 => to_unsigned(894, 10), 110 => to_unsigned(296, 10), 111 => to_unsigned(729, 10), 112 => to_unsigned(877, 10), 113 => to_unsigned(111, 10), 114 => to_unsigned(544, 10), 115 => to_unsigned(984, 10), 116 => to_unsigned(161, 10), 117 => to_unsigned(495, 10), 118 => to_unsigned(426, 10), 119 => to_unsigned(281, 10), 120 => to_unsigned(412, 10), 121 => to_unsigned(589, 10), 122 => to_unsigned(931, 10), 123 => to_unsigned(419, 10), 124 => to_unsigned(202, 10), 125 => to_unsigned(1010, 10), 126 => to_unsigned(24, 10), 127 => to_unsigned(162, 10), 128 => to_unsigned(743, 10), 129 => to_unsigned(695, 10), 130 => to_unsigned(849, 10), 131 => to_unsigned(764, 10), 132 => to_unsigned(286, 10), 133 => to_unsigned(756, 10), 134 => to_unsigned(750, 10), 135 => to_unsigned(740, 10), 136 => to_unsigned(187, 10), 137 => to_unsigned(350, 10), 138 => to_unsigned(128, 10), 139 => to_unsigned(656, 10), 140 => to_unsigned(582, 10), 141 => to_unsigned(536, 10), 142 => to_unsigned(350, 10), 143 => to_unsigned(440, 10), 144 => to_unsigned(347, 10), 145 => to_unsigned(611, 10), 146 => to_unsigned(287, 10), 147 => to_unsigned(211, 10), 148 => to_unsigned(610, 10), 149 => to_unsigned(583, 10), 150 => to_unsigned(408, 10), 151 => to_unsigned(855, 10), 152 => to_unsigned(130, 10), 153 => to_unsigned(946, 10), 154 => to_unsigned(925, 10), 155 => to_unsigned(805, 10), 156 => to_unsigned(100, 10), 157 => to_unsigned(832, 10), 158 => to_unsigned(337, 10), 159 => to_unsigned(402, 10), 160 => to_unsigned(584, 10), 161 => to_unsigned(902, 10), 162 => to_unsigned(630, 10), 163 => to_unsigned(720, 10), 164 => to_unsigned(416, 10), 165 => to_unsigned(162, 10), 166 => to_unsigned(778, 10), 167 => to_unsigned(832, 10), 168 => to_unsigned(595, 10), 169 => to_unsigned(300, 10), 170 => to_unsigned(442, 10), 171 => to_unsigned(158, 10), 172 => to_unsigned(482, 10), 173 => to_unsigned(71, 10), 174 => to_unsigned(515, 10), 175 => to_unsigned(712, 10), 176 => to_unsigned(907, 10), 177 => to_unsigned(3, 10), 178 => to_unsigned(886, 10), 179 => to_unsigned(976, 10), 180 => to_unsigned(341, 10), 181 => to_unsigned(634, 10), 182 => to_unsigned(991, 10), 183 => to_unsigned(994, 10), 184 => to_unsigned(24, 10), 185 => to_unsigned(356, 10), 186 => to_unsigned(191, 10), 187 => to_unsigned(799, 10), 188 => to_unsigned(505, 10), 189 => to_unsigned(635, 10), 190 => to_unsigned(392, 10), 191 => to_unsigned(849, 10), 192 => to_unsigned(542, 10), 193 => to_unsigned(38, 10), 194 => to_unsigned(764, 10), 195 => to_unsigned(675, 10), 196 => to_unsigned(568, 10), 197 => to_unsigned(669, 10), 198 => to_unsigned(656, 10), 199 => to_unsigned(755, 10), 200 => to_unsigned(435, 10), 201 => to_unsigned(554, 10), 202 => to_unsigned(486, 10), 203 => to_unsigned(671, 10), 204 => to_unsigned(419, 10), 205 => to_unsigned(508, 10), 206 => to_unsigned(462, 10), 207 => to_unsigned(578, 10), 208 => to_unsigned(706, 10), 209 => to_unsigned(322, 10), 210 => to_unsigned(372, 10), 211 => to_unsigned(443, 10), 212 => to_unsigned(104, 10), 213 => to_unsigned(688, 10), 214 => to_unsigned(341, 10), 215 => to_unsigned(418, 10), 216 => to_unsigned(360, 10), 217 => to_unsigned(858, 10), 218 => to_unsigned(859, 10), 219 => to_unsigned(395, 10), 220 => to_unsigned(659, 10), 221 => to_unsigned(946, 10), 222 => to_unsigned(804, 10), 223 => to_unsigned(875, 10), 224 => to_unsigned(367, 10), 225 => to_unsigned(212, 10), 226 => to_unsigned(372, 10), 227 => to_unsigned(800, 10), 228 => to_unsigned(291, 10), 229 => to_unsigned(747, 10), 230 => to_unsigned(885, 10), 231 => to_unsigned(28, 10), 232 => to_unsigned(441, 10), 233 => to_unsigned(433, 10), 234 => to_unsigned(378, 10), 235 => to_unsigned(177, 10), 236 => to_unsigned(810, 10), 237 => to_unsigned(981, 10), 238 => to_unsigned(935, 10), 239 => to_unsigned(692, 10), 240 => to_unsigned(591, 10), 241 => to_unsigned(539, 10), 242 => to_unsigned(802, 10), 243 => to_unsigned(959, 10), 244 => to_unsigned(74, 10), 245 => to_unsigned(591, 10), 246 => to_unsigned(272, 10), 247 => to_unsigned(867, 10), 248 => to_unsigned(543, 10), 249 => to_unsigned(814, 10), 250 => to_unsigned(171, 10), 251 => to_unsigned(69, 10), 252 => to_unsigned(322, 10), 253 => to_unsigned(258, 10), 254 => to_unsigned(915, 10), 255 => to_unsigned(414, 10), 256 => to_unsigned(633, 10), 257 => to_unsigned(805, 10), 258 => to_unsigned(936, 10), 259 => to_unsigned(257, 10), 260 => to_unsigned(103, 10), 261 => to_unsigned(437, 10), 262 => to_unsigned(772, 10), 263 => to_unsigned(546, 10), 264 => to_unsigned(277, 10), 265 => to_unsigned(490, 10), 266 => to_unsigned(179, 10), 267 => to_unsigned(716, 10), 268 => to_unsigned(737, 10), 269 => to_unsigned(1014, 10), 270 => to_unsigned(948, 10), 271 => to_unsigned(777, 10), 272 => to_unsigned(229, 10), 273 => to_unsigned(787, 10), 274 => to_unsigned(625, 10), 275 => to_unsigned(95, 10), 276 => to_unsigned(1005, 10), 277 => to_unsigned(68, 10), 278 => to_unsigned(5, 10), 279 => to_unsigned(91, 10), 280 => to_unsigned(102, 10), 281 => to_unsigned(437, 10), 282 => to_unsigned(977, 10), 283 => to_unsigned(846, 10), 284 => to_unsigned(361, 10), 285 => to_unsigned(840, 10), 286 => to_unsigned(209, 10), 287 => to_unsigned(208, 10), 288 => to_unsigned(964, 10), 289 => to_unsigned(237, 10), 290 => to_unsigned(41, 10), 291 => to_unsigned(413, 10), 292 => to_unsigned(176, 10), 293 => to_unsigned(667, 10), 294 => to_unsigned(578, 10), 295 => to_unsigned(356, 10), 296 => to_unsigned(603, 10), 297 => to_unsigned(949, 10), 298 => to_unsigned(687, 10), 299 => to_unsigned(123, 10), 300 => to_unsigned(581, 10), 301 => to_unsigned(750, 10), 302 => to_unsigned(764, 10), 303 => to_unsigned(475, 10), 304 => to_unsigned(501, 10), 305 => to_unsigned(123, 10), 306 => to_unsigned(912, 10), 307 => to_unsigned(178, 10), 308 => to_unsigned(739, 10), 309 => to_unsigned(682, 10), 310 => to_unsigned(640, 10), 311 => to_unsigned(332, 10), 312 => to_unsigned(263, 10), 313 => to_unsigned(602, 10), 314 => to_unsigned(656, 10), 315 => to_unsigned(696, 10), 316 => to_unsigned(96, 10), 317 => to_unsigned(983, 10), 318 => to_unsigned(826, 10), 319 => to_unsigned(15, 10), 320 => to_unsigned(185, 10), 321 => to_unsigned(427, 10), 322 => to_unsigned(381, 10), 323 => to_unsigned(344, 10), 324 => to_unsigned(486, 10), 325 => to_unsigned(268, 10), 326 => to_unsigned(361, 10), 327 => to_unsigned(225, 10), 328 => to_unsigned(648, 10), 329 => to_unsigned(668, 10), 330 => to_unsigned(139, 10), 331 => to_unsigned(672, 10), 332 => to_unsigned(589, 10), 333 => to_unsigned(338, 10), 334 => to_unsigned(589, 10), 335 => to_unsigned(518, 10), 336 => to_unsigned(722, 10), 337 => to_unsigned(1003, 10), 338 => to_unsigned(716, 10), 339 => to_unsigned(847, 10), 340 => to_unsigned(890, 10), 341 => to_unsigned(661, 10), 342 => to_unsigned(937, 10), 343 => to_unsigned(532, 10), 344 => to_unsigned(730, 10), 345 => to_unsigned(145, 10), 346 => to_unsigned(69, 10), 347 => to_unsigned(988, 10), 348 => to_unsigned(32, 10), 349 => to_unsigned(407, 10), 350 => to_unsigned(46, 10), 351 => to_unsigned(26, 10), 352 => to_unsigned(140, 10), 353 => to_unsigned(396, 10), 354 => to_unsigned(771, 10), 355 => to_unsigned(206, 10), 356 => to_unsigned(462, 10), 357 => to_unsigned(32, 10), 358 => to_unsigned(524, 10), 359 => to_unsigned(545, 10), 360 => to_unsigned(284, 10), 361 => to_unsigned(653, 10), 362 => to_unsigned(636, 10), 363 => to_unsigned(588, 10), 364 => to_unsigned(287, 10), 365 => to_unsigned(975, 10), 366 => to_unsigned(108, 10), 367 => to_unsigned(703, 10), 368 => to_unsigned(599, 10), 369 => to_unsigned(92, 10), 370 => to_unsigned(729, 10), 371 => to_unsigned(298, 10), 372 => to_unsigned(2, 10), 373 => to_unsigned(218, 10), 374 => to_unsigned(473, 10), 375 => to_unsigned(871, 10), 376 => to_unsigned(760, 10), 377 => to_unsigned(878, 10), 378 => to_unsigned(680, 10), 379 => to_unsigned(1004, 10), 380 => to_unsigned(705, 10), 381 => to_unsigned(947, 10), 382 => to_unsigned(829, 10), 383 => to_unsigned(613, 10), 384 => to_unsigned(695, 10), 385 => to_unsigned(598, 10), 386 => to_unsigned(719, 10), 387 => to_unsigned(199, 10), 388 => to_unsigned(892, 10), 389 => to_unsigned(742, 10), 390 => to_unsigned(699, 10), 391 => to_unsigned(676, 10), 392 => to_unsigned(822, 10), 393 => to_unsigned(599, 10), 394 => to_unsigned(384, 10), 395 => to_unsigned(535, 10), 396 => to_unsigned(707, 10), 397 => to_unsigned(391, 10), 398 => to_unsigned(660, 10), 399 => to_unsigned(760, 10), 400 => to_unsigned(626, 10), 401 => to_unsigned(918, 10), 402 => to_unsigned(114, 10), 403 => to_unsigned(358, 10), 404 => to_unsigned(862, 10), 405 => to_unsigned(539, 10), 406 => to_unsigned(427, 10), 407 => to_unsigned(123, 10), 408 => to_unsigned(65, 10), 409 => to_unsigned(27, 10), 410 => to_unsigned(223, 10), 411 => to_unsigned(838, 10), 412 => to_unsigned(935, 10), 413 => to_unsigned(501, 10), 414 => to_unsigned(52, 10), 415 => to_unsigned(389, 10), 416 => to_unsigned(82, 10), 417 => to_unsigned(584, 10), 418 => to_unsigned(870, 10), 419 => to_unsigned(404, 10), 420 => to_unsigned(89, 10), 421 => to_unsigned(98, 10), 422 => to_unsigned(399, 10), 423 => to_unsigned(512, 10), 424 => to_unsigned(466, 10), 425 => to_unsigned(32, 10), 426 => to_unsigned(180, 10), 427 => to_unsigned(707, 10), 428 => to_unsigned(765, 10), 429 => to_unsigned(211, 10), 430 => to_unsigned(118, 10), 431 => to_unsigned(303, 10), 432 => to_unsigned(637, 10), 433 => to_unsigned(788, 10), 434 => to_unsigned(987, 10), 435 => to_unsigned(684, 10), 436 => to_unsigned(240, 10), 437 => to_unsigned(743, 10), 438 => to_unsigned(526, 10), 439 => to_unsigned(612, 10), 440 => to_unsigned(421, 10), 441 => to_unsigned(927, 10), 442 => to_unsigned(647, 10), 443 => to_unsigned(601, 10), 444 => to_unsigned(706, 10), 445 => to_unsigned(248, 10), 446 => to_unsigned(411, 10), 447 => to_unsigned(244, 10), 448 => to_unsigned(840, 10), 449 => to_unsigned(285, 10), 450 => to_unsigned(906, 10), 451 => to_unsigned(897, 10), 452 => to_unsigned(843, 10), 453 => to_unsigned(576, 10), 454 => to_unsigned(295, 10), 455 => to_unsigned(475, 10), 456 => to_unsigned(847, 10), 457 => to_unsigned(526, 10), 458 => to_unsigned(245, 10), 459 => to_unsigned(1000, 10), 460 => to_unsigned(350, 10), 461 => to_unsigned(9, 10), 462 => to_unsigned(256, 10), 463 => to_unsigned(170, 10), 464 => to_unsigned(119, 10), 465 => to_unsigned(189, 10), 466 => to_unsigned(907, 10), 467 => to_unsigned(916, 10), 468 => to_unsigned(934, 10), 469 => to_unsigned(543, 10), 470 => to_unsigned(399, 10), 471 => to_unsigned(0, 10), 472 => to_unsigned(232, 10), 473 => to_unsigned(930, 10), 474 => to_unsigned(816, 10), 475 => to_unsigned(151, 10), 476 => to_unsigned(967, 10), 477 => to_unsigned(446, 10), 478 => to_unsigned(446, 10), 479 => to_unsigned(746, 10), 480 => to_unsigned(37, 10), 481 => to_unsigned(856, 10), 482 => to_unsigned(156, 10), 483 => to_unsigned(208, 10), 484 => to_unsigned(690, 10), 485 => to_unsigned(1023, 10), 486 => to_unsigned(842, 10), 487 => to_unsigned(366, 10), 488 => to_unsigned(981, 10), 489 => to_unsigned(333, 10), 490 => to_unsigned(92, 10), 491 => to_unsigned(1012, 10), 492 => to_unsigned(294, 10), 493 => to_unsigned(484, 10), 494 => to_unsigned(262, 10), 495 => to_unsigned(200, 10), 496 => to_unsigned(934, 10), 497 => to_unsigned(379, 10), 498 => to_unsigned(231, 10), 499 => to_unsigned(36, 10), 500 => to_unsigned(797, 10), 501 => to_unsigned(699, 10), 502 => to_unsigned(380, 10), 503 => to_unsigned(652, 10), 504 => to_unsigned(591, 10), 505 => to_unsigned(905, 10), 506 => to_unsigned(1009, 10), 507 => to_unsigned(932, 10), 508 => to_unsigned(153, 10), 509 => to_unsigned(781, 10), 510 => to_unsigned(689, 10), 511 => to_unsigned(582, 10), 512 => to_unsigned(370, 10), 513 => to_unsigned(613, 10), 514 => to_unsigned(926, 10), 515 => to_unsigned(433, 10), 516 => to_unsigned(19, 10), 517 => to_unsigned(540, 10), 518 => to_unsigned(972, 10), 519 => to_unsigned(635, 10), 520 => to_unsigned(40, 10), 521 => to_unsigned(1012, 10), 522 => to_unsigned(608, 10), 523 => to_unsigned(249, 10), 524 => to_unsigned(865, 10), 525 => to_unsigned(460, 10), 526 => to_unsigned(823, 10), 527 => to_unsigned(805, 10), 528 => to_unsigned(16, 10), 529 => to_unsigned(722, 10), 530 => to_unsigned(797, 10), 531 => to_unsigned(151, 10), 532 => to_unsigned(948, 10), 533 => to_unsigned(660, 10), 534 => to_unsigned(255, 10), 535 => to_unsigned(855, 10), 536 => to_unsigned(257, 10), 537 => to_unsigned(755, 10), 538 => to_unsigned(683, 10), 539 => to_unsigned(280, 10), 540 => to_unsigned(503, 10), 541 => to_unsigned(157, 10), 542 => to_unsigned(930, 10), 543 => to_unsigned(109, 10), 544 => to_unsigned(1001, 10), 545 => to_unsigned(882, 10), 546 => to_unsigned(454, 10), 547 => to_unsigned(98, 10), 548 => to_unsigned(203, 10), 549 => to_unsigned(608, 10), 550 => to_unsigned(387, 10), 551 => to_unsigned(626, 10), 552 => to_unsigned(81, 10), 553 => to_unsigned(712, 10), 554 => to_unsigned(812, 10), 555 => to_unsigned(218, 10), 556 => to_unsigned(58, 10), 557 => to_unsigned(202, 10), 558 => to_unsigned(848, 10), 559 => to_unsigned(602, 10), 560 => to_unsigned(815, 10), 561 => to_unsigned(15, 10), 562 => to_unsigned(642, 10), 563 => to_unsigned(666, 10), 564 => to_unsigned(954, 10), 565 => to_unsigned(278, 10), 566 => to_unsigned(332, 10), 567 => to_unsigned(144, 10), 568 => to_unsigned(405, 10), 569 => to_unsigned(403, 10), 570 => to_unsigned(133, 10), 571 => to_unsigned(689, 10), 572 => to_unsigned(504, 10), 573 => to_unsigned(275, 10), 574 => to_unsigned(35, 10), 575 => to_unsigned(183, 10), 576 => to_unsigned(531, 10), 577 => to_unsigned(518, 10), 578 => to_unsigned(502, 10), 579 => to_unsigned(339, 10), 580 => to_unsigned(798, 10), 581 => to_unsigned(625, 10), 582 => to_unsigned(491, 10), 583 => to_unsigned(92, 10), 584 => to_unsigned(383, 10), 585 => to_unsigned(903, 10), 586 => to_unsigned(265, 10), 587 => to_unsigned(733, 10), 588 => to_unsigned(829, 10), 589 => to_unsigned(606, 10), 590 => to_unsigned(890, 10), 591 => to_unsigned(634, 10), 592 => to_unsigned(913, 10), 593 => to_unsigned(903, 10), 594 => to_unsigned(307, 10), 595 => to_unsigned(689, 10), 596 => to_unsigned(64, 10), 597 => to_unsigned(854, 10), 598 => to_unsigned(797, 10), 599 => to_unsigned(823, 10), 600 => to_unsigned(483, 10), 601 => to_unsigned(884, 10), 602 => to_unsigned(945, 10), 603 => to_unsigned(693, 10), 604 => to_unsigned(669, 10), 605 => to_unsigned(268, 10), 606 => to_unsigned(600, 10), 607 => to_unsigned(228, 10), 608 => to_unsigned(686, 10), 609 => to_unsigned(304, 10), 610 => to_unsigned(942, 10), 611 => to_unsigned(457, 10), 612 => to_unsigned(222, 10), 613 => to_unsigned(144, 10), 614 => to_unsigned(122, 10), 615 => to_unsigned(632, 10), 616 => to_unsigned(905, 10), 617 => to_unsigned(1016, 10), 618 => to_unsigned(348, 10), 619 => to_unsigned(478, 10), 620 => to_unsigned(532, 10), 621 => to_unsigned(96, 10), 622 => to_unsigned(527, 10), 623 => to_unsigned(1010, 10), 624 => to_unsigned(934, 10), 625 => to_unsigned(620, 10), 626 => to_unsigned(780, 10), 627 => to_unsigned(114, 10), 628 => to_unsigned(591, 10), 629 => to_unsigned(651, 10), 630 => to_unsigned(843, 10), 631 => to_unsigned(157, 10), 632 => to_unsigned(659, 10), 633 => to_unsigned(103, 10), 634 => to_unsigned(346, 10), 635 => to_unsigned(10, 10), 636 => to_unsigned(572, 10), 637 => to_unsigned(1002, 10), 638 => to_unsigned(242, 10), 639 => to_unsigned(737, 10), 640 => to_unsigned(231, 10), 641 => to_unsigned(476, 10), 642 => to_unsigned(704, 10), 643 => to_unsigned(845, 10), 644 => to_unsigned(458, 10), 645 => to_unsigned(307, 10), 646 => to_unsigned(279, 10), 647 => to_unsigned(739, 10), 648 => to_unsigned(725, 10), 649 => to_unsigned(106, 10), 650 => to_unsigned(890, 10), 651 => to_unsigned(509, 10), 652 => to_unsigned(384, 10), 653 => to_unsigned(392, 10), 654 => to_unsigned(550, 10), 655 => to_unsigned(123, 10), 656 => to_unsigned(863, 10), 657 => to_unsigned(667, 10), 658 => to_unsigned(224, 10), 659 => to_unsigned(93, 10), 660 => to_unsigned(173, 10), 661 => to_unsigned(115, 10), 662 => to_unsigned(13, 10), 663 => to_unsigned(215, 10), 664 => to_unsigned(665, 10), 665 => to_unsigned(133, 10), 666 => to_unsigned(136, 10), 667 => to_unsigned(530, 10), 668 => to_unsigned(713, 10), 669 => to_unsigned(38, 10), 670 => to_unsigned(498, 10), 671 => to_unsigned(815, 10), 672 => to_unsigned(573, 10), 673 => to_unsigned(315, 10), 674 => to_unsigned(418, 10), 675 => to_unsigned(171, 10), 676 => to_unsigned(20, 10), 677 => to_unsigned(755, 10), 678 => to_unsigned(35, 10), 679 => to_unsigned(42, 10), 680 => to_unsigned(30, 10), 681 => to_unsigned(227, 10), 682 => to_unsigned(725, 10), 683 => to_unsigned(111, 10), 684 => to_unsigned(444, 10), 685 => to_unsigned(251, 10), 686 => to_unsigned(293, 10), 687 => to_unsigned(563, 10), 688 => to_unsigned(279, 10), 689 => to_unsigned(53, 10), 690 => to_unsigned(224, 10), 691 => to_unsigned(929, 10), 692 => to_unsigned(438, 10), 693 => to_unsigned(448, 10), 694 => to_unsigned(116, 10), 695 => to_unsigned(57, 10), 696 => to_unsigned(660, 10), 697 => to_unsigned(979, 10), 698 => to_unsigned(975, 10), 699 => to_unsigned(209, 10), 700 => to_unsigned(186, 10), 701 => to_unsigned(117, 10), 702 => to_unsigned(243, 10), 703 => to_unsigned(345, 10), 704 => to_unsigned(79, 10), 705 => to_unsigned(708, 10), 706 => to_unsigned(136, 10), 707 => to_unsigned(565, 10), 708 => to_unsigned(471, 10), 709 => to_unsigned(642, 10), 710 => to_unsigned(677, 10), 711 => to_unsigned(558, 10), 712 => to_unsigned(857, 10), 713 => to_unsigned(172, 10), 714 => to_unsigned(50, 10), 715 => to_unsigned(165, 10), 716 => to_unsigned(191, 10), 717 => to_unsigned(726, 10), 718 => to_unsigned(726, 10), 719 => to_unsigned(181, 10), 720 => to_unsigned(155, 10), 721 => to_unsigned(643, 10), 722 => to_unsigned(455, 10), 723 => to_unsigned(138, 10), 724 => to_unsigned(337, 10), 725 => to_unsigned(485, 10), 726 => to_unsigned(262, 10), 727 => to_unsigned(551, 10), 728 => to_unsigned(565, 10), 729 => to_unsigned(896, 10), 730 => to_unsigned(899, 10), 731 => to_unsigned(627, 10), 732 => to_unsigned(655, 10), 733 => to_unsigned(894, 10), 734 => to_unsigned(492, 10), 735 => to_unsigned(592, 10), 736 => to_unsigned(719, 10), 737 => to_unsigned(128, 10), 738 => to_unsigned(288, 10), 739 => to_unsigned(512, 10), 740 => to_unsigned(651, 10), 741 => to_unsigned(187, 10), 742 => to_unsigned(472, 10), 743 => to_unsigned(795, 10), 744 => to_unsigned(305, 10), 745 => to_unsigned(435, 10), 746 => to_unsigned(17, 10), 747 => to_unsigned(222, 10), 748 => to_unsigned(851, 10), 749 => to_unsigned(684, 10), 750 => to_unsigned(987, 10), 751 => to_unsigned(373, 10), 752 => to_unsigned(844, 10), 753 => to_unsigned(714, 10), 754 => to_unsigned(969, 10), 755 => to_unsigned(137, 10), 756 => to_unsigned(237, 10), 757 => to_unsigned(124, 10), 758 => to_unsigned(740, 10), 759 => to_unsigned(375, 10), 760 => to_unsigned(379, 10), 761 => to_unsigned(665, 10), 762 => to_unsigned(412, 10), 763 => to_unsigned(211, 10), 764 => to_unsigned(963, 10), 765 => to_unsigned(607, 10), 766 => to_unsigned(598, 10), 767 => to_unsigned(1005, 10), 768 => to_unsigned(861, 10), 769 => to_unsigned(992, 10), 770 => to_unsigned(864, 10), 771 => to_unsigned(38, 10), 772 => to_unsigned(541, 10), 773 => to_unsigned(50, 10), 774 => to_unsigned(111, 10), 775 => to_unsigned(670, 10), 776 => to_unsigned(617, 10), 777 => to_unsigned(526, 10), 778 => to_unsigned(359, 10), 779 => to_unsigned(37, 10), 780 => to_unsigned(132, 10), 781 => to_unsigned(617, 10), 782 => to_unsigned(571, 10), 783 => to_unsigned(20, 10), 784 => to_unsigned(151, 10), 785 => to_unsigned(784, 10), 786 => to_unsigned(308, 10), 787 => to_unsigned(534, 10), 788 => to_unsigned(518, 10), 789 => to_unsigned(536, 10), 790 => to_unsigned(283, 10), 791 => to_unsigned(343, 10), 792 => to_unsigned(1015, 10), 793 => to_unsigned(810, 10), 794 => to_unsigned(390, 10), 795 => to_unsigned(669, 10), 796 => to_unsigned(645, 10), 797 => to_unsigned(464, 10), 798 => to_unsigned(109, 10), 799 => to_unsigned(327, 10), 800 => to_unsigned(0, 10), 801 => to_unsigned(698, 10), 802 => to_unsigned(330, 10), 803 => to_unsigned(812, 10), 804 => to_unsigned(894, 10), 805 => to_unsigned(71, 10), 806 => to_unsigned(429, 10), 807 => to_unsigned(419, 10), 808 => to_unsigned(769, 10), 809 => to_unsigned(392, 10), 810 => to_unsigned(283, 10), 811 => to_unsigned(875, 10), 812 => to_unsigned(541, 10), 813 => to_unsigned(485, 10), 814 => to_unsigned(806, 10), 815 => to_unsigned(15, 10), 816 => to_unsigned(43, 10), 817 => to_unsigned(811, 10), 818 => to_unsigned(571, 10), 819 => to_unsigned(524, 10), 820 => to_unsigned(268, 10), 821 => to_unsigned(938, 10), 822 => to_unsigned(788, 10), 823 => to_unsigned(214, 10), 824 => to_unsigned(423, 10), 825 => to_unsigned(480, 10), 826 => to_unsigned(176, 10), 827 => to_unsigned(804, 10), 828 => to_unsigned(551, 10), 829 => to_unsigned(707, 10), 830 => to_unsigned(54, 10), 831 => to_unsigned(130, 10), 832 => to_unsigned(906, 10), 833 => to_unsigned(149, 10), 834 => to_unsigned(980, 10), 835 => to_unsigned(471, 10), 836 => to_unsigned(805, 10), 837 => to_unsigned(761, 10), 838 => to_unsigned(412, 10), 839 => to_unsigned(670, 10), 840 => to_unsigned(291, 10), 841 => to_unsigned(755, 10), 842 => to_unsigned(532, 10), 843 => to_unsigned(753, 10), 844 => to_unsigned(614, 10), 845 => to_unsigned(751, 10), 846 => to_unsigned(179, 10), 847 => to_unsigned(848, 10), 848 => to_unsigned(728, 10), 849 => to_unsigned(287, 10), 850 => to_unsigned(768, 10), 851 => to_unsigned(16, 10), 852 => to_unsigned(790, 10), 853 => to_unsigned(43, 10), 854 => to_unsigned(990, 10), 855 => to_unsigned(82, 10), 856 => to_unsigned(1019, 10), 857 => to_unsigned(370, 10), 858 => to_unsigned(894, 10), 859 => to_unsigned(798, 10), 860 => to_unsigned(633, 10), 861 => to_unsigned(833, 10), 862 => to_unsigned(38, 10), 863 => to_unsigned(806, 10), 864 => to_unsigned(83, 10), 865 => to_unsigned(362, 10), 866 => to_unsigned(309, 10), 867 => to_unsigned(667, 10), 868 => to_unsigned(443, 10), 869 => to_unsigned(270, 10), 870 => to_unsigned(210, 10), 871 => to_unsigned(749, 10), 872 => to_unsigned(302, 10), 873 => to_unsigned(756, 10), 874 => to_unsigned(369, 10), 875 => to_unsigned(565, 10), 876 => to_unsigned(125, 10), 877 => to_unsigned(689, 10), 878 => to_unsigned(465, 10), 879 => to_unsigned(17, 10), 880 => to_unsigned(917, 10), 881 => to_unsigned(709, 10), 882 => to_unsigned(17, 10), 883 => to_unsigned(899, 10), 884 => to_unsigned(803, 10), 885 => to_unsigned(951, 10), 886 => to_unsigned(910, 10), 887 => to_unsigned(371, 10), 888 => to_unsigned(556, 10), 889 => to_unsigned(804, 10), 890 => to_unsigned(4, 10), 891 => to_unsigned(834, 10), 892 => to_unsigned(120, 10), 893 => to_unsigned(107, 10), 894 => to_unsigned(555, 10), 895 => to_unsigned(509, 10), 896 => to_unsigned(70, 10), 897 => to_unsigned(546, 10), 898 => to_unsigned(477, 10), 899 => to_unsigned(543, 10), 900 => to_unsigned(322, 10), 901 => to_unsigned(725, 10), 902 => to_unsigned(361, 10), 903 => to_unsigned(1018, 10), 904 => to_unsigned(98, 10), 905 => to_unsigned(169, 10), 906 => to_unsigned(292, 10), 907 => to_unsigned(417, 10), 908 => to_unsigned(57, 10), 909 => to_unsigned(705, 10), 910 => to_unsigned(50, 10), 911 => to_unsigned(24, 10), 912 => to_unsigned(762, 10), 913 => to_unsigned(827, 10), 914 => to_unsigned(868, 10), 915 => to_unsigned(768, 10), 916 => to_unsigned(451, 10), 917 => to_unsigned(610, 10), 918 => to_unsigned(320, 10), 919 => to_unsigned(646, 10), 920 => to_unsigned(836, 10), 921 => to_unsigned(153, 10), 922 => to_unsigned(30, 10), 923 => to_unsigned(279, 10), 924 => to_unsigned(493, 10), 925 => to_unsigned(337, 10), 926 => to_unsigned(350, 10), 927 => to_unsigned(931, 10), 928 => to_unsigned(826, 10), 929 => to_unsigned(970, 10), 930 => to_unsigned(295, 10), 931 => to_unsigned(126, 10), 932 => to_unsigned(222, 10), 933 => to_unsigned(999, 10), 934 => to_unsigned(150, 10), 935 => to_unsigned(276, 10), 936 => to_unsigned(438, 10), 937 => to_unsigned(1010, 10), 938 => to_unsigned(668, 10), 939 => to_unsigned(429, 10), 940 => to_unsigned(699, 10), 941 => to_unsigned(574, 10), 942 => to_unsigned(997, 10), 943 => to_unsigned(176, 10), 944 => to_unsigned(485, 10), 945 => to_unsigned(835, 10), 946 => to_unsigned(371, 10), 947 => to_unsigned(121, 10), 948 => to_unsigned(1002, 10), 949 => to_unsigned(757, 10), 950 => to_unsigned(783, 10), 951 => to_unsigned(84, 10), 952 => to_unsigned(7, 10), 953 => to_unsigned(113, 10), 954 => to_unsigned(474, 10), 955 => to_unsigned(974, 10), 956 => to_unsigned(489, 10), 957 => to_unsigned(152, 10), 958 => to_unsigned(242, 10), 959 => to_unsigned(72, 10), 960 => to_unsigned(118, 10), 961 => to_unsigned(949, 10), 962 => to_unsigned(16, 10), 963 => to_unsigned(186, 10), 964 => to_unsigned(639, 10), 965 => to_unsigned(200, 10), 966 => to_unsigned(188, 10), 967 => to_unsigned(716, 10), 968 => to_unsigned(35, 10), 969 => to_unsigned(933, 10), 970 => to_unsigned(585, 10), 971 => to_unsigned(411, 10), 972 => to_unsigned(705, 10), 973 => to_unsigned(316, 10), 974 => to_unsigned(653, 10), 975 => to_unsigned(286, 10), 976 => to_unsigned(669, 10), 977 => to_unsigned(188, 10), 978 => to_unsigned(790, 10), 979 => to_unsigned(118, 10), 980 => to_unsigned(702, 10), 981 => to_unsigned(831, 10), 982 => to_unsigned(940, 10), 983 => to_unsigned(576, 10), 984 => to_unsigned(744, 10), 985 => to_unsigned(629, 10), 986 => to_unsigned(280, 10), 987 => to_unsigned(807, 10), 988 => to_unsigned(810, 10), 989 => to_unsigned(944, 10), 990 => to_unsigned(234, 10), 991 => to_unsigned(944, 10), 992 => to_unsigned(494, 10), 993 => to_unsigned(610, 10), 994 => to_unsigned(935, 10), 995 => to_unsigned(274, 10), 996 => to_unsigned(478, 10), 997 => to_unsigned(269, 10), 998 => to_unsigned(885, 10), 999 => to_unsigned(637, 10), 1000 => to_unsigned(27, 10), 1001 => to_unsigned(179, 10), 1002 => to_unsigned(664, 10), 1003 => to_unsigned(867, 10), 1004 => to_unsigned(535, 10), 1005 => to_unsigned(370, 10), 1006 => to_unsigned(312, 10), 1007 => to_unsigned(471, 10), 1008 => to_unsigned(230, 10), 1009 => to_unsigned(146, 10), 1010 => to_unsigned(677, 10), 1011 => to_unsigned(785, 10), 1012 => to_unsigned(440, 10), 1013 => to_unsigned(428, 10), 1014 => to_unsigned(505, 10), 1015 => to_unsigned(654, 10), 1016 => to_unsigned(882, 10), 1017 => to_unsigned(635, 10), 1018 => to_unsigned(312, 10), 1019 => to_unsigned(824, 10), 1020 => to_unsigned(744, 10), 1021 => to_unsigned(573, 10), 1022 => to_unsigned(199, 10), 1023 => to_unsigned(867, 10), 1024 => to_unsigned(456, 10), 1025 => to_unsigned(390, 10), 1026 => to_unsigned(38, 10), 1027 => to_unsigned(567, 10), 1028 => to_unsigned(649, 10), 1029 => to_unsigned(683, 10), 1030 => to_unsigned(774, 10), 1031 => to_unsigned(927, 10), 1032 => to_unsigned(830, 10), 1033 => to_unsigned(710, 10), 1034 => to_unsigned(915, 10), 1035 => to_unsigned(44, 10), 1036 => to_unsigned(555, 10), 1037 => to_unsigned(311, 10), 1038 => to_unsigned(414, 10), 1039 => to_unsigned(751, 10), 1040 => to_unsigned(638, 10), 1041 => to_unsigned(518, 10), 1042 => to_unsigned(241, 10), 1043 => to_unsigned(646, 10), 1044 => to_unsigned(400, 10), 1045 => to_unsigned(358, 10), 1046 => to_unsigned(446, 10), 1047 => to_unsigned(179, 10), 1048 => to_unsigned(203, 10), 1049 => to_unsigned(832, 10), 1050 => to_unsigned(253, 10), 1051 => to_unsigned(387, 10), 1052 => to_unsigned(730, 10), 1053 => to_unsigned(525, 10), 1054 => to_unsigned(79, 10), 1055 => to_unsigned(510, 10), 1056 => to_unsigned(30, 10), 1057 => to_unsigned(847, 10), 1058 => to_unsigned(497, 10), 1059 => to_unsigned(524, 10), 1060 => to_unsigned(639, 10), 1061 => to_unsigned(349, 10), 1062 => to_unsigned(554, 10), 1063 => to_unsigned(689, 10), 1064 => to_unsigned(270, 10), 1065 => to_unsigned(387, 10), 1066 => to_unsigned(58, 10), 1067 => to_unsigned(305, 10), 1068 => to_unsigned(138, 10), 1069 => to_unsigned(569, 10), 1070 => to_unsigned(184, 10), 1071 => to_unsigned(762, 10), 1072 => to_unsigned(976, 10), 1073 => to_unsigned(67, 10), 1074 => to_unsigned(13, 10), 1075 => to_unsigned(135, 10), 1076 => to_unsigned(755, 10), 1077 => to_unsigned(978, 10), 1078 => to_unsigned(879, 10), 1079 => to_unsigned(743, 10), 1080 => to_unsigned(528, 10), 1081 => to_unsigned(541, 10), 1082 => to_unsigned(70, 10), 1083 => to_unsigned(481, 10), 1084 => to_unsigned(565, 10), 1085 => to_unsigned(862, 10), 1086 => to_unsigned(43, 10), 1087 => to_unsigned(129, 10), 1088 => to_unsigned(392, 10), 1089 => to_unsigned(921, 10), 1090 => to_unsigned(446, 10), 1091 => to_unsigned(487, 10), 1092 => to_unsigned(227, 10), 1093 => to_unsigned(59, 10), 1094 => to_unsigned(645, 10), 1095 => to_unsigned(662, 10), 1096 => to_unsigned(251, 10), 1097 => to_unsigned(819, 10), 1098 => to_unsigned(764, 10), 1099 => to_unsigned(389, 10), 1100 => to_unsigned(882, 10), 1101 => to_unsigned(718, 10), 1102 => to_unsigned(868, 10), 1103 => to_unsigned(917, 10), 1104 => to_unsigned(276, 10), 1105 => to_unsigned(901, 10), 1106 => to_unsigned(382, 10), 1107 => to_unsigned(851, 10), 1108 => to_unsigned(782, 10), 1109 => to_unsigned(558, 10), 1110 => to_unsigned(75, 10), 1111 => to_unsigned(46, 10), 1112 => to_unsigned(135, 10), 1113 => to_unsigned(645, 10), 1114 => to_unsigned(914, 10), 1115 => to_unsigned(788, 10), 1116 => to_unsigned(392, 10), 1117 => to_unsigned(273, 10), 1118 => to_unsigned(825, 10), 1119 => to_unsigned(291, 10), 1120 => to_unsigned(437, 10), 1121 => to_unsigned(1020, 10), 1122 => to_unsigned(863, 10), 1123 => to_unsigned(864, 10), 1124 => to_unsigned(18, 10), 1125 => to_unsigned(96, 10), 1126 => to_unsigned(449, 10), 1127 => to_unsigned(740, 10), 1128 => to_unsigned(639, 10), 1129 => to_unsigned(564, 10), 1130 => to_unsigned(187, 10), 1131 => to_unsigned(824, 10), 1132 => to_unsigned(657, 10), 1133 => to_unsigned(295, 10), 1134 => to_unsigned(979, 10), 1135 => to_unsigned(799, 10), 1136 => to_unsigned(682, 10), 1137 => to_unsigned(903, 10), 1138 => to_unsigned(862, 10), 1139 => to_unsigned(324, 10), 1140 => to_unsigned(66, 10), 1141 => to_unsigned(827, 10), 1142 => to_unsigned(961, 10), 1143 => to_unsigned(38, 10), 1144 => to_unsigned(128, 10), 1145 => to_unsigned(502, 10), 1146 => to_unsigned(524, 10), 1147 => to_unsigned(379, 10), 1148 => to_unsigned(693, 10), 1149 => to_unsigned(942, 10), 1150 => to_unsigned(289, 10), 1151 => to_unsigned(729, 10), 1152 => to_unsigned(679, 10), 1153 => to_unsigned(746, 10), 1154 => to_unsigned(470, 10), 1155 => to_unsigned(108, 10), 1156 => to_unsigned(269, 10), 1157 => to_unsigned(775, 10), 1158 => to_unsigned(641, 10), 1159 => to_unsigned(418, 10), 1160 => to_unsigned(531, 10), 1161 => to_unsigned(583, 10), 1162 => to_unsigned(662, 10), 1163 => to_unsigned(543, 10), 1164 => to_unsigned(162, 10), 1165 => to_unsigned(39, 10), 1166 => to_unsigned(732, 10), 1167 => to_unsigned(649, 10), 1168 => to_unsigned(94, 10), 1169 => to_unsigned(903, 10), 1170 => to_unsigned(279, 10), 1171 => to_unsigned(615, 10), 1172 => to_unsigned(635, 10), 1173 => to_unsigned(546, 10), 1174 => to_unsigned(550, 10), 1175 => to_unsigned(329, 10), 1176 => to_unsigned(711, 10), 1177 => to_unsigned(100, 10), 1178 => to_unsigned(791, 10), 1179 => to_unsigned(100, 10), 1180 => to_unsigned(384, 10), 1181 => to_unsigned(171, 10), 1182 => to_unsigned(936, 10), 1183 => to_unsigned(486, 10), 1184 => to_unsigned(956, 10), 1185 => to_unsigned(550, 10), 1186 => to_unsigned(334, 10), 1187 => to_unsigned(233, 10), 1188 => to_unsigned(749, 10), 1189 => to_unsigned(165, 10), 1190 => to_unsigned(307, 10), 1191 => to_unsigned(586, 10), 1192 => to_unsigned(192, 10), 1193 => to_unsigned(734, 10), 1194 => to_unsigned(945, 10), 1195 => to_unsigned(919, 10), 1196 => to_unsigned(726, 10), 1197 => to_unsigned(77, 10), 1198 => to_unsigned(29, 10), 1199 => to_unsigned(669, 10), 1200 => to_unsigned(669, 10), 1201 => to_unsigned(626, 10), 1202 => to_unsigned(837, 10), 1203 => to_unsigned(571, 10), 1204 => to_unsigned(403, 10), 1205 => to_unsigned(384, 10), 1206 => to_unsigned(1001, 10), 1207 => to_unsigned(897, 10), 1208 => to_unsigned(751, 10), 1209 => to_unsigned(213, 10), 1210 => to_unsigned(547, 10), 1211 => to_unsigned(855, 10), 1212 => to_unsigned(236, 10), 1213 => to_unsigned(366, 10), 1214 => to_unsigned(729, 10), 1215 => to_unsigned(702, 10), 1216 => to_unsigned(796, 10), 1217 => to_unsigned(470, 10), 1218 => to_unsigned(397, 10), 1219 => to_unsigned(772, 10), 1220 => to_unsigned(813, 10), 1221 => to_unsigned(602, 10), 1222 => to_unsigned(872, 10), 1223 => to_unsigned(543, 10), 1224 => to_unsigned(603, 10), 1225 => to_unsigned(43, 10), 1226 => to_unsigned(50, 10), 1227 => to_unsigned(1021, 10), 1228 => to_unsigned(140, 10), 1229 => to_unsigned(937, 10), 1230 => to_unsigned(986, 10), 1231 => to_unsigned(206, 10), 1232 => to_unsigned(954, 10), 1233 => to_unsigned(444, 10), 1234 => to_unsigned(255, 10), 1235 => to_unsigned(54, 10), 1236 => to_unsigned(337, 10), 1237 => to_unsigned(594, 10), 1238 => to_unsigned(343, 10), 1239 => to_unsigned(774, 10), 1240 => to_unsigned(316, 10), 1241 => to_unsigned(285, 10), 1242 => to_unsigned(316, 10), 1243 => to_unsigned(868, 10), 1244 => to_unsigned(556, 10), 1245 => to_unsigned(814, 10), 1246 => to_unsigned(18, 10), 1247 => to_unsigned(859, 10), 1248 => to_unsigned(802, 10), 1249 => to_unsigned(615, 10), 1250 => to_unsigned(444, 10), 1251 => to_unsigned(929, 10), 1252 => to_unsigned(386, 10), 1253 => to_unsigned(327, 10), 1254 => to_unsigned(217, 10), 1255 => to_unsigned(704, 10), 1256 => to_unsigned(478, 10), 1257 => to_unsigned(156, 10), 1258 => to_unsigned(786, 10), 1259 => to_unsigned(988, 10), 1260 => to_unsigned(911, 10), 1261 => to_unsigned(89, 10), 1262 => to_unsigned(411, 10), 1263 => to_unsigned(349, 10), 1264 => to_unsigned(667, 10), 1265 => to_unsigned(110, 10), 1266 => to_unsigned(999, 10), 1267 => to_unsigned(765, 10), 1268 => to_unsigned(7, 10), 1269 => to_unsigned(361, 10), 1270 => to_unsigned(682, 10), 1271 => to_unsigned(804, 10), 1272 => to_unsigned(594, 10), 1273 => to_unsigned(801, 10), 1274 => to_unsigned(69, 10), 1275 => to_unsigned(828, 10), 1276 => to_unsigned(989, 10), 1277 => to_unsigned(463, 10), 1278 => to_unsigned(478, 10), 1279 => to_unsigned(718, 10), 1280 => to_unsigned(71, 10), 1281 => to_unsigned(337, 10), 1282 => to_unsigned(134, 10), 1283 => to_unsigned(744, 10), 1284 => to_unsigned(990, 10), 1285 => to_unsigned(0, 10), 1286 => to_unsigned(253, 10), 1287 => to_unsigned(234, 10), 1288 => to_unsigned(759, 10), 1289 => to_unsigned(474, 10), 1290 => to_unsigned(779, 10), 1291 => to_unsigned(824, 10), 1292 => to_unsigned(520, 10), 1293 => to_unsigned(732, 10), 1294 => to_unsigned(638, 10), 1295 => to_unsigned(819, 10), 1296 => to_unsigned(247, 10), 1297 => to_unsigned(593, 10), 1298 => to_unsigned(165, 10), 1299 => to_unsigned(36, 10), 1300 => to_unsigned(1019, 10), 1301 => to_unsigned(294, 10), 1302 => to_unsigned(740, 10), 1303 => to_unsigned(579, 10), 1304 => to_unsigned(192, 10), 1305 => to_unsigned(261, 10), 1306 => to_unsigned(917, 10), 1307 => to_unsigned(308, 10), 1308 => to_unsigned(954, 10), 1309 => to_unsigned(844, 10), 1310 => to_unsigned(723, 10), 1311 => to_unsigned(170, 10), 1312 => to_unsigned(390, 10), 1313 => to_unsigned(0, 10), 1314 => to_unsigned(88, 10), 1315 => to_unsigned(12, 10), 1316 => to_unsigned(55, 10), 1317 => to_unsigned(986, 10), 1318 => to_unsigned(319, 10), 1319 => to_unsigned(571, 10), 1320 => to_unsigned(372, 10), 1321 => to_unsigned(714, 10), 1322 => to_unsigned(546, 10), 1323 => to_unsigned(86, 10), 1324 => to_unsigned(690, 10), 1325 => to_unsigned(313, 10), 1326 => to_unsigned(590, 10), 1327 => to_unsigned(800, 10), 1328 => to_unsigned(219, 10), 1329 => to_unsigned(959, 10), 1330 => to_unsigned(792, 10), 1331 => to_unsigned(799, 10), 1332 => to_unsigned(76, 10), 1333 => to_unsigned(323, 10), 1334 => to_unsigned(858, 10), 1335 => to_unsigned(48, 10), 1336 => to_unsigned(343, 10), 1337 => to_unsigned(826, 10), 1338 => to_unsigned(448, 10), 1339 => to_unsigned(778, 10), 1340 => to_unsigned(285, 10), 1341 => to_unsigned(673, 10), 1342 => to_unsigned(487, 10), 1343 => to_unsigned(923, 10), 1344 => to_unsigned(533, 10), 1345 => to_unsigned(350, 10), 1346 => to_unsigned(847, 10), 1347 => to_unsigned(889, 10), 1348 => to_unsigned(497, 10), 1349 => to_unsigned(1001, 10), 1350 => to_unsigned(200, 10), 1351 => to_unsigned(487, 10), 1352 => to_unsigned(151, 10), 1353 => to_unsigned(419, 10), 1354 => to_unsigned(310, 10), 1355 => to_unsigned(247, 10), 1356 => to_unsigned(435, 10), 1357 => to_unsigned(946, 10), 1358 => to_unsigned(280, 10), 1359 => to_unsigned(282, 10), 1360 => to_unsigned(540, 10), 1361 => to_unsigned(78, 10), 1362 => to_unsigned(974, 10), 1363 => to_unsigned(123, 10), 1364 => to_unsigned(468, 10), 1365 => to_unsigned(942, 10), 1366 => to_unsigned(806, 10), 1367 => to_unsigned(451, 10), 1368 => to_unsigned(911, 10), 1369 => to_unsigned(279, 10), 1370 => to_unsigned(484, 10), 1371 => to_unsigned(254, 10), 1372 => to_unsigned(189, 10), 1373 => to_unsigned(216, 10), 1374 => to_unsigned(977, 10), 1375 => to_unsigned(862, 10), 1376 => to_unsigned(977, 10), 1377 => to_unsigned(145, 10), 1378 => to_unsigned(314, 10), 1379 => to_unsigned(678, 10), 1380 => to_unsigned(435, 10), 1381 => to_unsigned(80, 10), 1382 => to_unsigned(47, 10), 1383 => to_unsigned(778, 10), 1384 => to_unsigned(389, 10), 1385 => to_unsigned(194, 10), 1386 => to_unsigned(782, 10), 1387 => to_unsigned(741, 10), 1388 => to_unsigned(308, 10), 1389 => to_unsigned(448, 10), 1390 => to_unsigned(541, 10), 1391 => to_unsigned(916, 10), 1392 => to_unsigned(965, 10), 1393 => to_unsigned(259, 10), 1394 => to_unsigned(1012, 10), 1395 => to_unsigned(970, 10), 1396 => to_unsigned(462, 10), 1397 => to_unsigned(261, 10), 1398 => to_unsigned(406, 10), 1399 => to_unsigned(67, 10), 1400 => to_unsigned(780, 10), 1401 => to_unsigned(876, 10), 1402 => to_unsigned(512, 10), 1403 => to_unsigned(160, 10), 1404 => to_unsigned(38, 10), 1405 => to_unsigned(636, 10), 1406 => to_unsigned(196, 10), 1407 => to_unsigned(984, 10), 1408 => to_unsigned(734, 10), 1409 => to_unsigned(884, 10), 1410 => to_unsigned(296, 10), 1411 => to_unsigned(126, 10), 1412 => to_unsigned(68, 10), 1413 => to_unsigned(906, 10), 1414 => to_unsigned(732, 10), 1415 => to_unsigned(797, 10), 1416 => to_unsigned(656, 10), 1417 => to_unsigned(468, 10), 1418 => to_unsigned(16, 10), 1419 => to_unsigned(459, 10), 1420 => to_unsigned(852, 10), 1421 => to_unsigned(137, 10), 1422 => to_unsigned(661, 10), 1423 => to_unsigned(638, 10), 1424 => to_unsigned(82, 10), 1425 => to_unsigned(78, 10), 1426 => to_unsigned(375, 10), 1427 => to_unsigned(951, 10), 1428 => to_unsigned(27, 10), 1429 => to_unsigned(639, 10), 1430 => to_unsigned(425, 10), 1431 => to_unsigned(499, 10), 1432 => to_unsigned(457, 10), 1433 => to_unsigned(291, 10), 1434 => to_unsigned(959, 10), 1435 => to_unsigned(503, 10), 1436 => to_unsigned(83, 10), 1437 => to_unsigned(826, 10), 1438 => to_unsigned(10, 10), 1439 => to_unsigned(565, 10), 1440 => to_unsigned(704, 10), 1441 => to_unsigned(662, 10), 1442 => to_unsigned(998, 10), 1443 => to_unsigned(427, 10), 1444 => to_unsigned(894, 10), 1445 => to_unsigned(968, 10), 1446 => to_unsigned(203, 10), 1447 => to_unsigned(93, 10), 1448 => to_unsigned(668, 10), 1449 => to_unsigned(692, 10), 1450 => to_unsigned(128, 10), 1451 => to_unsigned(961, 10), 1452 => to_unsigned(81, 10), 1453 => to_unsigned(12, 10), 1454 => to_unsigned(44, 10), 1455 => to_unsigned(991, 10), 1456 => to_unsigned(691, 10), 1457 => to_unsigned(739, 10), 1458 => to_unsigned(873, 10), 1459 => to_unsigned(266, 10), 1460 => to_unsigned(761, 10), 1461 => to_unsigned(700, 10), 1462 => to_unsigned(617, 10), 1463 => to_unsigned(172, 10), 1464 => to_unsigned(659, 10), 1465 => to_unsigned(61, 10), 1466 => to_unsigned(434, 10), 1467 => to_unsigned(442, 10), 1468 => to_unsigned(629, 10), 1469 => to_unsigned(828, 10), 1470 => to_unsigned(890, 10), 1471 => to_unsigned(108, 10), 1472 => to_unsigned(403, 10), 1473 => to_unsigned(742, 10), 1474 => to_unsigned(201, 10), 1475 => to_unsigned(781, 10), 1476 => to_unsigned(590, 10), 1477 => to_unsigned(837, 10), 1478 => to_unsigned(243, 10), 1479 => to_unsigned(493, 10), 1480 => to_unsigned(243, 10), 1481 => to_unsigned(241, 10), 1482 => to_unsigned(186, 10), 1483 => to_unsigned(628, 10), 1484 => to_unsigned(723, 10), 1485 => to_unsigned(683, 10), 1486 => to_unsigned(124, 10), 1487 => to_unsigned(97, 10), 1488 => to_unsigned(804, 10), 1489 => to_unsigned(364, 10), 1490 => to_unsigned(739, 10), 1491 => to_unsigned(884, 10), 1492 => to_unsigned(670, 10), 1493 => to_unsigned(184, 10), 1494 => to_unsigned(248, 10), 1495 => to_unsigned(512, 10), 1496 => to_unsigned(925, 10), 1497 => to_unsigned(763, 10), 1498 => to_unsigned(371, 10), 1499 => to_unsigned(617, 10), 1500 => to_unsigned(353, 10), 1501 => to_unsigned(523, 10), 1502 => to_unsigned(817, 10), 1503 => to_unsigned(554, 10), 1504 => to_unsigned(261, 10), 1505 => to_unsigned(393, 10), 1506 => to_unsigned(411, 10), 1507 => to_unsigned(686, 10), 1508 => to_unsigned(171, 10), 1509 => to_unsigned(527, 10), 1510 => to_unsigned(447, 10), 1511 => to_unsigned(931, 10), 1512 => to_unsigned(10, 10), 1513 => to_unsigned(903, 10), 1514 => to_unsigned(526, 10), 1515 => to_unsigned(592, 10), 1516 => to_unsigned(163, 10), 1517 => to_unsigned(138, 10), 1518 => to_unsigned(492, 10), 1519 => to_unsigned(134, 10), 1520 => to_unsigned(539, 10), 1521 => to_unsigned(753, 10), 1522 => to_unsigned(239, 10), 1523 => to_unsigned(758, 10), 1524 => to_unsigned(918, 10), 1525 => to_unsigned(223, 10), 1526 => to_unsigned(50, 10), 1527 => to_unsigned(140, 10), 1528 => to_unsigned(127, 10), 1529 => to_unsigned(441, 10), 1530 => to_unsigned(290, 10), 1531 => to_unsigned(856, 10), 1532 => to_unsigned(1009, 10), 1533 => to_unsigned(298, 10), 1534 => to_unsigned(462, 10), 1535 => to_unsigned(496, 10), 1536 => to_unsigned(720, 10), 1537 => to_unsigned(622, 10), 1538 => to_unsigned(689, 10), 1539 => to_unsigned(660, 10), 1540 => to_unsigned(665, 10), 1541 => to_unsigned(784, 10), 1542 => to_unsigned(242, 10), 1543 => to_unsigned(998, 10), 1544 => to_unsigned(174, 10), 1545 => to_unsigned(704, 10), 1546 => to_unsigned(497, 10), 1547 => to_unsigned(853, 10), 1548 => to_unsigned(360, 10), 1549 => to_unsigned(412, 10), 1550 => to_unsigned(453, 10), 1551 => to_unsigned(352, 10), 1552 => to_unsigned(844, 10), 1553 => to_unsigned(476, 10), 1554 => to_unsigned(202, 10), 1555 => to_unsigned(248, 10), 1556 => to_unsigned(970, 10), 1557 => to_unsigned(251, 10), 1558 => to_unsigned(314, 10), 1559 => to_unsigned(922, 10), 1560 => to_unsigned(439, 10), 1561 => to_unsigned(132, 10), 1562 => to_unsigned(1012, 10), 1563 => to_unsigned(763, 10), 1564 => to_unsigned(709, 10), 1565 => to_unsigned(84, 10), 1566 => to_unsigned(196, 10), 1567 => to_unsigned(530, 10), 1568 => to_unsigned(412, 10), 1569 => to_unsigned(104, 10), 1570 => to_unsigned(955, 10), 1571 => to_unsigned(860, 10), 1572 => to_unsigned(321, 10), 1573 => to_unsigned(514, 10), 1574 => to_unsigned(605, 10), 1575 => to_unsigned(175, 10), 1576 => to_unsigned(362, 10), 1577 => to_unsigned(320, 10), 1578 => to_unsigned(327, 10), 1579 => to_unsigned(369, 10), 1580 => to_unsigned(197, 10), 1581 => to_unsigned(411, 10), 1582 => to_unsigned(962, 10), 1583 => to_unsigned(960, 10), 1584 => to_unsigned(388, 10), 1585 => to_unsigned(843, 10), 1586 => to_unsigned(682, 10), 1587 => to_unsigned(415, 10), 1588 => to_unsigned(476, 10), 1589 => to_unsigned(84, 10), 1590 => to_unsigned(168, 10), 1591 => to_unsigned(773, 10), 1592 => to_unsigned(100, 10), 1593 => to_unsigned(451, 10), 1594 => to_unsigned(535, 10), 1595 => to_unsigned(157, 10), 1596 => to_unsigned(884, 10), 1597 => to_unsigned(861, 10), 1598 => to_unsigned(290, 10), 1599 => to_unsigned(727, 10), 1600 => to_unsigned(189, 10), 1601 => to_unsigned(38, 10), 1602 => to_unsigned(435, 10), 1603 => to_unsigned(491, 10), 1604 => to_unsigned(567, 10), 1605 => to_unsigned(608, 10), 1606 => to_unsigned(327, 10), 1607 => to_unsigned(80, 10), 1608 => to_unsigned(360, 10), 1609 => to_unsigned(793, 10), 1610 => to_unsigned(430, 10), 1611 => to_unsigned(305, 10), 1612 => to_unsigned(176, 10), 1613 => to_unsigned(910, 10), 1614 => to_unsigned(68, 10), 1615 => to_unsigned(958, 10), 1616 => to_unsigned(132, 10), 1617 => to_unsigned(155, 10), 1618 => to_unsigned(253, 10), 1619 => to_unsigned(940, 10), 1620 => to_unsigned(68, 10), 1621 => to_unsigned(134, 10), 1622 => to_unsigned(938, 10), 1623 => to_unsigned(507, 10), 1624 => to_unsigned(152, 10), 1625 => to_unsigned(312, 10), 1626 => to_unsigned(308, 10), 1627 => to_unsigned(559, 10), 1628 => to_unsigned(816, 10), 1629 => to_unsigned(887, 10), 1630 => to_unsigned(159, 10), 1631 => to_unsigned(536, 10), 1632 => to_unsigned(212, 10), 1633 => to_unsigned(751, 10), 1634 => to_unsigned(493, 10), 1635 => to_unsigned(102, 10), 1636 => to_unsigned(438, 10), 1637 => to_unsigned(132, 10), 1638 => to_unsigned(422, 10), 1639 => to_unsigned(1000, 10), 1640 => to_unsigned(442, 10), 1641 => to_unsigned(315, 10), 1642 => to_unsigned(413, 10), 1643 => to_unsigned(122, 10), 1644 => to_unsigned(62, 10), 1645 => to_unsigned(612, 10), 1646 => to_unsigned(387, 10), 1647 => to_unsigned(898, 10), 1648 => to_unsigned(897, 10), 1649 => to_unsigned(178, 10), 1650 => to_unsigned(398, 10), 1651 => to_unsigned(1015, 10), 1652 => to_unsigned(230, 10), 1653 => to_unsigned(157, 10), 1654 => to_unsigned(997, 10), 1655 => to_unsigned(741, 10), 1656 => to_unsigned(445, 10), 1657 => to_unsigned(664, 10), 1658 => to_unsigned(663, 10), 1659 => to_unsigned(472, 10), 1660 => to_unsigned(808, 10), 1661 => to_unsigned(900, 10), 1662 => to_unsigned(910, 10), 1663 => to_unsigned(320, 10), 1664 => to_unsigned(795, 10), 1665 => to_unsigned(130, 10), 1666 => to_unsigned(938, 10), 1667 => to_unsigned(628, 10), 1668 => to_unsigned(475, 10), 1669 => to_unsigned(335, 10), 1670 => to_unsigned(471, 10), 1671 => to_unsigned(915, 10), 1672 => to_unsigned(195, 10), 1673 => to_unsigned(873, 10), 1674 => to_unsigned(408, 10), 1675 => to_unsigned(361, 10), 1676 => to_unsigned(118, 10), 1677 => to_unsigned(978, 10), 1678 => to_unsigned(38, 10), 1679 => to_unsigned(364, 10), 1680 => to_unsigned(395, 10), 1681 => to_unsigned(128, 10), 1682 => to_unsigned(49, 10), 1683 => to_unsigned(365, 10), 1684 => to_unsigned(113, 10), 1685 => to_unsigned(800, 10), 1686 => to_unsigned(478, 10), 1687 => to_unsigned(901, 10), 1688 => to_unsigned(125, 10), 1689 => to_unsigned(242, 10), 1690 => to_unsigned(509, 10), 1691 => to_unsigned(182, 10), 1692 => to_unsigned(0, 10), 1693 => to_unsigned(186, 10), 1694 => to_unsigned(27, 10), 1695 => to_unsigned(563, 10), 1696 => to_unsigned(490, 10), 1697 => to_unsigned(890, 10), 1698 => to_unsigned(958, 10), 1699 => to_unsigned(622, 10), 1700 => to_unsigned(829, 10), 1701 => to_unsigned(363, 10), 1702 => to_unsigned(606, 10), 1703 => to_unsigned(588, 10), 1704 => to_unsigned(955, 10), 1705 => to_unsigned(550, 10), 1706 => to_unsigned(430, 10), 1707 => to_unsigned(287, 10), 1708 => to_unsigned(758, 10), 1709 => to_unsigned(178, 10), 1710 => to_unsigned(549, 10), 1711 => to_unsigned(807, 10), 1712 => to_unsigned(108, 10), 1713 => to_unsigned(115, 10), 1714 => to_unsigned(478, 10), 1715 => to_unsigned(369, 10), 1716 => to_unsigned(896, 10), 1717 => to_unsigned(689, 10), 1718 => to_unsigned(640, 10), 1719 => to_unsigned(357, 10), 1720 => to_unsigned(497, 10), 1721 => to_unsigned(1015, 10), 1722 => to_unsigned(188, 10), 1723 => to_unsigned(107, 10), 1724 => to_unsigned(538, 10), 1725 => to_unsigned(740, 10), 1726 => to_unsigned(105, 10), 1727 => to_unsigned(960, 10), 1728 => to_unsigned(559, 10), 1729 => to_unsigned(564, 10), 1730 => to_unsigned(36, 10), 1731 => to_unsigned(215, 10), 1732 => to_unsigned(233, 10), 1733 => to_unsigned(57, 10), 1734 => to_unsigned(99, 10), 1735 => to_unsigned(410, 10), 1736 => to_unsigned(55, 10), 1737 => to_unsigned(825, 10), 1738 => to_unsigned(466, 10), 1739 => to_unsigned(661, 10), 1740 => to_unsigned(878, 10), 1741 => to_unsigned(1020, 10), 1742 => to_unsigned(765, 10), 1743 => to_unsigned(382, 10), 1744 => to_unsigned(453, 10), 1745 => to_unsigned(611, 10), 1746 => to_unsigned(54, 10), 1747 => to_unsigned(84, 10), 1748 => to_unsigned(149, 10), 1749 => to_unsigned(1020, 10), 1750 => to_unsigned(596, 10), 1751 => to_unsigned(1004, 10), 1752 => to_unsigned(627, 10), 1753 => to_unsigned(424, 10), 1754 => to_unsigned(375, 10), 1755 => to_unsigned(526, 10), 1756 => to_unsigned(69, 10), 1757 => to_unsigned(744, 10), 1758 => to_unsigned(658, 10), 1759 => to_unsigned(674, 10), 1760 => to_unsigned(536, 10), 1761 => to_unsigned(970, 10), 1762 => to_unsigned(782, 10), 1763 => to_unsigned(202, 10), 1764 => to_unsigned(271, 10), 1765 => to_unsigned(663, 10), 1766 => to_unsigned(873, 10), 1767 => to_unsigned(833, 10), 1768 => to_unsigned(702, 10), 1769 => to_unsigned(543, 10), 1770 => to_unsigned(896, 10), 1771 => to_unsigned(556, 10), 1772 => to_unsigned(694, 10), 1773 => to_unsigned(67, 10), 1774 => to_unsigned(321, 10), 1775 => to_unsigned(246, 10), 1776 => to_unsigned(360, 10), 1777 => to_unsigned(509, 10), 1778 => to_unsigned(296, 10), 1779 => to_unsigned(635, 10), 1780 => to_unsigned(536, 10), 1781 => to_unsigned(95, 10), 1782 => to_unsigned(27, 10), 1783 => to_unsigned(550, 10), 1784 => to_unsigned(305, 10), 1785 => to_unsigned(723, 10), 1786 => to_unsigned(922, 10), 1787 => to_unsigned(140, 10), 1788 => to_unsigned(341, 10), 1789 => to_unsigned(825, 10), 1790 => to_unsigned(919, 10), 1791 => to_unsigned(425, 10), 1792 => to_unsigned(673, 10), 1793 => to_unsigned(156, 10), 1794 => to_unsigned(940, 10), 1795 => to_unsigned(726, 10), 1796 => to_unsigned(75, 10), 1797 => to_unsigned(3, 10), 1798 => to_unsigned(750, 10), 1799 => to_unsigned(386, 10), 1800 => to_unsigned(691, 10), 1801 => to_unsigned(859, 10), 1802 => to_unsigned(742, 10), 1803 => to_unsigned(490, 10), 1804 => to_unsigned(250, 10), 1805 => to_unsigned(739, 10), 1806 => to_unsigned(855, 10), 1807 => to_unsigned(578, 10), 1808 => to_unsigned(65, 10), 1809 => to_unsigned(448, 10), 1810 => to_unsigned(1014, 10), 1811 => to_unsigned(248, 10), 1812 => to_unsigned(950, 10), 1813 => to_unsigned(620, 10), 1814 => to_unsigned(703, 10), 1815 => to_unsigned(740, 10), 1816 => to_unsigned(281, 10), 1817 => to_unsigned(925, 10), 1818 => to_unsigned(865, 10), 1819 => to_unsigned(218, 10), 1820 => to_unsigned(55, 10), 1821 => to_unsigned(202, 10), 1822 => to_unsigned(918, 10), 1823 => to_unsigned(245, 10), 1824 => to_unsigned(195, 10), 1825 => to_unsigned(484, 10), 1826 => to_unsigned(499, 10), 1827 => to_unsigned(424, 10), 1828 => to_unsigned(744, 10), 1829 => to_unsigned(751, 10), 1830 => to_unsigned(318, 10), 1831 => to_unsigned(538, 10), 1832 => to_unsigned(694, 10), 1833 => to_unsigned(692, 10), 1834 => to_unsigned(127, 10), 1835 => to_unsigned(81, 10), 1836 => to_unsigned(892, 10), 1837 => to_unsigned(745, 10), 1838 => to_unsigned(679, 10), 1839 => to_unsigned(443, 10), 1840 => to_unsigned(937, 10), 1841 => to_unsigned(525, 10), 1842 => to_unsigned(698, 10), 1843 => to_unsigned(188, 10), 1844 => to_unsigned(969, 10), 1845 => to_unsigned(821, 10), 1846 => to_unsigned(901, 10), 1847 => to_unsigned(859, 10), 1848 => to_unsigned(94, 10), 1849 => to_unsigned(601, 10), 1850 => to_unsigned(99, 10), 1851 => to_unsigned(447, 10), 1852 => to_unsigned(185, 10), 1853 => to_unsigned(624, 10), 1854 => to_unsigned(674, 10), 1855 => to_unsigned(967, 10), 1856 => to_unsigned(367, 10), 1857 => to_unsigned(925, 10), 1858 => to_unsigned(815, 10), 1859 => to_unsigned(684, 10), 1860 => to_unsigned(490, 10), 1861 => to_unsigned(412, 10), 1862 => to_unsigned(513, 10), 1863 => to_unsigned(762, 10), 1864 => to_unsigned(128, 10), 1865 => to_unsigned(945, 10), 1866 => to_unsigned(776, 10), 1867 => to_unsigned(457, 10), 1868 => to_unsigned(299, 10), 1869 => to_unsigned(932, 10), 1870 => to_unsigned(732, 10), 1871 => to_unsigned(221, 10), 1872 => to_unsigned(288, 10), 1873 => to_unsigned(368, 10), 1874 => to_unsigned(631, 10), 1875 => to_unsigned(640, 10), 1876 => to_unsigned(59, 10), 1877 => to_unsigned(969, 10), 1878 => to_unsigned(42, 10), 1879 => to_unsigned(0, 10), 1880 => to_unsigned(1015, 10), 1881 => to_unsigned(302, 10), 1882 => to_unsigned(288, 10), 1883 => to_unsigned(253, 10), 1884 => to_unsigned(987, 10), 1885 => to_unsigned(165, 10), 1886 => to_unsigned(618, 10), 1887 => to_unsigned(124, 10), 1888 => to_unsigned(869, 10), 1889 => to_unsigned(919, 10), 1890 => to_unsigned(488, 10), 1891 => to_unsigned(276, 10), 1892 => to_unsigned(136, 10), 1893 => to_unsigned(681, 10), 1894 => to_unsigned(398, 10), 1895 => to_unsigned(448, 10), 1896 => to_unsigned(592, 10), 1897 => to_unsigned(1013, 10), 1898 => to_unsigned(976, 10), 1899 => to_unsigned(435, 10), 1900 => to_unsigned(271, 10), 1901 => to_unsigned(395, 10), 1902 => to_unsigned(432, 10), 1903 => to_unsigned(907, 10), 1904 => to_unsigned(835, 10), 1905 => to_unsigned(354, 10), 1906 => to_unsigned(568, 10), 1907 => to_unsigned(630, 10), 1908 => to_unsigned(451, 10), 1909 => to_unsigned(332, 10), 1910 => to_unsigned(852, 10), 1911 => to_unsigned(418, 10), 1912 => to_unsigned(813, 10), 1913 => to_unsigned(655, 10), 1914 => to_unsigned(1015, 10), 1915 => to_unsigned(17, 10), 1916 => to_unsigned(972, 10), 1917 => to_unsigned(314, 10), 1918 => to_unsigned(23, 10), 1919 => to_unsigned(77, 10), 1920 => to_unsigned(355, 10), 1921 => to_unsigned(463, 10), 1922 => to_unsigned(289, 10), 1923 => to_unsigned(313, 10), 1924 => to_unsigned(73, 10), 1925 => to_unsigned(199, 10), 1926 => to_unsigned(693, 10), 1927 => to_unsigned(500, 10), 1928 => to_unsigned(289, 10), 1929 => to_unsigned(800, 10), 1930 => to_unsigned(15, 10), 1931 => to_unsigned(771, 10), 1932 => to_unsigned(283, 10), 1933 => to_unsigned(165, 10), 1934 => to_unsigned(878, 10), 1935 => to_unsigned(985, 10), 1936 => to_unsigned(305, 10), 1937 => to_unsigned(47, 10), 1938 => to_unsigned(121, 10), 1939 => to_unsigned(1006, 10), 1940 => to_unsigned(219, 10), 1941 => to_unsigned(497, 10), 1942 => to_unsigned(729, 10), 1943 => to_unsigned(235, 10), 1944 => to_unsigned(258, 10), 1945 => to_unsigned(950, 10), 1946 => to_unsigned(523, 10), 1947 => to_unsigned(882, 10), 1948 => to_unsigned(236, 10), 1949 => to_unsigned(780, 10), 1950 => to_unsigned(202, 10), 1951 => to_unsigned(107, 10), 1952 => to_unsigned(1006, 10), 1953 => to_unsigned(207, 10), 1954 => to_unsigned(832, 10), 1955 => to_unsigned(715, 10), 1956 => to_unsigned(11, 10), 1957 => to_unsigned(527, 10), 1958 => to_unsigned(935, 10), 1959 => to_unsigned(82, 10), 1960 => to_unsigned(950, 10), 1961 => to_unsigned(573, 10), 1962 => to_unsigned(312, 10), 1963 => to_unsigned(112, 10), 1964 => to_unsigned(364, 10), 1965 => to_unsigned(239, 10), 1966 => to_unsigned(432, 10), 1967 => to_unsigned(242, 10), 1968 => to_unsigned(762, 10), 1969 => to_unsigned(799, 10), 1970 => to_unsigned(576, 10), 1971 => to_unsigned(248, 10), 1972 => to_unsigned(547, 10), 1973 => to_unsigned(458, 10), 1974 => to_unsigned(849, 10), 1975 => to_unsigned(734, 10), 1976 => to_unsigned(291, 10), 1977 => to_unsigned(46, 10), 1978 => to_unsigned(90, 10), 1979 => to_unsigned(871, 10), 1980 => to_unsigned(346, 10), 1981 => to_unsigned(332, 10), 1982 => to_unsigned(421, 10), 1983 => to_unsigned(851, 10), 1984 => to_unsigned(582, 10), 1985 => to_unsigned(90, 10), 1986 => to_unsigned(566, 10), 1987 => to_unsigned(67, 10), 1988 => to_unsigned(666, 10), 1989 => to_unsigned(898, 10), 1990 => to_unsigned(297, 10), 1991 => to_unsigned(580, 10), 1992 => to_unsigned(747, 10), 1993 => to_unsigned(842, 10), 1994 => to_unsigned(627, 10), 1995 => to_unsigned(867, 10), 1996 => to_unsigned(543, 10), 1997 => to_unsigned(712, 10), 1998 => to_unsigned(294, 10), 1999 => to_unsigned(787, 10), 2000 => to_unsigned(656, 10), 2001 => to_unsigned(339, 10), 2002 => to_unsigned(99, 10), 2003 => to_unsigned(783, 10), 2004 => to_unsigned(320, 10), 2005 => to_unsigned(751, 10), 2006 => to_unsigned(444, 10), 2007 => to_unsigned(582, 10), 2008 => to_unsigned(270, 10), 2009 => to_unsigned(1019, 10), 2010 => to_unsigned(166, 10), 2011 => to_unsigned(786, 10), 2012 => to_unsigned(308, 10), 2013 => to_unsigned(478, 10), 2014 => to_unsigned(793, 10), 2015 => to_unsigned(347, 10), 2016 => to_unsigned(169, 10), 2017 => to_unsigned(876, 10), 2018 => to_unsigned(314, 10), 2019 => to_unsigned(294, 10), 2020 => to_unsigned(635, 10), 2021 => to_unsigned(176, 10), 2022 => to_unsigned(983, 10), 2023 => to_unsigned(41, 10), 2024 => to_unsigned(488, 10), 2025 => to_unsigned(438, 10), 2026 => to_unsigned(724, 10), 2027 => to_unsigned(331, 10), 2028 => to_unsigned(731, 10), 2029 => to_unsigned(853, 10), 2030 => to_unsigned(385, 10), 2031 => to_unsigned(905, 10), 2032 => to_unsigned(86, 10), 2033 => to_unsigned(242, 10), 2034 => to_unsigned(396, 10), 2035 => to_unsigned(225, 10), 2036 => to_unsigned(176, 10), 2037 => to_unsigned(693, 10), 2038 => to_unsigned(750, 10), 2039 => to_unsigned(837, 10), 2040 => to_unsigned(568, 10), 2041 => to_unsigned(955, 10), 2042 => to_unsigned(604, 10), 2043 => to_unsigned(797, 10), 2044 => to_unsigned(130, 10), 2045 => to_unsigned(381, 10), 2046 => to_unsigned(30, 10), 2047 => to_unsigned(290, 10))
        ),
        1 => (
            0 => (0 => to_unsigned(570, 10), 1 => to_unsigned(241, 10), 2 => to_unsigned(332, 10), 3 => to_unsigned(597, 10), 4 => to_unsigned(972, 10), 5 => to_unsigned(80, 10), 6 => to_unsigned(599, 10), 7 => to_unsigned(714, 10), 8 => to_unsigned(848, 10), 9 => to_unsigned(85, 10), 10 => to_unsigned(89, 10), 11 => to_unsigned(19, 10), 12 => to_unsigned(482, 10), 13 => to_unsigned(919, 10), 14 => to_unsigned(144, 10), 15 => to_unsigned(364, 10), 16 => to_unsigned(672, 10), 17 => to_unsigned(577, 10), 18 => to_unsigned(346, 10), 19 => to_unsigned(525, 10), 20 => to_unsigned(286, 10), 21 => to_unsigned(163, 10), 22 => to_unsigned(1001, 10), 23 => to_unsigned(300, 10), 24 => to_unsigned(543, 10), 25 => to_unsigned(169, 10), 26 => to_unsigned(952, 10), 27 => to_unsigned(470, 10), 28 => to_unsigned(513, 10), 29 => to_unsigned(510, 10), 30 => to_unsigned(767, 10), 31 => to_unsigned(399, 10), 32 => to_unsigned(415, 10), 33 => to_unsigned(126, 10), 34 => to_unsigned(322, 10), 35 => to_unsigned(717, 10), 36 => to_unsigned(512, 10), 37 => to_unsigned(768, 10), 38 => to_unsigned(10, 10), 39 => to_unsigned(784, 10), 40 => to_unsigned(760, 10), 41 => to_unsigned(523, 10), 42 => to_unsigned(444, 10), 43 => to_unsigned(985, 10), 44 => to_unsigned(278, 10), 45 => to_unsigned(255, 10), 46 => to_unsigned(575, 10), 47 => to_unsigned(837, 10), 48 => to_unsigned(323, 10), 49 => to_unsigned(622, 10), 50 => to_unsigned(252, 10), 51 => to_unsigned(275, 10), 52 => to_unsigned(582, 10), 53 => to_unsigned(307, 10), 54 => to_unsigned(401, 10), 55 => to_unsigned(311, 10), 56 => to_unsigned(400, 10), 57 => to_unsigned(921, 10), 58 => to_unsigned(508, 10), 59 => to_unsigned(482, 10), 60 => to_unsigned(182, 10), 61 => to_unsigned(169, 10), 62 => to_unsigned(977, 10), 63 => to_unsigned(876, 10), 64 => to_unsigned(408, 10), 65 => to_unsigned(266, 10), 66 => to_unsigned(626, 10), 67 => to_unsigned(362, 10), 68 => to_unsigned(282, 10), 69 => to_unsigned(1019, 10), 70 => to_unsigned(55, 10), 71 => to_unsigned(247, 10), 72 => to_unsigned(612, 10), 73 => to_unsigned(380, 10), 74 => to_unsigned(222, 10), 75 => to_unsigned(880, 10), 76 => to_unsigned(722, 10), 77 => to_unsigned(640, 10), 78 => to_unsigned(3, 10), 79 => to_unsigned(190, 10), 80 => to_unsigned(98, 10), 81 => to_unsigned(796, 10), 82 => to_unsigned(511, 10), 83 => to_unsigned(767, 10), 84 => to_unsigned(906, 10), 85 => to_unsigned(593, 10), 86 => to_unsigned(584, 10), 87 => to_unsigned(957, 10), 88 => to_unsigned(917, 10), 89 => to_unsigned(431, 10), 90 => to_unsigned(603, 10), 91 => to_unsigned(78, 10), 92 => to_unsigned(408, 10), 93 => to_unsigned(850, 10), 94 => to_unsigned(802, 10), 95 => to_unsigned(1007, 10), 96 => to_unsigned(1018, 10), 97 => to_unsigned(887, 10), 98 => to_unsigned(979, 10), 99 => to_unsigned(367, 10), 100 => to_unsigned(604, 10), 101 => to_unsigned(971, 10), 102 => to_unsigned(722, 10), 103 => to_unsigned(832, 10), 104 => to_unsigned(422, 10), 105 => to_unsigned(234, 10), 106 => to_unsigned(1007, 10), 107 => to_unsigned(45, 10), 108 => to_unsigned(292, 10), 109 => to_unsigned(513, 10), 110 => to_unsigned(40, 10), 111 => to_unsigned(364, 10), 112 => to_unsigned(95, 10), 113 => to_unsigned(875, 10), 114 => to_unsigned(625, 10), 115 => to_unsigned(352, 10), 116 => to_unsigned(408, 10), 117 => to_unsigned(192, 10), 118 => to_unsigned(157, 10), 119 => to_unsigned(958, 10), 120 => to_unsigned(503, 10), 121 => to_unsigned(108, 10), 122 => to_unsigned(226, 10), 123 => to_unsigned(495, 10), 124 => to_unsigned(1010, 10), 125 => to_unsigned(1004, 10), 126 => to_unsigned(684, 10), 127 => to_unsigned(322, 10), 128 => to_unsigned(530, 10), 129 => to_unsigned(717, 10), 130 => to_unsigned(501, 10), 131 => to_unsigned(200, 10), 132 => to_unsigned(516, 10), 133 => to_unsigned(275, 10), 134 => to_unsigned(905, 10), 135 => to_unsigned(93, 10), 136 => to_unsigned(576, 10), 137 => to_unsigned(294, 10), 138 => to_unsigned(1009, 10), 139 => to_unsigned(534, 10), 140 => to_unsigned(921, 10), 141 => to_unsigned(539, 10), 142 => to_unsigned(657, 10), 143 => to_unsigned(701, 10), 144 => to_unsigned(698, 10), 145 => to_unsigned(246, 10), 146 => to_unsigned(345, 10), 147 => to_unsigned(118, 10), 148 => to_unsigned(118, 10), 149 => to_unsigned(107, 10), 150 => to_unsigned(971, 10), 151 => to_unsigned(454, 10), 152 => to_unsigned(324, 10), 153 => to_unsigned(670, 10), 154 => to_unsigned(648, 10), 155 => to_unsigned(828, 10), 156 => to_unsigned(655, 10), 157 => to_unsigned(531, 10), 158 => to_unsigned(144, 10), 159 => to_unsigned(480, 10), 160 => to_unsigned(860, 10), 161 => to_unsigned(266, 10), 162 => to_unsigned(698, 10), 163 => to_unsigned(157, 10), 164 => to_unsigned(717, 10), 165 => to_unsigned(679, 10), 166 => to_unsigned(995, 10), 167 => to_unsigned(369, 10), 168 => to_unsigned(115, 10), 169 => to_unsigned(299, 10), 170 => to_unsigned(442, 10), 171 => to_unsigned(1003, 10), 172 => to_unsigned(646, 10), 173 => to_unsigned(106, 10), 174 => to_unsigned(518, 10), 175 => to_unsigned(947, 10), 176 => to_unsigned(476, 10), 177 => to_unsigned(41, 10), 178 => to_unsigned(717, 10), 179 => to_unsigned(740, 10), 180 => to_unsigned(678, 10), 181 => to_unsigned(753, 10), 182 => to_unsigned(660, 10), 183 => to_unsigned(113, 10), 184 => to_unsigned(795, 10), 185 => to_unsigned(981, 10), 186 => to_unsigned(99, 10), 187 => to_unsigned(782, 10), 188 => to_unsigned(994, 10), 189 => to_unsigned(882, 10), 190 => to_unsigned(1010, 10), 191 => to_unsigned(1000, 10), 192 => to_unsigned(400, 10), 193 => to_unsigned(316, 10), 194 => to_unsigned(782, 10), 195 => to_unsigned(161, 10), 196 => to_unsigned(821, 10), 197 => to_unsigned(404, 10), 198 => to_unsigned(1006, 10), 199 => to_unsigned(336, 10), 200 => to_unsigned(54, 10), 201 => to_unsigned(94, 10), 202 => to_unsigned(810, 10), 203 => to_unsigned(142, 10), 204 => to_unsigned(882, 10), 205 => to_unsigned(917, 10), 206 => to_unsigned(775, 10), 207 => to_unsigned(185, 10), 208 => to_unsigned(818, 10), 209 => to_unsigned(185, 10), 210 => to_unsigned(673, 10), 211 => to_unsigned(777, 10), 212 => to_unsigned(257, 10), 213 => to_unsigned(968, 10), 214 => to_unsigned(389, 10), 215 => to_unsigned(110, 10), 216 => to_unsigned(556, 10), 217 => to_unsigned(667, 10), 218 => to_unsigned(150, 10), 219 => to_unsigned(771, 10), 220 => to_unsigned(827, 10), 221 => to_unsigned(760, 10), 222 => to_unsigned(979, 10), 223 => to_unsigned(175, 10), 224 => to_unsigned(824, 10), 225 => to_unsigned(459, 10), 226 => to_unsigned(51, 10), 227 => to_unsigned(235, 10), 228 => to_unsigned(68, 10), 229 => to_unsigned(306, 10), 230 => to_unsigned(648, 10), 231 => to_unsigned(100, 10), 232 => to_unsigned(163, 10), 233 => to_unsigned(565, 10), 234 => to_unsigned(463, 10), 235 => to_unsigned(17, 10), 236 => to_unsigned(886, 10), 237 => to_unsigned(469, 10), 238 => to_unsigned(571, 10), 239 => to_unsigned(322, 10), 240 => to_unsigned(987, 10), 241 => to_unsigned(583, 10), 242 => to_unsigned(410, 10), 243 => to_unsigned(0, 10), 244 => to_unsigned(608, 10), 245 => to_unsigned(264, 10), 246 => to_unsigned(319, 10), 247 => to_unsigned(954, 10), 248 => to_unsigned(71, 10), 249 => to_unsigned(442, 10), 250 => to_unsigned(92, 10), 251 => to_unsigned(879, 10), 252 => to_unsigned(283, 10), 253 => to_unsigned(333, 10), 254 => to_unsigned(404, 10), 255 => to_unsigned(703, 10), 256 => to_unsigned(357, 10), 257 => to_unsigned(145, 10), 258 => to_unsigned(880, 10), 259 => to_unsigned(88, 10), 260 => to_unsigned(980, 10), 261 => to_unsigned(68, 10), 262 => to_unsigned(524, 10), 263 => to_unsigned(11, 10), 264 => to_unsigned(522, 10), 265 => to_unsigned(568, 10), 266 => to_unsigned(845, 10), 267 => to_unsigned(58, 10), 268 => to_unsigned(523, 10), 269 => to_unsigned(672, 10), 270 => to_unsigned(220, 10), 271 => to_unsigned(316, 10), 272 => to_unsigned(971, 10), 273 => to_unsigned(423, 10), 274 => to_unsigned(965, 10), 275 => to_unsigned(241, 10), 276 => to_unsigned(627, 10), 277 => to_unsigned(417, 10), 278 => to_unsigned(740, 10), 279 => to_unsigned(189, 10), 280 => to_unsigned(353, 10), 281 => to_unsigned(161, 10), 282 => to_unsigned(518, 10), 283 => to_unsigned(158, 10), 284 => to_unsigned(486, 10), 285 => to_unsigned(859, 10), 286 => to_unsigned(398, 10), 287 => to_unsigned(97, 10), 288 => to_unsigned(986, 10), 289 => to_unsigned(995, 10), 290 => to_unsigned(855, 10), 291 => to_unsigned(468, 10), 292 => to_unsigned(707, 10), 293 => to_unsigned(982, 10), 294 => to_unsigned(325, 10), 295 => to_unsigned(781, 10), 296 => to_unsigned(159, 10), 297 => to_unsigned(755, 10), 298 => to_unsigned(719, 10), 299 => to_unsigned(325, 10), 300 => to_unsigned(820, 10), 301 => to_unsigned(81, 10), 302 => to_unsigned(870, 10), 303 => to_unsigned(479, 10), 304 => to_unsigned(115, 10), 305 => to_unsigned(344, 10), 306 => to_unsigned(854, 10), 307 => to_unsigned(953, 10), 308 => to_unsigned(785, 10), 309 => to_unsigned(635, 10), 310 => to_unsigned(190, 10), 311 => to_unsigned(836, 10), 312 => to_unsigned(107, 10), 313 => to_unsigned(977, 10), 314 => to_unsigned(173, 10), 315 => to_unsigned(182, 10), 316 => to_unsigned(703, 10), 317 => to_unsigned(489, 10), 318 => to_unsigned(838, 10), 319 => to_unsigned(1004, 10), 320 => to_unsigned(187, 10), 321 => to_unsigned(725, 10), 322 => to_unsigned(390, 10), 323 => to_unsigned(812, 10), 324 => to_unsigned(798, 10), 325 => to_unsigned(564, 10), 326 => to_unsigned(406, 10), 327 => to_unsigned(496, 10), 328 => to_unsigned(790, 10), 329 => to_unsigned(938, 10), 330 => to_unsigned(53, 10), 331 => to_unsigned(305, 10), 332 => to_unsigned(90, 10), 333 => to_unsigned(424, 10), 334 => to_unsigned(1015, 10), 335 => to_unsigned(845, 10), 336 => to_unsigned(776, 10), 337 => to_unsigned(303, 10), 338 => to_unsigned(509, 10), 339 => to_unsigned(908, 10), 340 => to_unsigned(984, 10), 341 => to_unsigned(495, 10), 342 => to_unsigned(1023, 10), 343 => to_unsigned(663, 10), 344 => to_unsigned(626, 10), 345 => to_unsigned(805, 10), 346 => to_unsigned(9, 10), 347 => to_unsigned(289, 10), 348 => to_unsigned(1016, 10), 349 => to_unsigned(604, 10), 350 => to_unsigned(481, 10), 351 => to_unsigned(650, 10), 352 => to_unsigned(898, 10), 353 => to_unsigned(219, 10), 354 => to_unsigned(142, 10), 355 => to_unsigned(858, 10), 356 => to_unsigned(771, 10), 357 => to_unsigned(531, 10), 358 => to_unsigned(447, 10), 359 => to_unsigned(716, 10), 360 => to_unsigned(567, 10), 361 => to_unsigned(218, 10), 362 => to_unsigned(842, 10), 363 => to_unsigned(818, 10), 364 => to_unsigned(920, 10), 365 => to_unsigned(996, 10), 366 => to_unsigned(696, 10), 367 => to_unsigned(883, 10), 368 => to_unsigned(938, 10), 369 => to_unsigned(1022, 10), 370 => to_unsigned(997, 10), 371 => to_unsigned(388, 10), 372 => to_unsigned(515, 10), 373 => to_unsigned(964, 10), 374 => to_unsigned(521, 10), 375 => to_unsigned(105, 10), 376 => to_unsigned(975, 10), 377 => to_unsigned(163, 10), 378 => to_unsigned(618, 10), 379 => to_unsigned(380, 10), 380 => to_unsigned(643, 10), 381 => to_unsigned(966, 10), 382 => to_unsigned(78, 10), 383 => to_unsigned(792, 10), 384 => to_unsigned(325, 10), 385 => to_unsigned(808, 10), 386 => to_unsigned(584, 10), 387 => to_unsigned(680, 10), 388 => to_unsigned(142, 10), 389 => to_unsigned(776, 10), 390 => to_unsigned(744, 10), 391 => to_unsigned(624, 10), 392 => to_unsigned(35, 10), 393 => to_unsigned(149, 10), 394 => to_unsigned(643, 10), 395 => to_unsigned(678, 10), 396 => to_unsigned(214, 10), 397 => to_unsigned(197, 10), 398 => to_unsigned(125, 10), 399 => to_unsigned(512, 10), 400 => to_unsigned(48, 10), 401 => to_unsigned(149, 10), 402 => to_unsigned(559, 10), 403 => to_unsigned(608, 10), 404 => to_unsigned(816, 10), 405 => to_unsigned(952, 10), 406 => to_unsigned(903, 10), 407 => to_unsigned(407, 10), 408 => to_unsigned(388, 10), 409 => to_unsigned(542, 10), 410 => to_unsigned(369, 10), 411 => to_unsigned(397, 10), 412 => to_unsigned(690, 10), 413 => to_unsigned(753, 10), 414 => to_unsigned(515, 10), 415 => to_unsigned(954, 10), 416 => to_unsigned(196, 10), 417 => to_unsigned(682, 10), 418 => to_unsigned(665, 10), 419 => to_unsigned(850, 10), 420 => to_unsigned(28, 10), 421 => to_unsigned(848, 10), 422 => to_unsigned(49, 10), 423 => to_unsigned(945, 10), 424 => to_unsigned(398, 10), 425 => to_unsigned(619, 10), 426 => to_unsigned(868, 10), 427 => to_unsigned(714, 10), 428 => to_unsigned(871, 10), 429 => to_unsigned(353, 10), 430 => to_unsigned(574, 10), 431 => to_unsigned(89, 10), 432 => to_unsigned(438, 10), 433 => to_unsigned(757, 10), 434 => to_unsigned(987, 10), 435 => to_unsigned(628, 10), 436 => to_unsigned(335, 10), 437 => to_unsigned(939, 10), 438 => to_unsigned(753, 10), 439 => to_unsigned(626, 10), 440 => to_unsigned(248, 10), 441 => to_unsigned(427, 10), 442 => to_unsigned(809, 10), 443 => to_unsigned(414, 10), 444 => to_unsigned(698, 10), 445 => to_unsigned(725, 10), 446 => to_unsigned(325, 10), 447 => to_unsigned(404, 10), 448 => to_unsigned(925, 10), 449 => to_unsigned(993, 10), 450 => to_unsigned(825, 10), 451 => to_unsigned(255, 10), 452 => to_unsigned(562, 10), 453 => to_unsigned(460, 10), 454 => to_unsigned(844, 10), 455 => to_unsigned(102, 10), 456 => to_unsigned(537, 10), 457 => to_unsigned(518, 10), 458 => to_unsigned(162, 10), 459 => to_unsigned(805, 10), 460 => to_unsigned(938, 10), 461 => to_unsigned(753, 10), 462 => to_unsigned(614, 10), 463 => to_unsigned(816, 10), 464 => to_unsigned(438, 10), 465 => to_unsigned(946, 10), 466 => to_unsigned(95, 10), 467 => to_unsigned(710, 10), 468 => to_unsigned(365, 10), 469 => to_unsigned(776, 10), 470 => to_unsigned(955, 10), 471 => to_unsigned(125, 10), 472 => to_unsigned(670, 10), 473 => to_unsigned(678, 10), 474 => to_unsigned(990, 10), 475 => to_unsigned(889, 10), 476 => to_unsigned(925, 10), 477 => to_unsigned(350, 10), 478 => to_unsigned(514, 10), 479 => to_unsigned(126, 10), 480 => to_unsigned(634, 10), 481 => to_unsigned(212, 10), 482 => to_unsigned(441, 10), 483 => to_unsigned(82, 10), 484 => to_unsigned(756, 10), 485 => to_unsigned(311, 10), 486 => to_unsigned(472, 10), 487 => to_unsigned(731, 10), 488 => to_unsigned(544, 10), 489 => to_unsigned(852, 10), 490 => to_unsigned(165, 10), 491 => to_unsigned(501, 10), 492 => to_unsigned(577, 10), 493 => to_unsigned(766, 10), 494 => to_unsigned(166, 10), 495 => to_unsigned(461, 10), 496 => to_unsigned(13, 10), 497 => to_unsigned(470, 10), 498 => to_unsigned(887, 10), 499 => to_unsigned(837, 10), 500 => to_unsigned(481, 10), 501 => to_unsigned(899, 10), 502 => to_unsigned(681, 10), 503 => to_unsigned(773, 10), 504 => to_unsigned(414, 10), 505 => to_unsigned(388, 10), 506 => to_unsigned(759, 10), 507 => to_unsigned(1004, 10), 508 => to_unsigned(1008, 10), 509 => to_unsigned(868, 10), 510 => to_unsigned(890, 10), 511 => to_unsigned(51, 10), 512 => to_unsigned(614, 10), 513 => to_unsigned(897, 10), 514 => to_unsigned(779, 10), 515 => to_unsigned(946, 10), 516 => to_unsigned(632, 10), 517 => to_unsigned(339, 10), 518 => to_unsigned(468, 10), 519 => to_unsigned(847, 10), 520 => to_unsigned(64, 10), 521 => to_unsigned(1023, 10), 522 => to_unsigned(237, 10), 523 => to_unsigned(437, 10), 524 => to_unsigned(294, 10), 525 => to_unsigned(344, 10), 526 => to_unsigned(921, 10), 527 => to_unsigned(106, 10), 528 => to_unsigned(115, 10), 529 => to_unsigned(974, 10), 530 => to_unsigned(656, 10), 531 => to_unsigned(866, 10), 532 => to_unsigned(925, 10), 533 => to_unsigned(693, 10), 534 => to_unsigned(1009, 10), 535 => to_unsigned(344, 10), 536 => to_unsigned(184, 10), 537 => to_unsigned(921, 10), 538 => to_unsigned(254, 10), 539 => to_unsigned(270, 10), 540 => to_unsigned(92, 10), 541 => to_unsigned(83, 10), 542 => to_unsigned(959, 10), 543 => to_unsigned(136, 10), 544 => to_unsigned(126, 10), 545 => to_unsigned(83, 10), 546 => to_unsigned(764, 10), 547 => to_unsigned(160, 10), 548 => to_unsigned(150, 10), 549 => to_unsigned(272, 10), 550 => to_unsigned(41, 10), 551 => to_unsigned(159, 10), 552 => to_unsigned(708, 10), 553 => to_unsigned(20, 10), 554 => to_unsigned(622, 10), 555 => to_unsigned(77, 10), 556 => to_unsigned(62, 10), 557 => to_unsigned(272, 10), 558 => to_unsigned(973, 10), 559 => to_unsigned(218, 10), 560 => to_unsigned(1016, 10), 561 => to_unsigned(544, 10), 562 => to_unsigned(198, 10), 563 => to_unsigned(381, 10), 564 => to_unsigned(229, 10), 565 => to_unsigned(728, 10), 566 => to_unsigned(777, 10), 567 => to_unsigned(1012, 10), 568 => to_unsigned(469, 10), 569 => to_unsigned(276, 10), 570 => to_unsigned(668, 10), 571 => to_unsigned(847, 10), 572 => to_unsigned(15, 10), 573 => to_unsigned(364, 10), 574 => to_unsigned(524, 10), 575 => to_unsigned(351, 10), 576 => to_unsigned(44, 10), 577 => to_unsigned(814, 10), 578 => to_unsigned(119, 10), 579 => to_unsigned(823, 10), 580 => to_unsigned(589, 10), 581 => to_unsigned(338, 10), 582 => to_unsigned(473, 10), 583 => to_unsigned(900, 10), 584 => to_unsigned(325, 10), 585 => to_unsigned(414, 10), 586 => to_unsigned(264, 10), 587 => to_unsigned(742, 10), 588 => to_unsigned(642, 10), 589 => to_unsigned(929, 10), 590 => to_unsigned(290, 10), 591 => to_unsigned(847, 10), 592 => to_unsigned(546, 10), 593 => to_unsigned(864, 10), 594 => to_unsigned(515, 10), 595 => to_unsigned(570, 10), 596 => to_unsigned(948, 10), 597 => to_unsigned(234, 10), 598 => to_unsigned(57, 10), 599 => to_unsigned(763, 10), 600 => to_unsigned(451, 10), 601 => to_unsigned(853, 10), 602 => to_unsigned(823, 10), 603 => to_unsigned(804, 10), 604 => to_unsigned(957, 10), 605 => to_unsigned(186, 10), 606 => to_unsigned(582, 10), 607 => to_unsigned(85, 10), 608 => to_unsigned(377, 10), 609 => to_unsigned(782, 10), 610 => to_unsigned(373, 10), 611 => to_unsigned(14, 10), 612 => to_unsigned(721, 10), 613 => to_unsigned(350, 10), 614 => to_unsigned(59, 10), 615 => to_unsigned(467, 10), 616 => to_unsigned(876, 10), 617 => to_unsigned(493, 10), 618 => to_unsigned(610, 10), 619 => to_unsigned(352, 10), 620 => to_unsigned(608, 10), 621 => to_unsigned(477, 10), 622 => to_unsigned(54, 10), 623 => to_unsigned(23, 10), 624 => to_unsigned(326, 10), 625 => to_unsigned(362, 10), 626 => to_unsigned(55, 10), 627 => to_unsigned(991, 10), 628 => to_unsigned(48, 10), 629 => to_unsigned(662, 10), 630 => to_unsigned(86, 10), 631 => to_unsigned(950, 10), 632 => to_unsigned(1003, 10), 633 => to_unsigned(352, 10), 634 => to_unsigned(897, 10), 635 => to_unsigned(509, 10), 636 => to_unsigned(852, 10), 637 => to_unsigned(660, 10), 638 => to_unsigned(653, 10), 639 => to_unsigned(318, 10), 640 => to_unsigned(966, 10), 641 => to_unsigned(357, 10), 642 => to_unsigned(574, 10), 643 => to_unsigned(176, 10), 644 => to_unsigned(802, 10), 645 => to_unsigned(229, 10), 646 => to_unsigned(486, 10), 647 => to_unsigned(980, 10), 648 => to_unsigned(1005, 10), 649 => to_unsigned(546, 10), 650 => to_unsigned(307, 10), 651 => to_unsigned(138, 10), 652 => to_unsigned(597, 10), 653 => to_unsigned(350, 10), 654 => to_unsigned(170, 10), 655 => to_unsigned(897, 10), 656 => to_unsigned(518, 10), 657 => to_unsigned(156, 10), 658 => to_unsigned(844, 10), 659 => to_unsigned(944, 10), 660 => to_unsigned(315, 10), 661 => to_unsigned(434, 10), 662 => to_unsigned(191, 10), 663 => to_unsigned(331, 10), 664 => to_unsigned(746, 10), 665 => to_unsigned(692, 10), 666 => to_unsigned(373, 10), 667 => to_unsigned(76, 10), 668 => to_unsigned(751, 10), 669 => to_unsigned(48, 10), 670 => to_unsigned(389, 10), 671 => to_unsigned(302, 10), 672 => to_unsigned(759, 10), 673 => to_unsigned(852, 10), 674 => to_unsigned(527, 10), 675 => to_unsigned(16, 10), 676 => to_unsigned(883, 10), 677 => to_unsigned(492, 10), 678 => to_unsigned(320, 10), 679 => to_unsigned(409, 10), 680 => to_unsigned(359, 10), 681 => to_unsigned(356, 10), 682 => to_unsigned(360, 10), 683 => to_unsigned(191, 10), 684 => to_unsigned(37, 10), 685 => to_unsigned(879, 10), 686 => to_unsigned(797, 10), 687 => to_unsigned(425, 10), 688 => to_unsigned(331, 10), 689 => to_unsigned(937, 10), 690 => to_unsigned(90, 10), 691 => to_unsigned(646, 10), 692 => to_unsigned(726, 10), 693 => to_unsigned(488, 10), 694 => to_unsigned(225, 10), 695 => to_unsigned(364, 10), 696 => to_unsigned(285, 10), 697 => to_unsigned(850, 10), 698 => to_unsigned(986, 10), 699 => to_unsigned(587, 10), 700 => to_unsigned(1013, 10), 701 => to_unsigned(433, 10), 702 => to_unsigned(981, 10), 703 => to_unsigned(136, 10), 704 => to_unsigned(362, 10), 705 => to_unsigned(429, 10), 706 => to_unsigned(1001, 10), 707 => to_unsigned(944, 10), 708 => to_unsigned(160, 10), 709 => to_unsigned(410, 10), 710 => to_unsigned(271, 10), 711 => to_unsigned(690, 10), 712 => to_unsigned(208, 10), 713 => to_unsigned(640, 10), 714 => to_unsigned(585, 10), 715 => to_unsigned(616, 10), 716 => to_unsigned(903, 10), 717 => to_unsigned(221, 10), 718 => to_unsigned(483, 10), 719 => to_unsigned(384, 10), 720 => to_unsigned(1008, 10), 721 => to_unsigned(928, 10), 722 => to_unsigned(992, 10), 723 => to_unsigned(398, 10), 724 => to_unsigned(562, 10), 725 => to_unsigned(71, 10), 726 => to_unsigned(610, 10), 727 => to_unsigned(280, 10), 728 => to_unsigned(802, 10), 729 => to_unsigned(656, 10), 730 => to_unsigned(778, 10), 731 => to_unsigned(566, 10), 732 => to_unsigned(754, 10), 733 => to_unsigned(9, 10), 734 => to_unsigned(395, 10), 735 => to_unsigned(1004, 10), 736 => to_unsigned(660, 10), 737 => to_unsigned(446, 10), 738 => to_unsigned(531, 10), 739 => to_unsigned(429, 10), 740 => to_unsigned(340, 10), 741 => to_unsigned(992, 10), 742 => to_unsigned(242, 10), 743 => to_unsigned(278, 10), 744 => to_unsigned(983, 10), 745 => to_unsigned(241, 10), 746 => to_unsigned(861, 10), 747 => to_unsigned(855, 10), 748 => to_unsigned(63, 10), 749 => to_unsigned(944, 10), 750 => to_unsigned(454, 10), 751 => to_unsigned(629, 10), 752 => to_unsigned(434, 10), 753 => to_unsigned(183, 10), 754 => to_unsigned(325, 10), 755 => to_unsigned(654, 10), 756 => to_unsigned(75, 10), 757 => to_unsigned(26, 10), 758 => to_unsigned(716, 10), 759 => to_unsigned(806, 10), 760 => to_unsigned(931, 10), 761 => to_unsigned(813, 10), 762 => to_unsigned(933, 10), 763 => to_unsigned(33, 10), 764 => to_unsigned(923, 10), 765 => to_unsigned(299, 10), 766 => to_unsigned(318, 10), 767 => to_unsigned(344, 10), 768 => to_unsigned(555, 10), 769 => to_unsigned(804, 10), 770 => to_unsigned(104, 10), 771 => to_unsigned(557, 10), 772 => to_unsigned(672, 10), 773 => to_unsigned(130, 10), 774 => to_unsigned(258, 10), 775 => to_unsigned(204, 10), 776 => to_unsigned(791, 10), 777 => to_unsigned(597, 10), 778 => to_unsigned(496, 10), 779 => to_unsigned(903, 10), 780 => to_unsigned(610, 10), 781 => to_unsigned(479, 10), 782 => to_unsigned(323, 10), 783 => to_unsigned(954, 10), 784 => to_unsigned(454, 10), 785 => to_unsigned(924, 10), 786 => to_unsigned(296, 10), 787 => to_unsigned(466, 10), 788 => to_unsigned(944, 10), 789 => to_unsigned(564, 10), 790 => to_unsigned(716, 10), 791 => to_unsigned(193, 10), 792 => to_unsigned(141, 10), 793 => to_unsigned(456, 10), 794 => to_unsigned(30, 10), 795 => to_unsigned(719, 10), 796 => to_unsigned(56, 10), 797 => to_unsigned(49, 10), 798 => to_unsigned(997, 10), 799 => to_unsigned(860, 10), 800 => to_unsigned(229, 10), 801 => to_unsigned(608, 10), 802 => to_unsigned(795, 10), 803 => to_unsigned(733, 10), 804 => to_unsigned(857, 10), 805 => to_unsigned(676, 10), 806 => to_unsigned(139, 10), 807 => to_unsigned(82, 10), 808 => to_unsigned(825, 10), 809 => to_unsigned(716, 10), 810 => to_unsigned(213, 10), 811 => to_unsigned(838, 10), 812 => to_unsigned(969, 10), 813 => to_unsigned(485, 10), 814 => to_unsigned(421, 10), 815 => to_unsigned(555, 10), 816 => to_unsigned(256, 10), 817 => to_unsigned(105, 10), 818 => to_unsigned(965, 10), 819 => to_unsigned(346, 10), 820 => to_unsigned(36, 10), 821 => to_unsigned(397, 10), 822 => to_unsigned(14, 10), 823 => to_unsigned(563, 10), 824 => to_unsigned(551, 10), 825 => to_unsigned(572, 10), 826 => to_unsigned(658, 10), 827 => to_unsigned(507, 10), 828 => to_unsigned(377, 10), 829 => to_unsigned(936, 10), 830 => to_unsigned(389, 10), 831 => to_unsigned(766, 10), 832 => to_unsigned(214, 10), 833 => to_unsigned(630, 10), 834 => to_unsigned(776, 10), 835 => to_unsigned(760, 10), 836 => to_unsigned(227, 10), 837 => to_unsigned(782, 10), 838 => to_unsigned(363, 10), 839 => to_unsigned(691, 10), 840 => to_unsigned(969, 10), 841 => to_unsigned(365, 10), 842 => to_unsigned(105, 10), 843 => to_unsigned(956, 10), 844 => to_unsigned(656, 10), 845 => to_unsigned(618, 10), 846 => to_unsigned(786, 10), 847 => to_unsigned(302, 10), 848 => to_unsigned(292, 10), 849 => to_unsigned(349, 10), 850 => to_unsigned(1010, 10), 851 => to_unsigned(449, 10), 852 => to_unsigned(999, 10), 853 => to_unsigned(469, 10), 854 => to_unsigned(762, 10), 855 => to_unsigned(817, 10), 856 => to_unsigned(291, 10), 857 => to_unsigned(343, 10), 858 => to_unsigned(708, 10), 859 => to_unsigned(509, 10), 860 => to_unsigned(833, 10), 861 => to_unsigned(758, 10), 862 => to_unsigned(533, 10), 863 => to_unsigned(947, 10), 864 => to_unsigned(287, 10), 865 => to_unsigned(355, 10), 866 => to_unsigned(134, 10), 867 => to_unsigned(514, 10), 868 => to_unsigned(655, 10), 869 => to_unsigned(699, 10), 870 => to_unsigned(1013, 10), 871 => to_unsigned(698, 10), 872 => to_unsigned(250, 10), 873 => to_unsigned(551, 10), 874 => to_unsigned(916, 10), 875 => to_unsigned(288, 10), 876 => to_unsigned(216, 10), 877 => to_unsigned(930, 10), 878 => to_unsigned(710, 10), 879 => to_unsigned(827, 10), 880 => to_unsigned(438, 10), 881 => to_unsigned(756, 10), 882 => to_unsigned(744, 10), 883 => to_unsigned(137, 10), 884 => to_unsigned(43, 10), 885 => to_unsigned(525, 10), 886 => to_unsigned(201, 10), 887 => to_unsigned(120, 10), 888 => to_unsigned(852, 10), 889 => to_unsigned(845, 10), 890 => to_unsigned(758, 10), 891 => to_unsigned(141, 10), 892 => to_unsigned(500, 10), 893 => to_unsigned(716, 10), 894 => to_unsigned(469, 10), 895 => to_unsigned(634, 10), 896 => to_unsigned(293, 10), 897 => to_unsigned(204, 10), 898 => to_unsigned(78, 10), 899 => to_unsigned(457, 10), 900 => to_unsigned(871, 10), 901 => to_unsigned(283, 10), 902 => to_unsigned(485, 10), 903 => to_unsigned(990, 10), 904 => to_unsigned(787, 10), 905 => to_unsigned(356, 10), 906 => to_unsigned(277, 10), 907 => to_unsigned(6, 10), 908 => to_unsigned(611, 10), 909 => to_unsigned(834, 10), 910 => to_unsigned(757, 10), 911 => to_unsigned(294, 10), 912 => to_unsigned(531, 10), 913 => to_unsigned(772, 10), 914 => to_unsigned(720, 10), 915 => to_unsigned(209, 10), 916 => to_unsigned(678, 10), 917 => to_unsigned(589, 10), 918 => to_unsigned(382, 10), 919 => to_unsigned(747, 10), 920 => to_unsigned(942, 10), 921 => to_unsigned(677, 10), 922 => to_unsigned(281, 10), 923 => to_unsigned(525, 10), 924 => to_unsigned(981, 10), 925 => to_unsigned(444, 10), 926 => to_unsigned(293, 10), 927 => to_unsigned(298, 10), 928 => to_unsigned(361, 10), 929 => to_unsigned(744, 10), 930 => to_unsigned(260, 10), 931 => to_unsigned(602, 10), 932 => to_unsigned(953, 10), 933 => to_unsigned(982, 10), 934 => to_unsigned(334, 10), 935 => to_unsigned(241, 10), 936 => to_unsigned(846, 10), 937 => to_unsigned(42, 10), 938 => to_unsigned(723, 10), 939 => to_unsigned(921, 10), 940 => to_unsigned(862, 10), 941 => to_unsigned(176, 10), 942 => to_unsigned(36, 10), 943 => to_unsigned(907, 10), 944 => to_unsigned(950, 10), 945 => to_unsigned(734, 10), 946 => to_unsigned(570, 10), 947 => to_unsigned(534, 10), 948 => to_unsigned(577, 10), 949 => to_unsigned(875, 10), 950 => to_unsigned(628, 10), 951 => to_unsigned(410, 10), 952 => to_unsigned(976, 10), 953 => to_unsigned(656, 10), 954 => to_unsigned(736, 10), 955 => to_unsigned(208, 10), 956 => to_unsigned(837, 10), 957 => to_unsigned(138, 10), 958 => to_unsigned(971, 10), 959 => to_unsigned(533, 10), 960 => to_unsigned(228, 10), 961 => to_unsigned(419, 10), 962 => to_unsigned(752, 10), 963 => to_unsigned(60, 10), 964 => to_unsigned(726, 10), 965 => to_unsigned(480, 10), 966 => to_unsigned(441, 10), 967 => to_unsigned(480, 10), 968 => to_unsigned(529, 10), 969 => to_unsigned(77, 10), 970 => to_unsigned(403, 10), 971 => to_unsigned(853, 10), 972 => to_unsigned(759, 10), 973 => to_unsigned(746, 10), 974 => to_unsigned(580, 10), 975 => to_unsigned(600, 10), 976 => to_unsigned(343, 10), 977 => to_unsigned(897, 10), 978 => to_unsigned(903, 10), 979 => to_unsigned(554, 10), 980 => to_unsigned(74, 10), 981 => to_unsigned(769, 10), 982 => to_unsigned(790, 10), 983 => to_unsigned(306, 10), 984 => to_unsigned(967, 10), 985 => to_unsigned(649, 10), 986 => to_unsigned(220, 10), 987 => to_unsigned(763, 10), 988 => to_unsigned(812, 10), 989 => to_unsigned(891, 10), 990 => to_unsigned(233, 10), 991 => to_unsigned(814, 10), 992 => to_unsigned(915, 10), 993 => to_unsigned(250, 10), 994 => to_unsigned(103, 10), 995 => to_unsigned(453, 10), 996 => to_unsigned(90, 10), 997 => to_unsigned(264, 10), 998 => to_unsigned(569, 10), 999 => to_unsigned(44, 10), 1000 => to_unsigned(85, 10), 1001 => to_unsigned(145, 10), 1002 => to_unsigned(645, 10), 1003 => to_unsigned(974, 10), 1004 => to_unsigned(352, 10), 1005 => to_unsigned(293, 10), 1006 => to_unsigned(667, 10), 1007 => to_unsigned(990, 10), 1008 => to_unsigned(61, 10), 1009 => to_unsigned(828, 10), 1010 => to_unsigned(188, 10), 1011 => to_unsigned(442, 10), 1012 => to_unsigned(184, 10), 1013 => to_unsigned(966, 10), 1014 => to_unsigned(204, 10), 1015 => to_unsigned(587, 10), 1016 => to_unsigned(155, 10), 1017 => to_unsigned(628, 10), 1018 => to_unsigned(209, 10), 1019 => to_unsigned(722, 10), 1020 => to_unsigned(207, 10), 1021 => to_unsigned(772, 10), 1022 => to_unsigned(528, 10), 1023 => to_unsigned(891, 10), 1024 => to_unsigned(359, 10), 1025 => to_unsigned(584, 10), 1026 => to_unsigned(139, 10), 1027 => to_unsigned(937, 10), 1028 => to_unsigned(42, 10), 1029 => to_unsigned(958, 10), 1030 => to_unsigned(780, 10), 1031 => to_unsigned(125, 10), 1032 => to_unsigned(804, 10), 1033 => to_unsigned(534, 10), 1034 => to_unsigned(890, 10), 1035 => to_unsigned(981, 10), 1036 => to_unsigned(124, 10), 1037 => to_unsigned(683, 10), 1038 => to_unsigned(636, 10), 1039 => to_unsigned(318, 10), 1040 => to_unsigned(639, 10), 1041 => to_unsigned(329, 10), 1042 => to_unsigned(376, 10), 1043 => to_unsigned(123, 10), 1044 => to_unsigned(844, 10), 1045 => to_unsigned(977, 10), 1046 => to_unsigned(215, 10), 1047 => to_unsigned(692, 10), 1048 => to_unsigned(55, 10), 1049 => to_unsigned(143, 10), 1050 => to_unsigned(387, 10), 1051 => to_unsigned(351, 10), 1052 => to_unsigned(58, 10), 1053 => to_unsigned(253, 10), 1054 => to_unsigned(303, 10), 1055 => to_unsigned(189, 10), 1056 => to_unsigned(139, 10), 1057 => to_unsigned(416, 10), 1058 => to_unsigned(618, 10), 1059 => to_unsigned(463, 10), 1060 => to_unsigned(921, 10), 1061 => to_unsigned(143, 10), 1062 => to_unsigned(833, 10), 1063 => to_unsigned(605, 10), 1064 => to_unsigned(528, 10), 1065 => to_unsigned(29, 10), 1066 => to_unsigned(312, 10), 1067 => to_unsigned(356, 10), 1068 => to_unsigned(605, 10), 1069 => to_unsigned(448, 10), 1070 => to_unsigned(573, 10), 1071 => to_unsigned(759, 10), 1072 => to_unsigned(295, 10), 1073 => to_unsigned(854, 10), 1074 => to_unsigned(258, 10), 1075 => to_unsigned(357, 10), 1076 => to_unsigned(688, 10), 1077 => to_unsigned(254, 10), 1078 => to_unsigned(787, 10), 1079 => to_unsigned(711, 10), 1080 => to_unsigned(910, 10), 1081 => to_unsigned(482, 10), 1082 => to_unsigned(926, 10), 1083 => to_unsigned(387, 10), 1084 => to_unsigned(586, 10), 1085 => to_unsigned(632, 10), 1086 => to_unsigned(236, 10), 1087 => to_unsigned(534, 10), 1088 => to_unsigned(815, 10), 1089 => to_unsigned(746, 10), 1090 => to_unsigned(822, 10), 1091 => to_unsigned(238, 10), 1092 => to_unsigned(983, 10), 1093 => to_unsigned(944, 10), 1094 => to_unsigned(127, 10), 1095 => to_unsigned(73, 10), 1096 => to_unsigned(545, 10), 1097 => to_unsigned(881, 10), 1098 => to_unsigned(218, 10), 1099 => to_unsigned(136, 10), 1100 => to_unsigned(157, 10), 1101 => to_unsigned(348, 10), 1102 => to_unsigned(993, 10), 1103 => to_unsigned(177, 10), 1104 => to_unsigned(360, 10), 1105 => to_unsigned(245, 10), 1106 => to_unsigned(182, 10), 1107 => to_unsigned(940, 10), 1108 => to_unsigned(892, 10), 1109 => to_unsigned(146, 10), 1110 => to_unsigned(462, 10), 1111 => to_unsigned(770, 10), 1112 => to_unsigned(1000, 10), 1113 => to_unsigned(650, 10), 1114 => to_unsigned(217, 10), 1115 => to_unsigned(326, 10), 1116 => to_unsigned(156, 10), 1117 => to_unsigned(53, 10), 1118 => to_unsigned(476, 10), 1119 => to_unsigned(400, 10), 1120 => to_unsigned(743, 10), 1121 => to_unsigned(85, 10), 1122 => to_unsigned(86, 10), 1123 => to_unsigned(61, 10), 1124 => to_unsigned(504, 10), 1125 => to_unsigned(722, 10), 1126 => to_unsigned(128, 10), 1127 => to_unsigned(968, 10), 1128 => to_unsigned(369, 10), 1129 => to_unsigned(322, 10), 1130 => to_unsigned(699, 10), 1131 => to_unsigned(1014, 10), 1132 => to_unsigned(9, 10), 1133 => to_unsigned(291, 10), 1134 => to_unsigned(845, 10), 1135 => to_unsigned(362, 10), 1136 => to_unsigned(442, 10), 1137 => to_unsigned(604, 10), 1138 => to_unsigned(428, 10), 1139 => to_unsigned(917, 10), 1140 => to_unsigned(0, 10), 1141 => to_unsigned(723, 10), 1142 => to_unsigned(456, 10), 1143 => to_unsigned(290, 10), 1144 => to_unsigned(954, 10), 1145 => to_unsigned(88, 10), 1146 => to_unsigned(819, 10), 1147 => to_unsigned(330, 10), 1148 => to_unsigned(500, 10), 1149 => to_unsigned(109, 10), 1150 => to_unsigned(908, 10), 1151 => to_unsigned(773, 10), 1152 => to_unsigned(996, 10), 1153 => to_unsigned(681, 10), 1154 => to_unsigned(884, 10), 1155 => to_unsigned(584, 10), 1156 => to_unsigned(194, 10), 1157 => to_unsigned(631, 10), 1158 => to_unsigned(242, 10), 1159 => to_unsigned(728, 10), 1160 => to_unsigned(745, 10), 1161 => to_unsigned(874, 10), 1162 => to_unsigned(666, 10), 1163 => to_unsigned(594, 10), 1164 => to_unsigned(37, 10), 1165 => to_unsigned(42, 10), 1166 => to_unsigned(766, 10), 1167 => to_unsigned(207, 10), 1168 => to_unsigned(145, 10), 1169 => to_unsigned(360, 10), 1170 => to_unsigned(143, 10), 1171 => to_unsigned(241, 10), 1172 => to_unsigned(1008, 10), 1173 => to_unsigned(128, 10), 1174 => to_unsigned(617, 10), 1175 => to_unsigned(992, 10), 1176 => to_unsigned(366, 10), 1177 => to_unsigned(887, 10), 1178 => to_unsigned(726, 10), 1179 => to_unsigned(675, 10), 1180 => to_unsigned(398, 10), 1181 => to_unsigned(125, 10), 1182 => to_unsigned(544, 10), 1183 => to_unsigned(288, 10), 1184 => to_unsigned(717, 10), 1185 => to_unsigned(314, 10), 1186 => to_unsigned(149, 10), 1187 => to_unsigned(150, 10), 1188 => to_unsigned(522, 10), 1189 => to_unsigned(533, 10), 1190 => to_unsigned(375, 10), 1191 => to_unsigned(979, 10), 1192 => to_unsigned(641, 10), 1193 => to_unsigned(937, 10), 1194 => to_unsigned(739, 10), 1195 => to_unsigned(976, 10), 1196 => to_unsigned(456, 10), 1197 => to_unsigned(3, 10), 1198 => to_unsigned(118, 10), 1199 => to_unsigned(725, 10), 1200 => to_unsigned(271, 10), 1201 => to_unsigned(24, 10), 1202 => to_unsigned(413, 10), 1203 => to_unsigned(983, 10), 1204 => to_unsigned(448, 10), 1205 => to_unsigned(748, 10), 1206 => to_unsigned(896, 10), 1207 => to_unsigned(951, 10), 1208 => to_unsigned(191, 10), 1209 => to_unsigned(33, 10), 1210 => to_unsigned(647, 10), 1211 => to_unsigned(155, 10), 1212 => to_unsigned(470, 10), 1213 => to_unsigned(90, 10), 1214 => to_unsigned(725, 10), 1215 => to_unsigned(484, 10), 1216 => to_unsigned(820, 10), 1217 => to_unsigned(565, 10), 1218 => to_unsigned(51, 10), 1219 => to_unsigned(89, 10), 1220 => to_unsigned(219, 10), 1221 => to_unsigned(777, 10), 1222 => to_unsigned(569, 10), 1223 => to_unsigned(182, 10), 1224 => to_unsigned(688, 10), 1225 => to_unsigned(413, 10), 1226 => to_unsigned(346, 10), 1227 => to_unsigned(393, 10), 1228 => to_unsigned(688, 10), 1229 => to_unsigned(925, 10), 1230 => to_unsigned(884, 10), 1231 => to_unsigned(683, 10), 1232 => to_unsigned(906, 10), 1233 => to_unsigned(1023, 10), 1234 => to_unsigned(422, 10), 1235 => to_unsigned(1001, 10), 1236 => to_unsigned(698, 10), 1237 => to_unsigned(406, 10), 1238 => to_unsigned(272, 10), 1239 => to_unsigned(980, 10), 1240 => to_unsigned(101, 10), 1241 => to_unsigned(684, 10), 1242 => to_unsigned(411, 10), 1243 => to_unsigned(266, 10), 1244 => to_unsigned(365, 10), 1245 => to_unsigned(167, 10), 1246 => to_unsigned(45, 10), 1247 => to_unsigned(428, 10), 1248 => to_unsigned(937, 10), 1249 => to_unsigned(605, 10), 1250 => to_unsigned(635, 10), 1251 => to_unsigned(1021, 10), 1252 => to_unsigned(133, 10), 1253 => to_unsigned(642, 10), 1254 => to_unsigned(304, 10), 1255 => to_unsigned(530, 10), 1256 => to_unsigned(996, 10), 1257 => to_unsigned(102, 10), 1258 => to_unsigned(607, 10), 1259 => to_unsigned(560, 10), 1260 => to_unsigned(823, 10), 1261 => to_unsigned(445, 10), 1262 => to_unsigned(136, 10), 1263 => to_unsigned(470, 10), 1264 => to_unsigned(934, 10), 1265 => to_unsigned(19, 10), 1266 => to_unsigned(762, 10), 1267 => to_unsigned(87, 10), 1268 => to_unsigned(645, 10), 1269 => to_unsigned(702, 10), 1270 => to_unsigned(284, 10), 1271 => to_unsigned(375, 10), 1272 => to_unsigned(801, 10), 1273 => to_unsigned(705, 10), 1274 => to_unsigned(58, 10), 1275 => to_unsigned(67, 10), 1276 => to_unsigned(945, 10), 1277 => to_unsigned(340, 10), 1278 => to_unsigned(718, 10), 1279 => to_unsigned(134, 10), 1280 => to_unsigned(939, 10), 1281 => to_unsigned(757, 10), 1282 => to_unsigned(875, 10), 1283 => to_unsigned(828, 10), 1284 => to_unsigned(667, 10), 1285 => to_unsigned(146, 10), 1286 => to_unsigned(605, 10), 1287 => to_unsigned(177, 10), 1288 => to_unsigned(897, 10), 1289 => to_unsigned(587, 10), 1290 => to_unsigned(477, 10), 1291 => to_unsigned(438, 10), 1292 => to_unsigned(173, 10), 1293 => to_unsigned(767, 10), 1294 => to_unsigned(375, 10), 1295 => to_unsigned(11, 10), 1296 => to_unsigned(924, 10), 1297 => to_unsigned(923, 10), 1298 => to_unsigned(951, 10), 1299 => to_unsigned(534, 10), 1300 => to_unsigned(154, 10), 1301 => to_unsigned(885, 10), 1302 => to_unsigned(675, 10), 1303 => to_unsigned(366, 10), 1304 => to_unsigned(86, 10), 1305 => to_unsigned(472, 10), 1306 => to_unsigned(88, 10), 1307 => to_unsigned(845, 10), 1308 => to_unsigned(486, 10), 1309 => to_unsigned(839, 10), 1310 => to_unsigned(77, 10), 1311 => to_unsigned(782, 10), 1312 => to_unsigned(795, 10), 1313 => to_unsigned(583, 10), 1314 => to_unsigned(341, 10), 1315 => to_unsigned(372, 10), 1316 => to_unsigned(455, 10), 1317 => to_unsigned(152, 10), 1318 => to_unsigned(303, 10), 1319 => to_unsigned(469, 10), 1320 => to_unsigned(122, 10), 1321 => to_unsigned(473, 10), 1322 => to_unsigned(125, 10), 1323 => to_unsigned(115, 10), 1324 => to_unsigned(805, 10), 1325 => to_unsigned(944, 10), 1326 => to_unsigned(969, 10), 1327 => to_unsigned(826, 10), 1328 => to_unsigned(564, 10), 1329 => to_unsigned(391, 10), 1330 => to_unsigned(513, 10), 1331 => to_unsigned(683, 10), 1332 => to_unsigned(889, 10), 1333 => to_unsigned(131, 10), 1334 => to_unsigned(871, 10), 1335 => to_unsigned(31, 10), 1336 => to_unsigned(20, 10), 1337 => to_unsigned(469, 10), 1338 => to_unsigned(528, 10), 1339 => to_unsigned(332, 10), 1340 => to_unsigned(315, 10), 1341 => to_unsigned(405, 10), 1342 => to_unsigned(70, 10), 1343 => to_unsigned(375, 10), 1344 => to_unsigned(521, 10), 1345 => to_unsigned(294, 10), 1346 => to_unsigned(330, 10), 1347 => to_unsigned(816, 10), 1348 => to_unsigned(798, 10), 1349 => to_unsigned(152, 10), 1350 => to_unsigned(169, 10), 1351 => to_unsigned(50, 10), 1352 => to_unsigned(72, 10), 1353 => to_unsigned(495, 10), 1354 => to_unsigned(807, 10), 1355 => to_unsigned(122, 10), 1356 => to_unsigned(193, 10), 1357 => to_unsigned(971, 10), 1358 => to_unsigned(627, 10), 1359 => to_unsigned(444, 10), 1360 => to_unsigned(731, 10), 1361 => to_unsigned(744, 10), 1362 => to_unsigned(37, 10), 1363 => to_unsigned(161, 10), 1364 => to_unsigned(32, 10), 1365 => to_unsigned(333, 10), 1366 => to_unsigned(644, 10), 1367 => to_unsigned(355, 10), 1368 => to_unsigned(817, 10), 1369 => to_unsigned(797, 10), 1370 => to_unsigned(129, 10), 1371 => to_unsigned(190, 10), 1372 => to_unsigned(565, 10), 1373 => to_unsigned(10, 10), 1374 => to_unsigned(198, 10), 1375 => to_unsigned(602, 10), 1376 => to_unsigned(41, 10), 1377 => to_unsigned(507, 10), 1378 => to_unsigned(798, 10), 1379 => to_unsigned(628, 10), 1380 => to_unsigned(716, 10), 1381 => to_unsigned(645, 10), 1382 => to_unsigned(535, 10), 1383 => to_unsigned(1014, 10), 1384 => to_unsigned(224, 10), 1385 => to_unsigned(447, 10), 1386 => to_unsigned(928, 10), 1387 => to_unsigned(581, 10), 1388 => to_unsigned(226, 10), 1389 => to_unsigned(152, 10), 1390 => to_unsigned(793, 10), 1391 => to_unsigned(391, 10), 1392 => to_unsigned(465, 10), 1393 => to_unsigned(984, 10), 1394 => to_unsigned(462, 10), 1395 => to_unsigned(401, 10), 1396 => to_unsigned(820, 10), 1397 => to_unsigned(645, 10), 1398 => to_unsigned(299, 10), 1399 => to_unsigned(929, 10), 1400 => to_unsigned(940, 10), 1401 => to_unsigned(421, 10), 1402 => to_unsigned(660, 10), 1403 => to_unsigned(741, 10), 1404 => to_unsigned(385, 10), 1405 => to_unsigned(524, 10), 1406 => to_unsigned(293, 10), 1407 => to_unsigned(875, 10), 1408 => to_unsigned(208, 10), 1409 => to_unsigned(174, 10), 1410 => to_unsigned(618, 10), 1411 => to_unsigned(228, 10), 1412 => to_unsigned(738, 10), 1413 => to_unsigned(64, 10), 1414 => to_unsigned(419, 10), 1415 => to_unsigned(178, 10), 1416 => to_unsigned(398, 10), 1417 => to_unsigned(601, 10), 1418 => to_unsigned(300, 10), 1419 => to_unsigned(46, 10), 1420 => to_unsigned(645, 10), 1421 => to_unsigned(829, 10), 1422 => to_unsigned(28, 10), 1423 => to_unsigned(716, 10), 1424 => to_unsigned(176, 10), 1425 => to_unsigned(742, 10), 1426 => to_unsigned(455, 10), 1427 => to_unsigned(723, 10), 1428 => to_unsigned(41, 10), 1429 => to_unsigned(469, 10), 1430 => to_unsigned(168, 10), 1431 => to_unsigned(255, 10), 1432 => to_unsigned(25, 10), 1433 => to_unsigned(832, 10), 1434 => to_unsigned(598, 10), 1435 => to_unsigned(299, 10), 1436 => to_unsigned(38, 10), 1437 => to_unsigned(245, 10), 1438 => to_unsigned(537, 10), 1439 => to_unsigned(383, 10), 1440 => to_unsigned(568, 10), 1441 => to_unsigned(428, 10), 1442 => to_unsigned(476, 10), 1443 => to_unsigned(769, 10), 1444 => to_unsigned(194, 10), 1445 => to_unsigned(438, 10), 1446 => to_unsigned(138, 10), 1447 => to_unsigned(749, 10), 1448 => to_unsigned(877, 10), 1449 => to_unsigned(182, 10), 1450 => to_unsigned(299, 10), 1451 => to_unsigned(269, 10), 1452 => to_unsigned(988, 10), 1453 => to_unsigned(749, 10), 1454 => to_unsigned(1, 10), 1455 => to_unsigned(767, 10), 1456 => to_unsigned(764, 10), 1457 => to_unsigned(501, 10), 1458 => to_unsigned(805, 10), 1459 => to_unsigned(740, 10), 1460 => to_unsigned(870, 10), 1461 => to_unsigned(434, 10), 1462 => to_unsigned(633, 10), 1463 => to_unsigned(482, 10), 1464 => to_unsigned(872, 10), 1465 => to_unsigned(296, 10), 1466 => to_unsigned(482, 10), 1467 => to_unsigned(239, 10), 1468 => to_unsigned(154, 10), 1469 => to_unsigned(235, 10), 1470 => to_unsigned(729, 10), 1471 => to_unsigned(601, 10), 1472 => to_unsigned(569, 10), 1473 => to_unsigned(190, 10), 1474 => to_unsigned(646, 10), 1475 => to_unsigned(911, 10), 1476 => to_unsigned(570, 10), 1477 => to_unsigned(1015, 10), 1478 => to_unsigned(46, 10), 1479 => to_unsigned(350, 10), 1480 => to_unsigned(903, 10), 1481 => to_unsigned(205, 10), 1482 => to_unsigned(727, 10), 1483 => to_unsigned(236, 10), 1484 => to_unsigned(27, 10), 1485 => to_unsigned(842, 10), 1486 => to_unsigned(954, 10), 1487 => to_unsigned(420, 10), 1488 => to_unsigned(665, 10), 1489 => to_unsigned(1014, 10), 1490 => to_unsigned(334, 10), 1491 => to_unsigned(737, 10), 1492 => to_unsigned(888, 10), 1493 => to_unsigned(425, 10), 1494 => to_unsigned(183, 10), 1495 => to_unsigned(999, 10), 1496 => to_unsigned(870, 10), 1497 => to_unsigned(799, 10), 1498 => to_unsigned(633, 10), 1499 => to_unsigned(339, 10), 1500 => to_unsigned(522, 10), 1501 => to_unsigned(183, 10), 1502 => to_unsigned(409, 10), 1503 => to_unsigned(934, 10), 1504 => to_unsigned(712, 10), 1505 => to_unsigned(166, 10), 1506 => to_unsigned(136, 10), 1507 => to_unsigned(348, 10), 1508 => to_unsigned(564, 10), 1509 => to_unsigned(67, 10), 1510 => to_unsigned(328, 10), 1511 => to_unsigned(348, 10), 1512 => to_unsigned(938, 10), 1513 => to_unsigned(617, 10), 1514 => to_unsigned(190, 10), 1515 => to_unsigned(910, 10), 1516 => to_unsigned(273, 10), 1517 => to_unsigned(1001, 10), 1518 => to_unsigned(145, 10), 1519 => to_unsigned(650, 10), 1520 => to_unsigned(708, 10), 1521 => to_unsigned(895, 10), 1522 => to_unsigned(733, 10), 1523 => to_unsigned(544, 10), 1524 => to_unsigned(870, 10), 1525 => to_unsigned(696, 10), 1526 => to_unsigned(483, 10), 1527 => to_unsigned(77, 10), 1528 => to_unsigned(669, 10), 1529 => to_unsigned(958, 10), 1530 => to_unsigned(211, 10), 1531 => to_unsigned(236, 10), 1532 => to_unsigned(11, 10), 1533 => to_unsigned(677, 10), 1534 => to_unsigned(355, 10), 1535 => to_unsigned(771, 10), 1536 => to_unsigned(578, 10), 1537 => to_unsigned(122, 10), 1538 => to_unsigned(273, 10), 1539 => to_unsigned(193, 10), 1540 => to_unsigned(310, 10), 1541 => to_unsigned(257, 10), 1542 => to_unsigned(947, 10), 1543 => to_unsigned(779, 10), 1544 => to_unsigned(925, 10), 1545 => to_unsigned(130, 10), 1546 => to_unsigned(280, 10), 1547 => to_unsigned(695, 10), 1548 => to_unsigned(412, 10), 1549 => to_unsigned(285, 10), 1550 => to_unsigned(684, 10), 1551 => to_unsigned(196, 10), 1552 => to_unsigned(317, 10), 1553 => to_unsigned(798, 10), 1554 => to_unsigned(792, 10), 1555 => to_unsigned(935, 10), 1556 => to_unsigned(349, 10), 1557 => to_unsigned(532, 10), 1558 => to_unsigned(628, 10), 1559 => to_unsigned(854, 10), 1560 => to_unsigned(919, 10), 1561 => to_unsigned(267, 10), 1562 => to_unsigned(948, 10), 1563 => to_unsigned(605, 10), 1564 => to_unsigned(396, 10), 1565 => to_unsigned(750, 10), 1566 => to_unsigned(161, 10), 1567 => to_unsigned(3, 10), 1568 => to_unsigned(327, 10), 1569 => to_unsigned(826, 10), 1570 => to_unsigned(171, 10), 1571 => to_unsigned(357, 10), 1572 => to_unsigned(908, 10), 1573 => to_unsigned(24, 10), 1574 => to_unsigned(241, 10), 1575 => to_unsigned(986, 10), 1576 => to_unsigned(757, 10), 1577 => to_unsigned(15, 10), 1578 => to_unsigned(117, 10), 1579 => to_unsigned(662, 10), 1580 => to_unsigned(483, 10), 1581 => to_unsigned(353, 10), 1582 => to_unsigned(890, 10), 1583 => to_unsigned(592, 10), 1584 => to_unsigned(620, 10), 1585 => to_unsigned(125, 10), 1586 => to_unsigned(247, 10), 1587 => to_unsigned(192, 10), 1588 => to_unsigned(886, 10), 1589 => to_unsigned(196, 10), 1590 => to_unsigned(518, 10), 1591 => to_unsigned(434, 10), 1592 => to_unsigned(377, 10), 1593 => to_unsigned(926, 10), 1594 => to_unsigned(762, 10), 1595 => to_unsigned(723, 10), 1596 => to_unsigned(528, 10), 1597 => to_unsigned(81, 10), 1598 => to_unsigned(413, 10), 1599 => to_unsigned(365, 10), 1600 => to_unsigned(588, 10), 1601 => to_unsigned(330, 10), 1602 => to_unsigned(401, 10), 1603 => to_unsigned(501, 10), 1604 => to_unsigned(694, 10), 1605 => to_unsigned(994, 10), 1606 => to_unsigned(808, 10), 1607 => to_unsigned(472, 10), 1608 => to_unsigned(27, 10), 1609 => to_unsigned(546, 10), 1610 => to_unsigned(442, 10), 1611 => to_unsigned(782, 10), 1612 => to_unsigned(776, 10), 1613 => to_unsigned(52, 10), 1614 => to_unsigned(812, 10), 1615 => to_unsigned(914, 10), 1616 => to_unsigned(475, 10), 1617 => to_unsigned(218, 10), 1618 => to_unsigned(1010, 10), 1619 => to_unsigned(727, 10), 1620 => to_unsigned(455, 10), 1621 => to_unsigned(970, 10), 1622 => to_unsigned(962, 10), 1623 => to_unsigned(21, 10), 1624 => to_unsigned(716, 10), 1625 => to_unsigned(102, 10), 1626 => to_unsigned(395, 10), 1627 => to_unsigned(662, 10), 1628 => to_unsigned(956, 10), 1629 => to_unsigned(679, 10), 1630 => to_unsigned(461, 10), 1631 => to_unsigned(1017, 10), 1632 => to_unsigned(289, 10), 1633 => to_unsigned(1001, 10), 1634 => to_unsigned(984, 10), 1635 => to_unsigned(757, 10), 1636 => to_unsigned(251, 10), 1637 => to_unsigned(695, 10), 1638 => to_unsigned(471, 10), 1639 => to_unsigned(599, 10), 1640 => to_unsigned(220, 10), 1641 => to_unsigned(270, 10), 1642 => to_unsigned(989, 10), 1643 => to_unsigned(189, 10), 1644 => to_unsigned(427, 10), 1645 => to_unsigned(167, 10), 1646 => to_unsigned(961, 10), 1647 => to_unsigned(348, 10), 1648 => to_unsigned(757, 10), 1649 => to_unsigned(432, 10), 1650 => to_unsigned(574, 10), 1651 => to_unsigned(626, 10), 1652 => to_unsigned(758, 10), 1653 => to_unsigned(478, 10), 1654 => to_unsigned(143, 10), 1655 => to_unsigned(351, 10), 1656 => to_unsigned(412, 10), 1657 => to_unsigned(264, 10), 1658 => to_unsigned(356, 10), 1659 => to_unsigned(876, 10), 1660 => to_unsigned(467, 10), 1661 => to_unsigned(527, 10), 1662 => to_unsigned(1014, 10), 1663 => to_unsigned(82, 10), 1664 => to_unsigned(873, 10), 1665 => to_unsigned(699, 10), 1666 => to_unsigned(320, 10), 1667 => to_unsigned(576, 10), 1668 => to_unsigned(567, 10), 1669 => to_unsigned(689, 10), 1670 => to_unsigned(317, 10), 1671 => to_unsigned(961, 10), 1672 => to_unsigned(330, 10), 1673 => to_unsigned(222, 10), 1674 => to_unsigned(906, 10), 1675 => to_unsigned(419, 10), 1676 => to_unsigned(514, 10), 1677 => to_unsigned(769, 10), 1678 => to_unsigned(457, 10), 1679 => to_unsigned(1014, 10), 1680 => to_unsigned(938, 10), 1681 => to_unsigned(112, 10), 1682 => to_unsigned(884, 10), 1683 => to_unsigned(451, 10), 1684 => to_unsigned(494, 10), 1685 => to_unsigned(363, 10), 1686 => to_unsigned(36, 10), 1687 => to_unsigned(525, 10), 1688 => to_unsigned(163, 10), 1689 => to_unsigned(245, 10), 1690 => to_unsigned(783, 10), 1691 => to_unsigned(690, 10), 1692 => to_unsigned(878, 10), 1693 => to_unsigned(969, 10), 1694 => to_unsigned(871, 10), 1695 => to_unsigned(978, 10), 1696 => to_unsigned(962, 10), 1697 => to_unsigned(941, 10), 1698 => to_unsigned(553, 10), 1699 => to_unsigned(4, 10), 1700 => to_unsigned(764, 10), 1701 => to_unsigned(108, 10), 1702 => to_unsigned(462, 10), 1703 => to_unsigned(911, 10), 1704 => to_unsigned(108, 10), 1705 => to_unsigned(980, 10), 1706 => to_unsigned(473, 10), 1707 => to_unsigned(554, 10), 1708 => to_unsigned(978, 10), 1709 => to_unsigned(854, 10), 1710 => to_unsigned(916, 10), 1711 => to_unsigned(382, 10), 1712 => to_unsigned(491, 10), 1713 => to_unsigned(885, 10), 1714 => to_unsigned(302, 10), 1715 => to_unsigned(828, 10), 1716 => to_unsigned(1002, 10), 1717 => to_unsigned(818, 10), 1718 => to_unsigned(450, 10), 1719 => to_unsigned(967, 10), 1720 => to_unsigned(944, 10), 1721 => to_unsigned(914, 10), 1722 => to_unsigned(77, 10), 1723 => to_unsigned(321, 10), 1724 => to_unsigned(307, 10), 1725 => to_unsigned(372, 10), 1726 => to_unsigned(608, 10), 1727 => to_unsigned(451, 10), 1728 => to_unsigned(1014, 10), 1729 => to_unsigned(868, 10), 1730 => to_unsigned(176, 10), 1731 => to_unsigned(1008, 10), 1732 => to_unsigned(541, 10), 1733 => to_unsigned(67, 10), 1734 => to_unsigned(581, 10), 1735 => to_unsigned(667, 10), 1736 => to_unsigned(394, 10), 1737 => to_unsigned(52, 10), 1738 => to_unsigned(238, 10), 1739 => to_unsigned(774, 10), 1740 => to_unsigned(780, 10), 1741 => to_unsigned(321, 10), 1742 => to_unsigned(323, 10), 1743 => to_unsigned(703, 10), 1744 => to_unsigned(8, 10), 1745 => to_unsigned(356, 10), 1746 => to_unsigned(395, 10), 1747 => to_unsigned(465, 10), 1748 => to_unsigned(872, 10), 1749 => to_unsigned(34, 10), 1750 => to_unsigned(259, 10), 1751 => to_unsigned(673, 10), 1752 => to_unsigned(659, 10), 1753 => to_unsigned(643, 10), 1754 => to_unsigned(237, 10), 1755 => to_unsigned(93, 10), 1756 => to_unsigned(282, 10), 1757 => to_unsigned(731, 10), 1758 => to_unsigned(359, 10), 1759 => to_unsigned(499, 10), 1760 => to_unsigned(1008, 10), 1761 => to_unsigned(837, 10), 1762 => to_unsigned(662, 10), 1763 => to_unsigned(468, 10), 1764 => to_unsigned(589, 10), 1765 => to_unsigned(218, 10), 1766 => to_unsigned(927, 10), 1767 => to_unsigned(242, 10), 1768 => to_unsigned(38, 10), 1769 => to_unsigned(901, 10), 1770 => to_unsigned(689, 10), 1771 => to_unsigned(742, 10), 1772 => to_unsigned(137, 10), 1773 => to_unsigned(231, 10), 1774 => to_unsigned(349, 10), 1775 => to_unsigned(876, 10), 1776 => to_unsigned(184, 10), 1777 => to_unsigned(189, 10), 1778 => to_unsigned(648, 10), 1779 => to_unsigned(992, 10), 1780 => to_unsigned(946, 10), 1781 => to_unsigned(656, 10), 1782 => to_unsigned(405, 10), 1783 => to_unsigned(735, 10), 1784 => to_unsigned(107, 10), 1785 => to_unsigned(504, 10), 1786 => to_unsigned(248, 10), 1787 => to_unsigned(938, 10), 1788 => to_unsigned(965, 10), 1789 => to_unsigned(242, 10), 1790 => to_unsigned(131, 10), 1791 => to_unsigned(59, 10), 1792 => to_unsigned(88, 10), 1793 => to_unsigned(478, 10), 1794 => to_unsigned(11, 10), 1795 => to_unsigned(633, 10), 1796 => to_unsigned(748, 10), 1797 => to_unsigned(425, 10), 1798 => to_unsigned(547, 10), 1799 => to_unsigned(247, 10), 1800 => to_unsigned(538, 10), 1801 => to_unsigned(627, 10), 1802 => to_unsigned(176, 10), 1803 => to_unsigned(130, 10), 1804 => to_unsigned(390, 10), 1805 => to_unsigned(305, 10), 1806 => to_unsigned(623, 10), 1807 => to_unsigned(11, 10), 1808 => to_unsigned(42, 10), 1809 => to_unsigned(533, 10), 1810 => to_unsigned(126, 10), 1811 => to_unsigned(789, 10), 1812 => to_unsigned(80, 10), 1813 => to_unsigned(776, 10), 1814 => to_unsigned(215, 10), 1815 => to_unsigned(871, 10), 1816 => to_unsigned(1008, 10), 1817 => to_unsigned(725, 10), 1818 => to_unsigned(960, 10), 1819 => to_unsigned(485, 10), 1820 => to_unsigned(239, 10), 1821 => to_unsigned(523, 10), 1822 => to_unsigned(675, 10), 1823 => to_unsigned(738, 10), 1824 => to_unsigned(346, 10), 1825 => to_unsigned(544, 10), 1826 => to_unsigned(97, 10), 1827 => to_unsigned(107, 10), 1828 => to_unsigned(764, 10), 1829 => to_unsigned(470, 10), 1830 => to_unsigned(403, 10), 1831 => to_unsigned(1000, 10), 1832 => to_unsigned(486, 10), 1833 => to_unsigned(565, 10), 1834 => to_unsigned(744, 10), 1835 => to_unsigned(56, 10), 1836 => to_unsigned(509, 10), 1837 => to_unsigned(701, 10), 1838 => to_unsigned(441, 10), 1839 => to_unsigned(66, 10), 1840 => to_unsigned(604, 10), 1841 => to_unsigned(544, 10), 1842 => to_unsigned(263, 10), 1843 => to_unsigned(253, 10), 1844 => to_unsigned(655, 10), 1845 => to_unsigned(619, 10), 1846 => to_unsigned(863, 10), 1847 => to_unsigned(1009, 10), 1848 => to_unsigned(734, 10), 1849 => to_unsigned(428, 10), 1850 => to_unsigned(469, 10), 1851 => to_unsigned(209, 10), 1852 => to_unsigned(205, 10), 1853 => to_unsigned(482, 10), 1854 => to_unsigned(816, 10), 1855 => to_unsigned(987, 10), 1856 => to_unsigned(200, 10), 1857 => to_unsigned(676, 10), 1858 => to_unsigned(468, 10), 1859 => to_unsigned(612, 10), 1860 => to_unsigned(666, 10), 1861 => to_unsigned(823, 10), 1862 => to_unsigned(37, 10), 1863 => to_unsigned(178, 10), 1864 => to_unsigned(620, 10), 1865 => to_unsigned(674, 10), 1866 => to_unsigned(10, 10), 1867 => to_unsigned(735, 10), 1868 => to_unsigned(340, 10), 1869 => to_unsigned(783, 10), 1870 => to_unsigned(875, 10), 1871 => to_unsigned(45, 10), 1872 => to_unsigned(889, 10), 1873 => to_unsigned(682, 10), 1874 => to_unsigned(279, 10), 1875 => to_unsigned(444, 10), 1876 => to_unsigned(942, 10), 1877 => to_unsigned(779, 10), 1878 => to_unsigned(917, 10), 1879 => to_unsigned(522, 10), 1880 => to_unsigned(961, 10), 1881 => to_unsigned(579, 10), 1882 => to_unsigned(307, 10), 1883 => to_unsigned(889, 10), 1884 => to_unsigned(292, 10), 1885 => to_unsigned(305, 10), 1886 => to_unsigned(481, 10), 1887 => to_unsigned(892, 10), 1888 => to_unsigned(452, 10), 1889 => to_unsigned(712, 10), 1890 => to_unsigned(323, 10), 1891 => to_unsigned(867, 10), 1892 => to_unsigned(847, 10), 1893 => to_unsigned(820, 10), 1894 => to_unsigned(350, 10), 1895 => to_unsigned(168, 10), 1896 => to_unsigned(895, 10), 1897 => to_unsigned(849, 10), 1898 => to_unsigned(801, 10), 1899 => to_unsigned(530, 10), 1900 => to_unsigned(639, 10), 1901 => to_unsigned(323, 10), 1902 => to_unsigned(1017, 10), 1903 => to_unsigned(533, 10), 1904 => to_unsigned(696, 10), 1905 => to_unsigned(563, 10), 1906 => to_unsigned(500, 10), 1907 => to_unsigned(237, 10), 1908 => to_unsigned(726, 10), 1909 => to_unsigned(464, 10), 1910 => to_unsigned(718, 10), 1911 => to_unsigned(729, 10), 1912 => to_unsigned(525, 10), 1913 => to_unsigned(387, 10), 1914 => to_unsigned(985, 10), 1915 => to_unsigned(762, 10), 1916 => to_unsigned(465, 10), 1917 => to_unsigned(460, 10), 1918 => to_unsigned(29, 10), 1919 => to_unsigned(686, 10), 1920 => to_unsigned(173, 10), 1921 => to_unsigned(217, 10), 1922 => to_unsigned(325, 10), 1923 => to_unsigned(492, 10), 1924 => to_unsigned(520, 10), 1925 => to_unsigned(942, 10), 1926 => to_unsigned(249, 10), 1927 => to_unsigned(176, 10), 1928 => to_unsigned(250, 10), 1929 => to_unsigned(704, 10), 1930 => to_unsigned(66, 10), 1931 => to_unsigned(61, 10), 1932 => to_unsigned(393, 10), 1933 => to_unsigned(11, 10), 1934 => to_unsigned(319, 10), 1935 => to_unsigned(799, 10), 1936 => to_unsigned(918, 10), 1937 => to_unsigned(801, 10), 1938 => to_unsigned(447, 10), 1939 => to_unsigned(943, 10), 1940 => to_unsigned(84, 10), 1941 => to_unsigned(713, 10), 1942 => to_unsigned(854, 10), 1943 => to_unsigned(347, 10), 1944 => to_unsigned(329, 10), 1945 => to_unsigned(147, 10), 1946 => to_unsigned(983, 10), 1947 => to_unsigned(185, 10), 1948 => to_unsigned(951, 10), 1949 => to_unsigned(820, 10), 1950 => to_unsigned(252, 10), 1951 => to_unsigned(984, 10), 1952 => to_unsigned(372, 10), 1953 => to_unsigned(217, 10), 1954 => to_unsigned(626, 10), 1955 => to_unsigned(198, 10), 1956 => to_unsigned(819, 10), 1957 => to_unsigned(291, 10), 1958 => to_unsigned(592, 10), 1959 => to_unsigned(479, 10), 1960 => to_unsigned(545, 10), 1961 => to_unsigned(389, 10), 1962 => to_unsigned(700, 10), 1963 => to_unsigned(909, 10), 1964 => to_unsigned(267, 10), 1965 => to_unsigned(363, 10), 1966 => to_unsigned(683, 10), 1967 => to_unsigned(965, 10), 1968 => to_unsigned(458, 10), 1969 => to_unsigned(210, 10), 1970 => to_unsigned(834, 10), 1971 => to_unsigned(702, 10), 1972 => to_unsigned(119, 10), 1973 => to_unsigned(656, 10), 1974 => to_unsigned(256, 10), 1975 => to_unsigned(269, 10), 1976 => to_unsigned(48, 10), 1977 => to_unsigned(918, 10), 1978 => to_unsigned(929, 10), 1979 => to_unsigned(768, 10), 1980 => to_unsigned(490, 10), 1981 => to_unsigned(585, 10), 1982 => to_unsigned(665, 10), 1983 => to_unsigned(104, 10), 1984 => to_unsigned(313, 10), 1985 => to_unsigned(570, 10), 1986 => to_unsigned(450, 10), 1987 => to_unsigned(526, 10), 1988 => to_unsigned(374, 10), 1989 => to_unsigned(826, 10), 1990 => to_unsigned(924, 10), 1991 => to_unsigned(725, 10), 1992 => to_unsigned(962, 10), 1993 => to_unsigned(406, 10), 1994 => to_unsigned(509, 10), 1995 => to_unsigned(200, 10), 1996 => to_unsigned(239, 10), 1997 => to_unsigned(464, 10), 1998 => to_unsigned(291, 10), 1999 => to_unsigned(493, 10), 2000 => to_unsigned(923, 10), 2001 => to_unsigned(866, 10), 2002 => to_unsigned(313, 10), 2003 => to_unsigned(647, 10), 2004 => to_unsigned(925, 10), 2005 => to_unsigned(394, 10), 2006 => to_unsigned(605, 10), 2007 => to_unsigned(71, 10), 2008 => to_unsigned(496, 10), 2009 => to_unsigned(135, 10), 2010 => to_unsigned(833, 10), 2011 => to_unsigned(409, 10), 2012 => to_unsigned(909, 10), 2013 => to_unsigned(205, 10), 2014 => to_unsigned(192, 10), 2015 => to_unsigned(809, 10), 2016 => to_unsigned(684, 10), 2017 => to_unsigned(147, 10), 2018 => to_unsigned(323, 10), 2019 => to_unsigned(889, 10), 2020 => to_unsigned(167, 10), 2021 => to_unsigned(117, 10), 2022 => to_unsigned(321, 10), 2023 => to_unsigned(81, 10), 2024 => to_unsigned(59, 10), 2025 => to_unsigned(246, 10), 2026 => to_unsigned(738, 10), 2027 => to_unsigned(106, 10), 2028 => to_unsigned(261, 10), 2029 => to_unsigned(834, 10), 2030 => to_unsigned(843, 10), 2031 => to_unsigned(63, 10), 2032 => to_unsigned(747, 10), 2033 => to_unsigned(965, 10), 2034 => to_unsigned(458, 10), 2035 => to_unsigned(1012, 10), 2036 => to_unsigned(644, 10), 2037 => to_unsigned(301, 10), 2038 => to_unsigned(383, 10), 2039 => to_unsigned(288, 10), 2040 => to_unsigned(308, 10), 2041 => to_unsigned(944, 10), 2042 => to_unsigned(723, 10), 2043 => to_unsigned(342, 10), 2044 => to_unsigned(68, 10), 2045 => to_unsigned(405, 10), 2046 => to_unsigned(995, 10), 2047 => to_unsigned(460, 10)),
            1 => (0 => to_unsigned(671, 10), 1 => to_unsigned(352, 10), 2 => to_unsigned(731, 10), 3 => to_unsigned(573, 10), 4 => to_unsigned(717, 10), 5 => to_unsigned(670, 10), 6 => to_unsigned(82, 10), 7 => to_unsigned(331, 10), 8 => to_unsigned(992, 10), 9 => to_unsigned(694, 10), 10 => to_unsigned(370, 10), 11 => to_unsigned(779, 10), 12 => to_unsigned(82, 10), 13 => to_unsigned(369, 10), 14 => to_unsigned(112, 10), 15 => to_unsigned(732, 10), 16 => to_unsigned(491, 10), 17 => to_unsigned(530, 10), 18 => to_unsigned(213, 10), 19 => to_unsigned(451, 10), 20 => to_unsigned(925, 10), 21 => to_unsigned(545, 10), 22 => to_unsigned(941, 10), 23 => to_unsigned(632, 10), 24 => to_unsigned(42, 10), 25 => to_unsigned(221, 10), 26 => to_unsigned(715, 10), 27 => to_unsigned(979, 10), 28 => to_unsigned(1011, 10), 29 => to_unsigned(56, 10), 30 => to_unsigned(978, 10), 31 => to_unsigned(35, 10), 32 => to_unsigned(173, 10), 33 => to_unsigned(486, 10), 34 => to_unsigned(687, 10), 35 => to_unsigned(770, 10), 36 => to_unsigned(643, 10), 37 => to_unsigned(58, 10), 38 => to_unsigned(899, 10), 39 => to_unsigned(980, 10), 40 => to_unsigned(166, 10), 41 => to_unsigned(272, 10), 42 => to_unsigned(607, 10), 43 => to_unsigned(141, 10), 44 => to_unsigned(495, 10), 45 => to_unsigned(779, 10), 46 => to_unsigned(481, 10), 47 => to_unsigned(733, 10), 48 => to_unsigned(594, 10), 49 => to_unsigned(842, 10), 50 => to_unsigned(109, 10), 51 => to_unsigned(88, 10), 52 => to_unsigned(368, 10), 53 => to_unsigned(916, 10), 54 => to_unsigned(706, 10), 55 => to_unsigned(81, 10), 56 => to_unsigned(330, 10), 57 => to_unsigned(156, 10), 58 => to_unsigned(732, 10), 59 => to_unsigned(755, 10), 60 => to_unsigned(101, 10), 61 => to_unsigned(969, 10), 62 => to_unsigned(132, 10), 63 => to_unsigned(975, 10), 64 => to_unsigned(439, 10), 65 => to_unsigned(732, 10), 66 => to_unsigned(684, 10), 67 => to_unsigned(268, 10), 68 => to_unsigned(194, 10), 69 => to_unsigned(95, 10), 70 => to_unsigned(680, 10), 71 => to_unsigned(319, 10), 72 => to_unsigned(116, 10), 73 => to_unsigned(571, 10), 74 => to_unsigned(482, 10), 75 => to_unsigned(401, 10), 76 => to_unsigned(72, 10), 77 => to_unsigned(354, 10), 78 => to_unsigned(670, 10), 79 => to_unsigned(456, 10), 80 => to_unsigned(398, 10), 81 => to_unsigned(25, 10), 82 => to_unsigned(525, 10), 83 => to_unsigned(425, 10), 84 => to_unsigned(278, 10), 85 => to_unsigned(356, 10), 86 => to_unsigned(740, 10), 87 => to_unsigned(81, 10), 88 => to_unsigned(708, 10), 89 => to_unsigned(512, 10), 90 => to_unsigned(534, 10), 91 => to_unsigned(420, 10), 92 => to_unsigned(865, 10), 93 => to_unsigned(395, 10), 94 => to_unsigned(892, 10), 95 => to_unsigned(564, 10), 96 => to_unsigned(118, 10), 97 => to_unsigned(644, 10), 98 => to_unsigned(498, 10), 99 => to_unsigned(1004, 10), 100 => to_unsigned(327, 10), 101 => to_unsigned(706, 10), 102 => to_unsigned(76, 10), 103 => to_unsigned(767, 10), 104 => to_unsigned(143, 10), 105 => to_unsigned(792, 10), 106 => to_unsigned(2, 10), 107 => to_unsigned(97, 10), 108 => to_unsigned(507, 10), 109 => to_unsigned(721, 10), 110 => to_unsigned(112, 10), 111 => to_unsigned(35, 10), 112 => to_unsigned(270, 10), 113 => to_unsigned(251, 10), 114 => to_unsigned(458, 10), 115 => to_unsigned(817, 10), 116 => to_unsigned(949, 10), 117 => to_unsigned(1002, 10), 118 => to_unsigned(623, 10), 119 => to_unsigned(1022, 10), 120 => to_unsigned(176, 10), 121 => to_unsigned(232, 10), 122 => to_unsigned(71, 10), 123 => to_unsigned(74, 10), 124 => to_unsigned(1021, 10), 125 => to_unsigned(61, 10), 126 => to_unsigned(671, 10), 127 => to_unsigned(207, 10), 128 => to_unsigned(984, 10), 129 => to_unsigned(785, 10), 130 => to_unsigned(758, 10), 131 => to_unsigned(571, 10), 132 => to_unsigned(656, 10), 133 => to_unsigned(856, 10), 134 => to_unsigned(342, 10), 135 => to_unsigned(940, 10), 136 => to_unsigned(842, 10), 137 => to_unsigned(230, 10), 138 => to_unsigned(277, 10), 139 => to_unsigned(761, 10), 140 => to_unsigned(823, 10), 141 => to_unsigned(832, 10), 142 => to_unsigned(198, 10), 143 => to_unsigned(239, 10), 144 => to_unsigned(500, 10), 145 => to_unsigned(58, 10), 146 => to_unsigned(432, 10), 147 => to_unsigned(435, 10), 148 => to_unsigned(732, 10), 149 => to_unsigned(592, 10), 150 => to_unsigned(179, 10), 151 => to_unsigned(189, 10), 152 => to_unsigned(263, 10), 153 => to_unsigned(1006, 10), 154 => to_unsigned(197, 10), 155 => to_unsigned(641, 10), 156 => to_unsigned(512, 10), 157 => to_unsigned(739, 10), 158 => to_unsigned(965, 10), 159 => to_unsigned(11, 10), 160 => to_unsigned(967, 10), 161 => to_unsigned(112, 10), 162 => to_unsigned(834, 10), 163 => to_unsigned(563, 10), 164 => to_unsigned(831, 10), 165 => to_unsigned(849, 10), 166 => to_unsigned(609, 10), 167 => to_unsigned(508, 10), 168 => to_unsigned(431, 10), 169 => to_unsigned(715, 10), 170 => to_unsigned(567, 10), 171 => to_unsigned(236, 10), 172 => to_unsigned(307, 10), 173 => to_unsigned(847, 10), 174 => to_unsigned(417, 10), 175 => to_unsigned(220, 10), 176 => to_unsigned(564, 10), 177 => to_unsigned(107, 10), 178 => to_unsigned(534, 10), 179 => to_unsigned(629, 10), 180 => to_unsigned(910, 10), 181 => to_unsigned(4, 10), 182 => to_unsigned(351, 10), 183 => to_unsigned(294, 10), 184 => to_unsigned(429, 10), 185 => to_unsigned(353, 10), 186 => to_unsigned(839, 10), 187 => to_unsigned(893, 10), 188 => to_unsigned(740, 10), 189 => to_unsigned(708, 10), 190 => to_unsigned(244, 10), 191 => to_unsigned(358, 10), 192 => to_unsigned(121, 10), 193 => to_unsigned(554, 10), 194 => to_unsigned(157, 10), 195 => to_unsigned(767, 10), 196 => to_unsigned(500, 10), 197 => to_unsigned(59, 10), 198 => to_unsigned(905, 10), 199 => to_unsigned(223, 10), 200 => to_unsigned(436, 10), 201 => to_unsigned(53, 10), 202 => to_unsigned(361, 10), 203 => to_unsigned(262, 10), 204 => to_unsigned(616, 10), 205 => to_unsigned(871, 10), 206 => to_unsigned(662, 10), 207 => to_unsigned(626, 10), 208 => to_unsigned(784, 10), 209 => to_unsigned(348, 10), 210 => to_unsigned(527, 10), 211 => to_unsigned(38, 10), 212 => to_unsigned(905, 10), 213 => to_unsigned(668, 10), 214 => to_unsigned(308, 10), 215 => to_unsigned(909, 10), 216 => to_unsigned(327, 10), 217 => to_unsigned(55, 10), 218 => to_unsigned(566, 10), 219 => to_unsigned(43, 10), 220 => to_unsigned(186, 10), 221 => to_unsigned(983, 10), 222 => to_unsigned(875, 10), 223 => to_unsigned(182, 10), 224 => to_unsigned(618, 10), 225 => to_unsigned(881, 10), 226 => to_unsigned(378, 10), 227 => to_unsigned(466, 10), 228 => to_unsigned(123, 10), 229 => to_unsigned(630, 10), 230 => to_unsigned(65, 10), 231 => to_unsigned(479, 10), 232 => to_unsigned(357, 10), 233 => to_unsigned(306, 10), 234 => to_unsigned(90, 10), 235 => to_unsigned(816, 10), 236 => to_unsigned(234, 10), 237 => to_unsigned(484, 10), 238 => to_unsigned(428, 10), 239 => to_unsigned(157, 10), 240 => to_unsigned(747, 10), 241 => to_unsigned(930, 10), 242 => to_unsigned(609, 10), 243 => to_unsigned(109, 10), 244 => to_unsigned(784, 10), 245 => to_unsigned(485, 10), 246 => to_unsigned(93, 10), 247 => to_unsigned(896, 10), 248 => to_unsigned(515, 10), 249 => to_unsigned(563, 10), 250 => to_unsigned(210, 10), 251 => to_unsigned(651, 10), 252 => to_unsigned(357, 10), 253 => to_unsigned(453, 10), 254 => to_unsigned(608, 10), 255 => to_unsigned(1000, 10), 256 => to_unsigned(876, 10), 257 => to_unsigned(931, 10), 258 => to_unsigned(379, 10), 259 => to_unsigned(357, 10), 260 => to_unsigned(581, 10), 261 => to_unsigned(808, 10), 262 => to_unsigned(690, 10), 263 => to_unsigned(216, 10), 264 => to_unsigned(74, 10), 265 => to_unsigned(746, 10), 266 => to_unsigned(459, 10), 267 => to_unsigned(371, 10), 268 => to_unsigned(959, 10), 269 => to_unsigned(98, 10), 270 => to_unsigned(500, 10), 271 => to_unsigned(409, 10), 272 => to_unsigned(233, 10), 273 => to_unsigned(165, 10), 274 => to_unsigned(227, 10), 275 => to_unsigned(27, 10), 276 => to_unsigned(709, 10), 277 => to_unsigned(238, 10), 278 => to_unsigned(739, 10), 279 => to_unsigned(843, 10), 280 => to_unsigned(870, 10), 281 => to_unsigned(82, 10), 282 => to_unsigned(955, 10), 283 => to_unsigned(15, 10), 284 => to_unsigned(886, 10), 285 => to_unsigned(602, 10), 286 => to_unsigned(10, 10), 287 => to_unsigned(524, 10), 288 => to_unsigned(592, 10), 289 => to_unsigned(611, 10), 290 => to_unsigned(606, 10), 291 => to_unsigned(45, 10), 292 => to_unsigned(896, 10), 293 => to_unsigned(458, 10), 294 => to_unsigned(132, 10), 295 => to_unsigned(384, 10), 296 => to_unsigned(76, 10), 297 => to_unsigned(690, 10), 298 => to_unsigned(1021, 10), 299 => to_unsigned(949, 10), 300 => to_unsigned(383, 10), 301 => to_unsigned(495, 10), 302 => to_unsigned(203, 10), 303 => to_unsigned(328, 10), 304 => to_unsigned(971, 10), 305 => to_unsigned(160, 10), 306 => to_unsigned(31, 10), 307 => to_unsigned(893, 10), 308 => to_unsigned(783, 10), 309 => to_unsigned(807, 10), 310 => to_unsigned(213, 10), 311 => to_unsigned(238, 10), 312 => to_unsigned(50, 10), 313 => to_unsigned(123, 10), 314 => to_unsigned(653, 10), 315 => to_unsigned(528, 10), 316 => to_unsigned(731, 10), 317 => to_unsigned(718, 10), 318 => to_unsigned(519, 10), 319 => to_unsigned(531, 10), 320 => to_unsigned(806, 10), 321 => to_unsigned(243, 10), 322 => to_unsigned(190, 10), 323 => to_unsigned(819, 10), 324 => to_unsigned(761, 10), 325 => to_unsigned(901, 10), 326 => to_unsigned(89, 10), 327 => to_unsigned(342, 10), 328 => to_unsigned(836, 10), 329 => to_unsigned(542, 10), 330 => to_unsigned(799, 10), 331 => to_unsigned(856, 10), 332 => to_unsigned(134, 10), 333 => to_unsigned(900, 10), 334 => to_unsigned(577, 10), 335 => to_unsigned(585, 10), 336 => to_unsigned(492, 10), 337 => to_unsigned(976, 10), 338 => to_unsigned(452, 10), 339 => to_unsigned(708, 10), 340 => to_unsigned(896, 10), 341 => to_unsigned(22, 10), 342 => to_unsigned(908, 10), 343 => to_unsigned(402, 10), 344 => to_unsigned(611, 10), 345 => to_unsigned(14, 10), 346 => to_unsigned(365, 10), 347 => to_unsigned(813, 10), 348 => to_unsigned(981, 10), 349 => to_unsigned(38, 10), 350 => to_unsigned(9, 10), 351 => to_unsigned(627, 10), 352 => to_unsigned(809, 10), 353 => to_unsigned(688, 10), 354 => to_unsigned(501, 10), 355 => to_unsigned(835, 10), 356 => to_unsigned(525, 10), 357 => to_unsigned(503, 10), 358 => to_unsigned(846, 10), 359 => to_unsigned(567, 10), 360 => to_unsigned(135, 10), 361 => to_unsigned(441, 10), 362 => to_unsigned(793, 10), 363 => to_unsigned(486, 10), 364 => to_unsigned(185, 10), 365 => to_unsigned(15, 10), 366 => to_unsigned(634, 10), 367 => to_unsigned(486, 10), 368 => to_unsigned(256, 10), 369 => to_unsigned(676, 10), 370 => to_unsigned(835, 10), 371 => to_unsigned(502, 10), 372 => to_unsigned(872, 10), 373 => to_unsigned(675, 10), 374 => to_unsigned(714, 10), 375 => to_unsigned(261, 10), 376 => to_unsigned(972, 10), 377 => to_unsigned(542, 10), 378 => to_unsigned(116, 10), 379 => to_unsigned(361, 10), 380 => to_unsigned(195, 10), 381 => to_unsigned(619, 10), 382 => to_unsigned(690, 10), 383 => to_unsigned(953, 10), 384 => to_unsigned(847, 10), 385 => to_unsigned(334, 10), 386 => to_unsigned(561, 10), 387 => to_unsigned(299, 10), 388 => to_unsigned(311, 10), 389 => to_unsigned(320, 10), 390 => to_unsigned(749, 10), 391 => to_unsigned(915, 10), 392 => to_unsigned(539, 10), 393 => to_unsigned(759, 10), 394 => to_unsigned(216, 10), 395 => to_unsigned(115, 10), 396 => to_unsigned(240, 10), 397 => to_unsigned(954, 10), 398 => to_unsigned(232, 10), 399 => to_unsigned(296, 10), 400 => to_unsigned(765, 10), 401 => to_unsigned(909, 10), 402 => to_unsigned(788, 10), 403 => to_unsigned(279, 10), 404 => to_unsigned(913, 10), 405 => to_unsigned(887, 10), 406 => to_unsigned(511, 10), 407 => to_unsigned(801, 10), 408 => to_unsigned(274, 10), 409 => to_unsigned(36, 10), 410 => to_unsigned(743, 10), 411 => to_unsigned(58, 10), 412 => to_unsigned(105, 10), 413 => to_unsigned(94, 10), 414 => to_unsigned(2, 10), 415 => to_unsigned(35, 10), 416 => to_unsigned(804, 10), 417 => to_unsigned(823, 10), 418 => to_unsigned(659, 10), 419 => to_unsigned(136, 10), 420 => to_unsigned(754, 10), 421 => to_unsigned(23, 10), 422 => to_unsigned(43, 10), 423 => to_unsigned(386, 10), 424 => to_unsigned(135, 10), 425 => to_unsigned(20, 10), 426 => to_unsigned(242, 10), 427 => to_unsigned(263, 10), 428 => to_unsigned(755, 10), 429 => to_unsigned(888, 10), 430 => to_unsigned(639, 10), 431 => to_unsigned(184, 10), 432 => to_unsigned(176, 10), 433 => to_unsigned(763, 10), 434 => to_unsigned(394, 10), 435 => to_unsigned(310, 10), 436 => to_unsigned(848, 10), 437 => to_unsigned(766, 10), 438 => to_unsigned(192, 10), 439 => to_unsigned(707, 10), 440 => to_unsigned(295, 10), 441 => to_unsigned(719, 10), 442 => to_unsigned(415, 10), 443 => to_unsigned(64, 10), 444 => to_unsigned(830, 10), 445 => to_unsigned(106, 10), 446 => to_unsigned(360, 10), 447 => to_unsigned(299, 10), 448 => to_unsigned(1001, 10), 449 => to_unsigned(815, 10), 450 => to_unsigned(165, 10), 451 => to_unsigned(588, 10), 452 => to_unsigned(404, 10), 453 => to_unsigned(426, 10), 454 => to_unsigned(352, 10), 455 => to_unsigned(94, 10), 456 => to_unsigned(185, 10), 457 => to_unsigned(169, 10), 458 => to_unsigned(852, 10), 459 => to_unsigned(972, 10), 460 => to_unsigned(586, 10), 461 => to_unsigned(7, 10), 462 => to_unsigned(587, 10), 463 => to_unsigned(581, 10), 464 => to_unsigned(518, 10), 465 => to_unsigned(617, 10), 466 => to_unsigned(42, 10), 467 => to_unsigned(731, 10), 468 => to_unsigned(876, 10), 469 => to_unsigned(217, 10), 470 => to_unsigned(804, 10), 471 => to_unsigned(1016, 10), 472 => to_unsigned(324, 10), 473 => to_unsigned(299, 10), 474 => to_unsigned(176, 10), 475 => to_unsigned(644, 10), 476 => to_unsigned(381, 10), 477 => to_unsigned(1003, 10), 478 => to_unsigned(549, 10), 479 => to_unsigned(837, 10), 480 => to_unsigned(72, 10), 481 => to_unsigned(334, 10), 482 => to_unsigned(598, 10), 483 => to_unsigned(984, 10), 484 => to_unsigned(697, 10), 485 => to_unsigned(971, 10), 486 => to_unsigned(907, 10), 487 => to_unsigned(804, 10), 488 => to_unsigned(246, 10), 489 => to_unsigned(255, 10), 490 => to_unsigned(969, 10), 491 => to_unsigned(815, 10), 492 => to_unsigned(52, 10), 493 => to_unsigned(807, 10), 494 => to_unsigned(64, 10), 495 => to_unsigned(69, 10), 496 => to_unsigned(335, 10), 497 => to_unsigned(373, 10), 498 => to_unsigned(343, 10), 499 => to_unsigned(274, 10), 500 => to_unsigned(377, 10), 501 => to_unsigned(117, 10), 502 => to_unsigned(694, 10), 503 => to_unsigned(777, 10), 504 => to_unsigned(662, 10), 505 => to_unsigned(41, 10), 506 => to_unsigned(913, 10), 507 => to_unsigned(912, 10), 508 => to_unsigned(890, 10), 509 => to_unsigned(341, 10), 510 => to_unsigned(811, 10), 511 => to_unsigned(946, 10), 512 => to_unsigned(695, 10), 513 => to_unsigned(801, 10), 514 => to_unsigned(85, 10), 515 => to_unsigned(586, 10), 516 => to_unsigned(689, 10), 517 => to_unsigned(79, 10), 518 => to_unsigned(368, 10), 519 => to_unsigned(664, 10), 520 => to_unsigned(799, 10), 521 => to_unsigned(36, 10), 522 => to_unsigned(20, 10), 523 => to_unsigned(180, 10), 524 => to_unsigned(575, 10), 525 => to_unsigned(637, 10), 526 => to_unsigned(180, 10), 527 => to_unsigned(954, 10), 528 => to_unsigned(611, 10), 529 => to_unsigned(6, 10), 530 => to_unsigned(299, 10), 531 => to_unsigned(339, 10), 532 => to_unsigned(972, 10), 533 => to_unsigned(756, 10), 534 => to_unsigned(287, 10), 535 => to_unsigned(258, 10), 536 => to_unsigned(792, 10), 537 => to_unsigned(555, 10), 538 => to_unsigned(702, 10), 539 => to_unsigned(577, 10), 540 => to_unsigned(157, 10), 541 => to_unsigned(798, 10), 542 => to_unsigned(410, 10), 543 => to_unsigned(389, 10), 544 => to_unsigned(738, 10), 545 => to_unsigned(440, 10), 546 => to_unsigned(969, 10), 547 => to_unsigned(392, 10), 548 => to_unsigned(376, 10), 549 => to_unsigned(618, 10), 550 => to_unsigned(313, 10), 551 => to_unsigned(717, 10), 552 => to_unsigned(382, 10), 553 => to_unsigned(874, 10), 554 => to_unsigned(863, 10), 555 => to_unsigned(432, 10), 556 => to_unsigned(343, 10), 557 => to_unsigned(505, 10), 558 => to_unsigned(424, 10), 559 => to_unsigned(141, 10), 560 => to_unsigned(66, 10), 561 => to_unsigned(1010, 10), 562 => to_unsigned(214, 10), 563 => to_unsigned(684, 10), 564 => to_unsigned(181, 10), 565 => to_unsigned(761, 10), 566 => to_unsigned(657, 10), 567 => to_unsigned(837, 10), 568 => to_unsigned(573, 10), 569 => to_unsigned(975, 10), 570 => to_unsigned(697, 10), 571 => to_unsigned(174, 10), 572 => to_unsigned(88, 10), 573 => to_unsigned(531, 10), 574 => to_unsigned(900, 10), 575 => to_unsigned(871, 10), 576 => to_unsigned(0, 10), 577 => to_unsigned(448, 10), 578 => to_unsigned(743, 10), 579 => to_unsigned(235, 10), 580 => to_unsigned(970, 10), 581 => to_unsigned(120, 10), 582 => to_unsigned(605, 10), 583 => to_unsigned(344, 10), 584 => to_unsigned(137, 10), 585 => to_unsigned(139, 10), 586 => to_unsigned(724, 10), 587 => to_unsigned(444, 10), 588 => to_unsigned(577, 10), 589 => to_unsigned(779, 10), 590 => to_unsigned(517, 10), 591 => to_unsigned(986, 10), 592 => to_unsigned(653, 10), 593 => to_unsigned(515, 10), 594 => to_unsigned(224, 10), 595 => to_unsigned(608, 10), 596 => to_unsigned(260, 10), 597 => to_unsigned(492, 10), 598 => to_unsigned(356, 10), 599 => to_unsigned(420, 10), 600 => to_unsigned(449, 10), 601 => to_unsigned(929, 10), 602 => to_unsigned(1017, 10), 603 => to_unsigned(347, 10), 604 => to_unsigned(824, 10), 605 => to_unsigned(630, 10), 606 => to_unsigned(875, 10), 607 => to_unsigned(375, 10), 608 => to_unsigned(43, 10), 609 => to_unsigned(474, 10), 610 => to_unsigned(21, 10), 611 => to_unsigned(808, 10), 612 => to_unsigned(534, 10), 613 => to_unsigned(355, 10), 614 => to_unsigned(206, 10), 615 => to_unsigned(203, 10), 616 => to_unsigned(852, 10), 617 => to_unsigned(183, 10), 618 => to_unsigned(15, 10), 619 => to_unsigned(194, 10), 620 => to_unsigned(82, 10), 621 => to_unsigned(841, 10), 622 => to_unsigned(222, 10), 623 => to_unsigned(215, 10), 624 => to_unsigned(310, 10), 625 => to_unsigned(945, 10), 626 => to_unsigned(440, 10), 627 => to_unsigned(281, 10), 628 => to_unsigned(391, 10), 629 => to_unsigned(758, 10), 630 => to_unsigned(138, 10), 631 => to_unsigned(87, 10), 632 => to_unsigned(934, 10), 633 => to_unsigned(68, 10), 634 => to_unsigned(52, 10), 635 => to_unsigned(784, 10), 636 => to_unsigned(973, 10), 637 => to_unsigned(1009, 10), 638 => to_unsigned(510, 10), 639 => to_unsigned(800, 10), 640 => to_unsigned(199, 10), 641 => to_unsigned(366, 10), 642 => to_unsigned(865, 10), 643 => to_unsigned(799, 10), 644 => to_unsigned(354, 10), 645 => to_unsigned(924, 10), 646 => to_unsigned(877, 10), 647 => to_unsigned(766, 10), 648 => to_unsigned(698, 10), 649 => to_unsigned(429, 10), 650 => to_unsigned(848, 10), 651 => to_unsigned(903, 10), 652 => to_unsigned(438, 10), 653 => to_unsigned(474, 10), 654 => to_unsigned(755, 10), 655 => to_unsigned(25, 10), 656 => to_unsigned(87, 10), 657 => to_unsigned(518, 10), 658 => to_unsigned(542, 10), 659 => to_unsigned(139, 10), 660 => to_unsigned(113, 10), 661 => to_unsigned(23, 10), 662 => to_unsigned(468, 10), 663 => to_unsigned(71, 10), 664 => to_unsigned(320, 10), 665 => to_unsigned(238, 10), 666 => to_unsigned(635, 10), 667 => to_unsigned(462, 10), 668 => to_unsigned(330, 10), 669 => to_unsigned(774, 10), 670 => to_unsigned(339, 10), 671 => to_unsigned(579, 10), 672 => to_unsigned(220, 10), 673 => to_unsigned(479, 10), 674 => to_unsigned(387, 10), 675 => to_unsigned(677, 10), 676 => to_unsigned(101, 10), 677 => to_unsigned(583, 10), 678 => to_unsigned(200, 10), 679 => to_unsigned(241, 10), 680 => to_unsigned(300, 10), 681 => to_unsigned(880, 10), 682 => to_unsigned(260, 10), 683 => to_unsigned(709, 10), 684 => to_unsigned(907, 10), 685 => to_unsigned(659, 10), 686 => to_unsigned(800, 10), 687 => to_unsigned(1014, 10), 688 => to_unsigned(464, 10), 689 => to_unsigned(553, 10), 690 => to_unsigned(752, 10), 691 => to_unsigned(301, 10), 692 => to_unsigned(710, 10), 693 => to_unsigned(470, 10), 694 => to_unsigned(354, 10), 695 => to_unsigned(321, 10), 696 => to_unsigned(762, 10), 697 => to_unsigned(30, 10), 698 => to_unsigned(815, 10), 699 => to_unsigned(636, 10), 700 => to_unsigned(117, 10), 701 => to_unsigned(353, 10), 702 => to_unsigned(193, 10), 703 => to_unsigned(417, 10), 704 => to_unsigned(234, 10), 705 => to_unsigned(65, 10), 706 => to_unsigned(509, 10), 707 => to_unsigned(942, 10), 708 => to_unsigned(530, 10), 709 => to_unsigned(185, 10), 710 => to_unsigned(717, 10), 711 => to_unsigned(23, 10), 712 => to_unsigned(63, 10), 713 => to_unsigned(528, 10), 714 => to_unsigned(7, 10), 715 => to_unsigned(354, 10), 716 => to_unsigned(1002, 10), 717 => to_unsigned(362, 10), 718 => to_unsigned(802, 10), 719 => to_unsigned(674, 10), 720 => to_unsigned(772, 10), 721 => to_unsigned(604, 10), 722 => to_unsigned(701, 10), 723 => to_unsigned(1003, 10), 724 => to_unsigned(552, 10), 725 => to_unsigned(367, 10), 726 => to_unsigned(80, 10), 727 => to_unsigned(122, 10), 728 => to_unsigned(20, 10), 729 => to_unsigned(585, 10), 730 => to_unsigned(827, 10), 731 => to_unsigned(549, 10), 732 => to_unsigned(291, 10), 733 => to_unsigned(253, 10), 734 => to_unsigned(862, 10), 735 => to_unsigned(505, 10), 736 => to_unsigned(293, 10), 737 => to_unsigned(508, 10), 738 => to_unsigned(690, 10), 739 => to_unsigned(37, 10), 740 => to_unsigned(913, 10), 741 => to_unsigned(623, 10), 742 => to_unsigned(690, 10), 743 => to_unsigned(742, 10), 744 => to_unsigned(176, 10), 745 => to_unsigned(441, 10), 746 => to_unsigned(565, 10), 747 => to_unsigned(291, 10), 748 => to_unsigned(561, 10), 749 => to_unsigned(270, 10), 750 => to_unsigned(40, 10), 751 => to_unsigned(133, 10), 752 => to_unsigned(934, 10), 753 => to_unsigned(92, 10), 754 => to_unsigned(90, 10), 755 => to_unsigned(65, 10), 756 => to_unsigned(955, 10), 757 => to_unsigned(742, 10), 758 => to_unsigned(629, 10), 759 => to_unsigned(345, 10), 760 => to_unsigned(724, 10), 761 => to_unsigned(778, 10), 762 => to_unsigned(581, 10), 763 => to_unsigned(62, 10), 764 => to_unsigned(102, 10), 765 => to_unsigned(824, 10), 766 => to_unsigned(65, 10), 767 => to_unsigned(112, 10), 768 => to_unsigned(187, 10), 769 => to_unsigned(618, 10), 770 => to_unsigned(813, 10), 771 => to_unsigned(260, 10), 772 => to_unsigned(418, 10), 773 => to_unsigned(35, 10), 774 => to_unsigned(560, 10), 775 => to_unsigned(591, 10), 776 => to_unsigned(681, 10), 777 => to_unsigned(488, 10), 778 => to_unsigned(944, 10), 779 => to_unsigned(195, 10), 780 => to_unsigned(371, 10), 781 => to_unsigned(972, 10), 782 => to_unsigned(326, 10), 783 => to_unsigned(892, 10), 784 => to_unsigned(83, 10), 785 => to_unsigned(1014, 10), 786 => to_unsigned(322, 10), 787 => to_unsigned(384, 10), 788 => to_unsigned(585, 10), 789 => to_unsigned(81, 10), 790 => to_unsigned(533, 10), 791 => to_unsigned(327, 10), 792 => to_unsigned(689, 10), 793 => to_unsigned(395, 10), 794 => to_unsigned(84, 10), 795 => to_unsigned(1016, 10), 796 => to_unsigned(1010, 10), 797 => to_unsigned(395, 10), 798 => to_unsigned(463, 10), 799 => to_unsigned(190, 10), 800 => to_unsigned(983, 10), 801 => to_unsigned(831, 10), 802 => to_unsigned(847, 10), 803 => to_unsigned(374, 10), 804 => to_unsigned(531, 10), 805 => to_unsigned(614, 10), 806 => to_unsigned(19, 10), 807 => to_unsigned(545, 10), 808 => to_unsigned(111, 10), 809 => to_unsigned(639, 10), 810 => to_unsigned(660, 10), 811 => to_unsigned(981, 10), 812 => to_unsigned(463, 10), 813 => to_unsigned(109, 10), 814 => to_unsigned(938, 10), 815 => to_unsigned(135, 10), 816 => to_unsigned(802, 10), 817 => to_unsigned(653, 10), 818 => to_unsigned(111, 10), 819 => to_unsigned(111, 10), 820 => to_unsigned(151, 10), 821 => to_unsigned(486, 10), 822 => to_unsigned(603, 10), 823 => to_unsigned(803, 10), 824 => to_unsigned(945, 10), 825 => to_unsigned(582, 10), 826 => to_unsigned(382, 10), 827 => to_unsigned(114, 10), 828 => to_unsigned(216, 10), 829 => to_unsigned(847, 10), 830 => to_unsigned(964, 10), 831 => to_unsigned(902, 10), 832 => to_unsigned(839, 10), 833 => to_unsigned(449, 10), 834 => to_unsigned(725, 10), 835 => to_unsigned(580, 10), 836 => to_unsigned(868, 10), 837 => to_unsigned(716, 10), 838 => to_unsigned(299, 10), 839 => to_unsigned(559, 10), 840 => to_unsigned(308, 10), 841 => to_unsigned(670, 10), 842 => to_unsigned(75, 10), 843 => to_unsigned(150, 10), 844 => to_unsigned(899, 10), 845 => to_unsigned(1015, 10), 846 => to_unsigned(989, 10), 847 => to_unsigned(492, 10), 848 => to_unsigned(131, 10), 849 => to_unsigned(945, 10), 850 => to_unsigned(662, 10), 851 => to_unsigned(66, 10), 852 => to_unsigned(549, 10), 853 => to_unsigned(658, 10), 854 => to_unsigned(891, 10), 855 => to_unsigned(184, 10), 856 => to_unsigned(981, 10), 857 => to_unsigned(699, 10), 858 => to_unsigned(835, 10), 859 => to_unsigned(39, 10), 860 => to_unsigned(388, 10), 861 => to_unsigned(844, 10), 862 => to_unsigned(308, 10), 863 => to_unsigned(817, 10), 864 => to_unsigned(864, 10), 865 => to_unsigned(594, 10), 866 => to_unsigned(376, 10), 867 => to_unsigned(187, 10), 868 => to_unsigned(675, 10), 869 => to_unsigned(582, 10), 870 => to_unsigned(860, 10), 871 => to_unsigned(599, 10), 872 => to_unsigned(408, 10), 873 => to_unsigned(603, 10), 874 => to_unsigned(146, 10), 875 => to_unsigned(656, 10), 876 => to_unsigned(377, 10), 877 => to_unsigned(420, 10), 878 => to_unsigned(560, 10), 879 => to_unsigned(745, 10), 880 => to_unsigned(432, 10), 881 => to_unsigned(959, 10), 882 => to_unsigned(385, 10), 883 => to_unsigned(692, 10), 884 => to_unsigned(270, 10), 885 => to_unsigned(27, 10), 886 => to_unsigned(13, 10), 887 => to_unsigned(118, 10), 888 => to_unsigned(690, 10), 889 => to_unsigned(845, 10), 890 => to_unsigned(236, 10), 891 => to_unsigned(794, 10), 892 => to_unsigned(916, 10), 893 => to_unsigned(762, 10), 894 => to_unsigned(910, 10), 895 => to_unsigned(723, 10), 896 => to_unsigned(999, 10), 897 => to_unsigned(218, 10), 898 => to_unsigned(657, 10), 899 => to_unsigned(85, 10), 900 => to_unsigned(928, 10), 901 => to_unsigned(344, 10), 902 => to_unsigned(102, 10), 903 => to_unsigned(711, 10), 904 => to_unsigned(731, 10), 905 => to_unsigned(584, 10), 906 => to_unsigned(558, 10), 907 => to_unsigned(86, 10), 908 => to_unsigned(269, 10), 909 => to_unsigned(621, 10), 910 => to_unsigned(687, 10), 911 => to_unsigned(286, 10), 912 => to_unsigned(898, 10), 913 => to_unsigned(495, 10), 914 => to_unsigned(537, 10), 915 => to_unsigned(872, 10), 916 => to_unsigned(1019, 10), 917 => to_unsigned(487, 10), 918 => to_unsigned(237, 10), 919 => to_unsigned(884, 10), 920 => to_unsigned(635, 10), 921 => to_unsigned(77, 10), 922 => to_unsigned(478, 10), 923 => to_unsigned(551, 10), 924 => to_unsigned(606, 10), 925 => to_unsigned(685, 10), 926 => to_unsigned(832, 10), 927 => to_unsigned(291, 10), 928 => to_unsigned(46, 10), 929 => to_unsigned(643, 10), 930 => to_unsigned(685, 10), 931 => to_unsigned(845, 10), 932 => to_unsigned(892, 10), 933 => to_unsigned(265, 10), 934 => to_unsigned(23, 10), 935 => to_unsigned(712, 10), 936 => to_unsigned(45, 10), 937 => to_unsigned(623, 10), 938 => to_unsigned(442, 10), 939 => to_unsigned(528, 10), 940 => to_unsigned(444, 10), 941 => to_unsigned(549, 10), 942 => to_unsigned(870, 10), 943 => to_unsigned(45, 10), 944 => to_unsigned(373, 10), 945 => to_unsigned(249, 10), 946 => to_unsigned(930, 10), 947 => to_unsigned(748, 10), 948 => to_unsigned(775, 10), 949 => to_unsigned(378, 10), 950 => to_unsigned(479, 10), 951 => to_unsigned(326, 10), 952 => to_unsigned(875, 10), 953 => to_unsigned(585, 10), 954 => to_unsigned(283, 10), 955 => to_unsigned(970, 10), 956 => to_unsigned(263, 10), 957 => to_unsigned(1003, 10), 958 => to_unsigned(856, 10), 959 => to_unsigned(399, 10), 960 => to_unsigned(764, 10), 961 => to_unsigned(543, 10), 962 => to_unsigned(483, 10), 963 => to_unsigned(227, 10), 964 => to_unsigned(702, 10), 965 => to_unsigned(742, 10), 966 => to_unsigned(345, 10), 967 => to_unsigned(585, 10), 968 => to_unsigned(174, 10), 969 => to_unsigned(679, 10), 970 => to_unsigned(251, 10), 971 => to_unsigned(319, 10), 972 => to_unsigned(30, 10), 973 => to_unsigned(29, 10), 974 => to_unsigned(915, 10), 975 => to_unsigned(161, 10), 976 => to_unsigned(590, 10), 977 => to_unsigned(967, 10), 978 => to_unsigned(613, 10), 979 => to_unsigned(272, 10), 980 => to_unsigned(233, 10), 981 => to_unsigned(126, 10), 982 => to_unsigned(886, 10), 983 => to_unsigned(508, 10), 984 => to_unsigned(75, 10), 985 => to_unsigned(730, 10), 986 => to_unsigned(28, 10), 987 => to_unsigned(134, 10), 988 => to_unsigned(407, 10), 989 => to_unsigned(209, 10), 990 => to_unsigned(732, 10), 991 => to_unsigned(959, 10), 992 => to_unsigned(878, 10), 993 => to_unsigned(168, 10), 994 => to_unsigned(291, 10), 995 => to_unsigned(92, 10), 996 => to_unsigned(563, 10), 997 => to_unsigned(401, 10), 998 => to_unsigned(690, 10), 999 => to_unsigned(690, 10), 1000 => to_unsigned(925, 10), 1001 => to_unsigned(844, 10), 1002 => to_unsigned(1021, 10), 1003 => to_unsigned(597, 10), 1004 => to_unsigned(238, 10), 1005 => to_unsigned(517, 10), 1006 => to_unsigned(810, 10), 1007 => to_unsigned(644, 10), 1008 => to_unsigned(170, 10), 1009 => to_unsigned(761, 10), 1010 => to_unsigned(280, 10), 1011 => to_unsigned(263, 10), 1012 => to_unsigned(665, 10), 1013 => to_unsigned(935, 10), 1014 => to_unsigned(78, 10), 1015 => to_unsigned(556, 10), 1016 => to_unsigned(145, 10), 1017 => to_unsigned(835, 10), 1018 => to_unsigned(669, 10), 1019 => to_unsigned(54, 10), 1020 => to_unsigned(301, 10), 1021 => to_unsigned(739, 10), 1022 => to_unsigned(865, 10), 1023 => to_unsigned(572, 10), 1024 => to_unsigned(767, 10), 1025 => to_unsigned(852, 10), 1026 => to_unsigned(150, 10), 1027 => to_unsigned(690, 10), 1028 => to_unsigned(302, 10), 1029 => to_unsigned(474, 10), 1030 => to_unsigned(952, 10), 1031 => to_unsigned(642, 10), 1032 => to_unsigned(1003, 10), 1033 => to_unsigned(107, 10), 1034 => to_unsigned(428, 10), 1035 => to_unsigned(302, 10), 1036 => to_unsigned(18, 10), 1037 => to_unsigned(2, 10), 1038 => to_unsigned(1008, 10), 1039 => to_unsigned(769, 10), 1040 => to_unsigned(58, 10), 1041 => to_unsigned(850, 10), 1042 => to_unsigned(192, 10), 1043 => to_unsigned(881, 10), 1044 => to_unsigned(271, 10), 1045 => to_unsigned(782, 10), 1046 => to_unsigned(849, 10), 1047 => to_unsigned(234, 10), 1048 => to_unsigned(818, 10), 1049 => to_unsigned(956, 10), 1050 => to_unsigned(301, 10), 1051 => to_unsigned(266, 10), 1052 => to_unsigned(464, 10), 1053 => to_unsigned(236, 10), 1054 => to_unsigned(746, 10), 1055 => to_unsigned(964, 10), 1056 => to_unsigned(872, 10), 1057 => to_unsigned(778, 10), 1058 => to_unsigned(996, 10), 1059 => to_unsigned(694, 10), 1060 => to_unsigned(630, 10), 1061 => to_unsigned(951, 10), 1062 => to_unsigned(436, 10), 1063 => to_unsigned(986, 10), 1064 => to_unsigned(750, 10), 1065 => to_unsigned(715, 10), 1066 => to_unsigned(304, 10), 1067 => to_unsigned(950, 10), 1068 => to_unsigned(288, 10), 1069 => to_unsigned(75, 10), 1070 => to_unsigned(556, 10), 1071 => to_unsigned(895, 10), 1072 => to_unsigned(897, 10), 1073 => to_unsigned(200, 10), 1074 => to_unsigned(326, 10), 1075 => to_unsigned(446, 10), 1076 => to_unsigned(291, 10), 1077 => to_unsigned(589, 10), 1078 => to_unsigned(668, 10), 1079 => to_unsigned(874, 10), 1080 => to_unsigned(217, 10), 1081 => to_unsigned(703, 10), 1082 => to_unsigned(539, 10), 1083 => to_unsigned(722, 10), 1084 => to_unsigned(894, 10), 1085 => to_unsigned(22, 10), 1086 => to_unsigned(874, 10), 1087 => to_unsigned(138, 10), 1088 => to_unsigned(569, 10), 1089 => to_unsigned(151, 10), 1090 => to_unsigned(107, 10), 1091 => to_unsigned(825, 10), 1092 => to_unsigned(286, 10), 1093 => to_unsigned(46, 10), 1094 => to_unsigned(643, 10), 1095 => to_unsigned(262, 10), 1096 => to_unsigned(899, 10), 1097 => to_unsigned(740, 10), 1098 => to_unsigned(208, 10), 1099 => to_unsigned(80, 10), 1100 => to_unsigned(35, 10), 1101 => to_unsigned(889, 10), 1102 => to_unsigned(252, 10), 1103 => to_unsigned(210, 10), 1104 => to_unsigned(298, 10), 1105 => to_unsigned(103, 10), 1106 => to_unsigned(255, 10), 1107 => to_unsigned(361, 10), 1108 => to_unsigned(111, 10), 1109 => to_unsigned(490, 10), 1110 => to_unsigned(602, 10), 1111 => to_unsigned(726, 10), 1112 => to_unsigned(991, 10), 1113 => to_unsigned(638, 10), 1114 => to_unsigned(100, 10), 1115 => to_unsigned(172, 10), 1116 => to_unsigned(910, 10), 1117 => to_unsigned(869, 10), 1118 => to_unsigned(269, 10), 1119 => to_unsigned(190, 10), 1120 => to_unsigned(155, 10), 1121 => to_unsigned(923, 10), 1122 => to_unsigned(1008, 10), 1123 => to_unsigned(503, 10), 1124 => to_unsigned(879, 10), 1125 => to_unsigned(725, 10), 1126 => to_unsigned(1023, 10), 1127 => to_unsigned(433, 10), 1128 => to_unsigned(29, 10), 1129 => to_unsigned(749, 10), 1130 => to_unsigned(946, 10), 1131 => to_unsigned(458, 10), 1132 => to_unsigned(689, 10), 1133 => to_unsigned(298, 10), 1134 => to_unsigned(305, 10), 1135 => to_unsigned(874, 10), 1136 => to_unsigned(225, 10), 1137 => to_unsigned(228, 10), 1138 => to_unsigned(97, 10), 1139 => to_unsigned(407, 10), 1140 => to_unsigned(951, 10), 1141 => to_unsigned(714, 10), 1142 => to_unsigned(759, 10), 1143 => to_unsigned(342, 10), 1144 => to_unsigned(157, 10), 1145 => to_unsigned(642, 10), 1146 => to_unsigned(252, 10), 1147 => to_unsigned(995, 10), 1148 => to_unsigned(1022, 10), 1149 => to_unsigned(792, 10), 1150 => to_unsigned(649, 10), 1151 => to_unsigned(738, 10), 1152 => to_unsigned(672, 10), 1153 => to_unsigned(233, 10), 1154 => to_unsigned(689, 10), 1155 => to_unsigned(215, 10), 1156 => to_unsigned(254, 10), 1157 => to_unsigned(927, 10), 1158 => to_unsigned(320, 10), 1159 => to_unsigned(698, 10), 1160 => to_unsigned(453, 10), 1161 => to_unsigned(145, 10), 1162 => to_unsigned(828, 10), 1163 => to_unsigned(767, 10), 1164 => to_unsigned(511, 10), 1165 => to_unsigned(355, 10), 1166 => to_unsigned(878, 10), 1167 => to_unsigned(372, 10), 1168 => to_unsigned(692, 10), 1169 => to_unsigned(898, 10), 1170 => to_unsigned(28, 10), 1171 => to_unsigned(255, 10), 1172 => to_unsigned(178, 10), 1173 => to_unsigned(555, 10), 1174 => to_unsigned(910, 10), 1175 => to_unsigned(80, 10), 1176 => to_unsigned(476, 10), 1177 => to_unsigned(328, 10), 1178 => to_unsigned(815, 10), 1179 => to_unsigned(191, 10), 1180 => to_unsigned(761, 10), 1181 => to_unsigned(199, 10), 1182 => to_unsigned(241, 10), 1183 => to_unsigned(370, 10), 1184 => to_unsigned(476, 10), 1185 => to_unsigned(279, 10), 1186 => to_unsigned(776, 10), 1187 => to_unsigned(972, 10), 1188 => to_unsigned(309, 10), 1189 => to_unsigned(276, 10), 1190 => to_unsigned(634, 10), 1191 => to_unsigned(629, 10), 1192 => to_unsigned(729, 10), 1193 => to_unsigned(670, 10), 1194 => to_unsigned(95, 10), 1195 => to_unsigned(661, 10), 1196 => to_unsigned(158, 10), 1197 => to_unsigned(963, 10), 1198 => to_unsigned(406, 10), 1199 => to_unsigned(653, 10), 1200 => to_unsigned(1008, 10), 1201 => to_unsigned(619, 10), 1202 => to_unsigned(759, 10), 1203 => to_unsigned(450, 10), 1204 => to_unsigned(796, 10), 1205 => to_unsigned(180, 10), 1206 => to_unsigned(93, 10), 1207 => to_unsigned(34, 10), 1208 => to_unsigned(665, 10), 1209 => to_unsigned(341, 10), 1210 => to_unsigned(693, 10), 1211 => to_unsigned(71, 10), 1212 => to_unsigned(514, 10), 1213 => to_unsigned(111, 10), 1214 => to_unsigned(848, 10), 1215 => to_unsigned(272, 10), 1216 => to_unsigned(493, 10), 1217 => to_unsigned(542, 10), 1218 => to_unsigned(35, 10), 1219 => to_unsigned(129, 10), 1220 => to_unsigned(681, 10), 1221 => to_unsigned(90, 10), 1222 => to_unsigned(688, 10), 1223 => to_unsigned(953, 10), 1224 => to_unsigned(376, 10), 1225 => to_unsigned(42, 10), 1226 => to_unsigned(298, 10), 1227 => to_unsigned(398, 10), 1228 => to_unsigned(120, 10), 1229 => to_unsigned(192, 10), 1230 => to_unsigned(941, 10), 1231 => to_unsigned(487, 10), 1232 => to_unsigned(300, 10), 1233 => to_unsigned(693, 10), 1234 => to_unsigned(283, 10), 1235 => to_unsigned(525, 10), 1236 => to_unsigned(161, 10), 1237 => to_unsigned(63, 10), 1238 => to_unsigned(215, 10), 1239 => to_unsigned(95, 10), 1240 => to_unsigned(37, 10), 1241 => to_unsigned(274, 10), 1242 => to_unsigned(975, 10), 1243 => to_unsigned(858, 10), 1244 => to_unsigned(889, 10), 1245 => to_unsigned(579, 10), 1246 => to_unsigned(7, 10), 1247 => to_unsigned(181, 10), 1248 => to_unsigned(507, 10), 1249 => to_unsigned(139, 10), 1250 => to_unsigned(481, 10), 1251 => to_unsigned(136, 10), 1252 => to_unsigned(452, 10), 1253 => to_unsigned(44, 10), 1254 => to_unsigned(536, 10), 1255 => to_unsigned(970, 10), 1256 => to_unsigned(540, 10), 1257 => to_unsigned(52, 10), 1258 => to_unsigned(736, 10), 1259 => to_unsigned(526, 10), 1260 => to_unsigned(811, 10), 1261 => to_unsigned(712, 10), 1262 => to_unsigned(777, 10), 1263 => to_unsigned(434, 10), 1264 => to_unsigned(366, 10), 1265 => to_unsigned(995, 10), 1266 => to_unsigned(514, 10), 1267 => to_unsigned(959, 10), 1268 => to_unsigned(106, 10), 1269 => to_unsigned(861, 10), 1270 => to_unsigned(232, 10), 1271 => to_unsigned(157, 10), 1272 => to_unsigned(632, 10), 1273 => to_unsigned(585, 10), 1274 => to_unsigned(864, 10), 1275 => to_unsigned(965, 10), 1276 => to_unsigned(868, 10), 1277 => to_unsigned(921, 10), 1278 => to_unsigned(42, 10), 1279 => to_unsigned(482, 10), 1280 => to_unsigned(385, 10), 1281 => to_unsigned(251, 10), 1282 => to_unsigned(827, 10), 1283 => to_unsigned(105, 10), 1284 => to_unsigned(334, 10), 1285 => to_unsigned(128, 10), 1286 => to_unsigned(783, 10), 1287 => to_unsigned(969, 10), 1288 => to_unsigned(119, 10), 1289 => to_unsigned(736, 10), 1290 => to_unsigned(397, 10), 1291 => to_unsigned(848, 10), 1292 => to_unsigned(579, 10), 1293 => to_unsigned(102, 10), 1294 => to_unsigned(437, 10), 1295 => to_unsigned(779, 10), 1296 => to_unsigned(749, 10), 1297 => to_unsigned(336, 10), 1298 => to_unsigned(441, 10), 1299 => to_unsigned(462, 10), 1300 => to_unsigned(625, 10), 1301 => to_unsigned(100, 10), 1302 => to_unsigned(190, 10), 1303 => to_unsigned(997, 10), 1304 => to_unsigned(27, 10), 1305 => to_unsigned(705, 10), 1306 => to_unsigned(194, 10), 1307 => to_unsigned(449, 10), 1308 => to_unsigned(641, 10), 1309 => to_unsigned(932, 10), 1310 => to_unsigned(228, 10), 1311 => to_unsigned(418, 10), 1312 => to_unsigned(453, 10), 1313 => to_unsigned(613, 10), 1314 => to_unsigned(739, 10), 1315 => to_unsigned(206, 10), 1316 => to_unsigned(1016, 10), 1317 => to_unsigned(266, 10), 1318 => to_unsigned(116, 10), 1319 => to_unsigned(584, 10), 1320 => to_unsigned(531, 10), 1321 => to_unsigned(534, 10), 1322 => to_unsigned(330, 10), 1323 => to_unsigned(592, 10), 1324 => to_unsigned(989, 10), 1325 => to_unsigned(443, 10), 1326 => to_unsigned(822, 10), 1327 => to_unsigned(632, 10), 1328 => to_unsigned(687, 10), 1329 => to_unsigned(967, 10), 1330 => to_unsigned(669, 10), 1331 => to_unsigned(712, 10), 1332 => to_unsigned(602, 10), 1333 => to_unsigned(734, 10), 1334 => to_unsigned(960, 10), 1335 => to_unsigned(716, 10), 1336 => to_unsigned(453, 10), 1337 => to_unsigned(758, 10), 1338 => to_unsigned(240, 10), 1339 => to_unsigned(598, 10), 1340 => to_unsigned(490, 10), 1341 => to_unsigned(425, 10), 1342 => to_unsigned(354, 10), 1343 => to_unsigned(871, 10), 1344 => to_unsigned(473, 10), 1345 => to_unsigned(314, 10), 1346 => to_unsigned(460, 10), 1347 => to_unsigned(619, 10), 1348 => to_unsigned(82, 10), 1349 => to_unsigned(299, 10), 1350 => to_unsigned(300, 10), 1351 => to_unsigned(467, 10), 1352 => to_unsigned(373, 10), 1353 => to_unsigned(474, 10), 1354 => to_unsigned(598, 10), 1355 => to_unsigned(715, 10), 1356 => to_unsigned(61, 10), 1357 => to_unsigned(765, 10), 1358 => to_unsigned(632, 10), 1359 => to_unsigned(856, 10), 1360 => to_unsigned(903, 10), 1361 => to_unsigned(534, 10), 1362 => to_unsigned(298, 10), 1363 => to_unsigned(332, 10), 1364 => to_unsigned(757, 10), 1365 => to_unsigned(164, 10), 1366 => to_unsigned(97, 10), 1367 => to_unsigned(362, 10), 1368 => to_unsigned(939, 10), 1369 => to_unsigned(828, 10), 1370 => to_unsigned(578, 10), 1371 => to_unsigned(456, 10), 1372 => to_unsigned(738, 10), 1373 => to_unsigned(124, 10), 1374 => to_unsigned(893, 10), 1375 => to_unsigned(447, 10), 1376 => to_unsigned(223, 10), 1377 => to_unsigned(44, 10), 1378 => to_unsigned(225, 10), 1379 => to_unsigned(11, 10), 1380 => to_unsigned(314, 10), 1381 => to_unsigned(196, 10), 1382 => to_unsigned(825, 10), 1383 => to_unsigned(917, 10), 1384 => to_unsigned(949, 10), 1385 => to_unsigned(262, 10), 1386 => to_unsigned(615, 10), 1387 => to_unsigned(25, 10), 1388 => to_unsigned(803, 10), 1389 => to_unsigned(276, 10), 1390 => to_unsigned(563, 10), 1391 => to_unsigned(631, 10), 1392 => to_unsigned(522, 10), 1393 => to_unsigned(469, 10), 1394 => to_unsigned(541, 10), 1395 => to_unsigned(800, 10), 1396 => to_unsigned(505, 10), 1397 => to_unsigned(482, 10), 1398 => to_unsigned(388, 10), 1399 => to_unsigned(242, 10), 1400 => to_unsigned(596, 10), 1401 => to_unsigned(286, 10), 1402 => to_unsigned(942, 10), 1403 => to_unsigned(14, 10), 1404 => to_unsigned(380, 10), 1405 => to_unsigned(987, 10), 1406 => to_unsigned(822, 10), 1407 => to_unsigned(485, 10), 1408 => to_unsigned(307, 10), 1409 => to_unsigned(461, 10), 1410 => to_unsigned(594, 10), 1411 => to_unsigned(350, 10), 1412 => to_unsigned(124, 10), 1413 => to_unsigned(33, 10), 1414 => to_unsigned(125, 10), 1415 => to_unsigned(719, 10), 1416 => to_unsigned(997, 10), 1417 => to_unsigned(426, 10), 1418 => to_unsigned(53, 10), 1419 => to_unsigned(432, 10), 1420 => to_unsigned(772, 10), 1421 => to_unsigned(958, 10), 1422 => to_unsigned(918, 10), 1423 => to_unsigned(973, 10), 1424 => to_unsigned(455, 10), 1425 => to_unsigned(330, 10), 1426 => to_unsigned(491, 10), 1427 => to_unsigned(304, 10), 1428 => to_unsigned(320, 10), 1429 => to_unsigned(963, 10), 1430 => to_unsigned(855, 10), 1431 => to_unsigned(268, 10), 1432 => to_unsigned(305, 10), 1433 => to_unsigned(672, 10), 1434 => to_unsigned(338, 10), 1435 => to_unsigned(759, 10), 1436 => to_unsigned(824, 10), 1437 => to_unsigned(717, 10), 1438 => to_unsigned(721, 10), 1439 => to_unsigned(25, 10), 1440 => to_unsigned(287, 10), 1441 => to_unsigned(798, 10), 1442 => to_unsigned(280, 10), 1443 => to_unsigned(630, 10), 1444 => to_unsigned(367, 10), 1445 => to_unsigned(509, 10), 1446 => to_unsigned(560, 10), 1447 => to_unsigned(904, 10), 1448 => to_unsigned(724, 10), 1449 => to_unsigned(303, 10), 1450 => to_unsigned(886, 10), 1451 => to_unsigned(1, 10), 1452 => to_unsigned(459, 10), 1453 => to_unsigned(250, 10), 1454 => to_unsigned(865, 10), 1455 => to_unsigned(138, 10), 1456 => to_unsigned(378, 10), 1457 => to_unsigned(803, 10), 1458 => to_unsigned(555, 10), 1459 => to_unsigned(874, 10), 1460 => to_unsigned(391, 10), 1461 => to_unsigned(894, 10), 1462 => to_unsigned(325, 10), 1463 => to_unsigned(270, 10), 1464 => to_unsigned(664, 10), 1465 => to_unsigned(788, 10), 1466 => to_unsigned(554, 10), 1467 => to_unsigned(901, 10), 1468 => to_unsigned(175, 10), 1469 => to_unsigned(573, 10), 1470 => to_unsigned(419, 10), 1471 => to_unsigned(463, 10), 1472 => to_unsigned(192, 10), 1473 => to_unsigned(15, 10), 1474 => to_unsigned(198, 10), 1475 => to_unsigned(606, 10), 1476 => to_unsigned(630, 10), 1477 => to_unsigned(118, 10), 1478 => to_unsigned(13, 10), 1479 => to_unsigned(483, 10), 1480 => to_unsigned(8, 10), 1481 => to_unsigned(564, 10), 1482 => to_unsigned(479, 10), 1483 => to_unsigned(228, 10), 1484 => to_unsigned(933, 10), 1485 => to_unsigned(28, 10), 1486 => to_unsigned(717, 10), 1487 => to_unsigned(753, 10), 1488 => to_unsigned(1009, 10), 1489 => to_unsigned(461, 10), 1490 => to_unsigned(349, 10), 1491 => to_unsigned(655, 10), 1492 => to_unsigned(622, 10), 1493 => to_unsigned(491, 10), 1494 => to_unsigned(412, 10), 1495 => to_unsigned(145, 10), 1496 => to_unsigned(676, 10), 1497 => to_unsigned(16, 10), 1498 => to_unsigned(379, 10), 1499 => to_unsigned(757, 10), 1500 => to_unsigned(434, 10), 1501 => to_unsigned(900, 10), 1502 => to_unsigned(107, 10), 1503 => to_unsigned(204, 10), 1504 => to_unsigned(719, 10), 1505 => to_unsigned(650, 10), 1506 => to_unsigned(543, 10), 1507 => to_unsigned(1006, 10), 1508 => to_unsigned(11, 10), 1509 => to_unsigned(860, 10), 1510 => to_unsigned(154, 10), 1511 => to_unsigned(851, 10), 1512 => to_unsigned(3, 10), 1513 => to_unsigned(101, 10), 1514 => to_unsigned(579, 10), 1515 => to_unsigned(872, 10), 1516 => to_unsigned(846, 10), 1517 => to_unsigned(213, 10), 1518 => to_unsigned(526, 10), 1519 => to_unsigned(424, 10), 1520 => to_unsigned(24, 10), 1521 => to_unsigned(388, 10), 1522 => to_unsigned(201, 10), 1523 => to_unsigned(251, 10), 1524 => to_unsigned(404, 10), 1525 => to_unsigned(23, 10), 1526 => to_unsigned(114, 10), 1527 => to_unsigned(1017, 10), 1528 => to_unsigned(368, 10), 1529 => to_unsigned(685, 10), 1530 => to_unsigned(242, 10), 1531 => to_unsigned(519, 10), 1532 => to_unsigned(280, 10), 1533 => to_unsigned(221, 10), 1534 => to_unsigned(258, 10), 1535 => to_unsigned(372, 10), 1536 => to_unsigned(1010, 10), 1537 => to_unsigned(297, 10), 1538 => to_unsigned(711, 10), 1539 => to_unsigned(50, 10), 1540 => to_unsigned(775, 10), 1541 => to_unsigned(4, 10), 1542 => to_unsigned(31, 10), 1543 => to_unsigned(247, 10), 1544 => to_unsigned(687, 10), 1545 => to_unsigned(667, 10), 1546 => to_unsigned(11, 10), 1547 => to_unsigned(71, 10), 1548 => to_unsigned(1, 10), 1549 => to_unsigned(173, 10), 1550 => to_unsigned(823, 10), 1551 => to_unsigned(854, 10), 1552 => to_unsigned(533, 10), 1553 => to_unsigned(542, 10), 1554 => to_unsigned(117, 10), 1555 => to_unsigned(616, 10), 1556 => to_unsigned(27, 10), 1557 => to_unsigned(156, 10), 1558 => to_unsigned(956, 10), 1559 => to_unsigned(47, 10), 1560 => to_unsigned(596, 10), 1561 => to_unsigned(449, 10), 1562 => to_unsigned(948, 10), 1563 => to_unsigned(479, 10), 1564 => to_unsigned(77, 10), 1565 => to_unsigned(1005, 10), 1566 => to_unsigned(325, 10), 1567 => to_unsigned(433, 10), 1568 => to_unsigned(810, 10), 1569 => to_unsigned(824, 10), 1570 => to_unsigned(266, 10), 1571 => to_unsigned(778, 10), 1572 => to_unsigned(177, 10), 1573 => to_unsigned(440, 10), 1574 => to_unsigned(42, 10), 1575 => to_unsigned(893, 10), 1576 => to_unsigned(424, 10), 1577 => to_unsigned(718, 10), 1578 => to_unsigned(736, 10), 1579 => to_unsigned(307, 10), 1580 => to_unsigned(1009, 10), 1581 => to_unsigned(772, 10), 1582 => to_unsigned(564, 10), 1583 => to_unsigned(858, 10), 1584 => to_unsigned(168, 10), 1585 => to_unsigned(278, 10), 1586 => to_unsigned(902, 10), 1587 => to_unsigned(944, 10), 1588 => to_unsigned(703, 10), 1589 => to_unsigned(454, 10), 1590 => to_unsigned(496, 10), 1591 => to_unsigned(248, 10), 1592 => to_unsigned(262, 10), 1593 => to_unsigned(877, 10), 1594 => to_unsigned(381, 10), 1595 => to_unsigned(39, 10), 1596 => to_unsigned(52, 10), 1597 => to_unsigned(496, 10), 1598 => to_unsigned(195, 10), 1599 => to_unsigned(502, 10), 1600 => to_unsigned(215, 10), 1601 => to_unsigned(1010, 10), 1602 => to_unsigned(322, 10), 1603 => to_unsigned(823, 10), 1604 => to_unsigned(773, 10), 1605 => to_unsigned(723, 10), 1606 => to_unsigned(261, 10), 1607 => to_unsigned(499, 10), 1608 => to_unsigned(843, 10), 1609 => to_unsigned(668, 10), 1610 => to_unsigned(86, 10), 1611 => to_unsigned(918, 10), 1612 => to_unsigned(761, 10), 1613 => to_unsigned(414, 10), 1614 => to_unsigned(232, 10), 1615 => to_unsigned(421, 10), 1616 => to_unsigned(630, 10), 1617 => to_unsigned(998, 10), 1618 => to_unsigned(878, 10), 1619 => to_unsigned(15, 10), 1620 => to_unsigned(280, 10), 1621 => to_unsigned(922, 10), 1622 => to_unsigned(357, 10), 1623 => to_unsigned(929, 10), 1624 => to_unsigned(917, 10), 1625 => to_unsigned(306, 10), 1626 => to_unsigned(582, 10), 1627 => to_unsigned(19, 10), 1628 => to_unsigned(265, 10), 1629 => to_unsigned(108, 10), 1630 => to_unsigned(212, 10), 1631 => to_unsigned(139, 10), 1632 => to_unsigned(283, 10), 1633 => to_unsigned(152, 10), 1634 => to_unsigned(106, 10), 1635 => to_unsigned(56, 10), 1636 => to_unsigned(719, 10), 1637 => to_unsigned(800, 10), 1638 => to_unsigned(124, 10), 1639 => to_unsigned(301, 10), 1640 => to_unsigned(367, 10), 1641 => to_unsigned(871, 10), 1642 => to_unsigned(596, 10), 1643 => to_unsigned(802, 10), 1644 => to_unsigned(451, 10), 1645 => to_unsigned(994, 10), 1646 => to_unsigned(994, 10), 1647 => to_unsigned(906, 10), 1648 => to_unsigned(200, 10), 1649 => to_unsigned(453, 10), 1650 => to_unsigned(403, 10), 1651 => to_unsigned(951, 10), 1652 => to_unsigned(706, 10), 1653 => to_unsigned(693, 10), 1654 => to_unsigned(823, 10), 1655 => to_unsigned(904, 10), 1656 => to_unsigned(507, 10), 1657 => to_unsigned(445, 10), 1658 => to_unsigned(59, 10), 1659 => to_unsigned(176, 10), 1660 => to_unsigned(172, 10), 1661 => to_unsigned(758, 10), 1662 => to_unsigned(301, 10), 1663 => to_unsigned(682, 10), 1664 => to_unsigned(561, 10), 1665 => to_unsigned(773, 10), 1666 => to_unsigned(222, 10), 1667 => to_unsigned(206, 10), 1668 => to_unsigned(524, 10), 1669 => to_unsigned(291, 10), 1670 => to_unsigned(713, 10), 1671 => to_unsigned(314, 10), 1672 => to_unsigned(432, 10), 1673 => to_unsigned(619, 10), 1674 => to_unsigned(235, 10), 1675 => to_unsigned(791, 10), 1676 => to_unsigned(701, 10), 1677 => to_unsigned(461, 10), 1678 => to_unsigned(460, 10), 1679 => to_unsigned(593, 10), 1680 => to_unsigned(584, 10), 1681 => to_unsigned(20, 10), 1682 => to_unsigned(209, 10), 1683 => to_unsigned(100, 10), 1684 => to_unsigned(985, 10), 1685 => to_unsigned(817, 10), 1686 => to_unsigned(373, 10), 1687 => to_unsigned(938, 10), 1688 => to_unsigned(266, 10), 1689 => to_unsigned(547, 10), 1690 => to_unsigned(577, 10), 1691 => to_unsigned(521, 10), 1692 => to_unsigned(174, 10), 1693 => to_unsigned(838, 10), 1694 => to_unsigned(270, 10), 1695 => to_unsigned(711, 10), 1696 => to_unsigned(854, 10), 1697 => to_unsigned(217, 10), 1698 => to_unsigned(133, 10), 1699 => to_unsigned(583, 10), 1700 => to_unsigned(730, 10), 1701 => to_unsigned(492, 10), 1702 => to_unsigned(513, 10), 1703 => to_unsigned(1012, 10), 1704 => to_unsigned(199, 10), 1705 => to_unsigned(165, 10), 1706 => to_unsigned(292, 10), 1707 => to_unsigned(650, 10), 1708 => to_unsigned(258, 10), 1709 => to_unsigned(363, 10), 1710 => to_unsigned(153, 10), 1711 => to_unsigned(879, 10), 1712 => to_unsigned(300, 10), 1713 => to_unsigned(222, 10), 1714 => to_unsigned(882, 10), 1715 => to_unsigned(583, 10), 1716 => to_unsigned(674, 10), 1717 => to_unsigned(700, 10), 1718 => to_unsigned(9, 10), 1719 => to_unsigned(998, 10), 1720 => to_unsigned(13, 10), 1721 => to_unsigned(549, 10), 1722 => to_unsigned(118, 10), 1723 => to_unsigned(949, 10), 1724 => to_unsigned(445, 10), 1725 => to_unsigned(853, 10), 1726 => to_unsigned(915, 10), 1727 => to_unsigned(122, 10), 1728 => to_unsigned(720, 10), 1729 => to_unsigned(235, 10), 1730 => to_unsigned(267, 10), 1731 => to_unsigned(89, 10), 1732 => to_unsigned(135, 10), 1733 => to_unsigned(354, 10), 1734 => to_unsigned(178, 10), 1735 => to_unsigned(538, 10), 1736 => to_unsigned(605, 10), 1737 => to_unsigned(969, 10), 1738 => to_unsigned(137, 10), 1739 => to_unsigned(182, 10), 1740 => to_unsigned(434, 10), 1741 => to_unsigned(10, 10), 1742 => to_unsigned(77, 10), 1743 => to_unsigned(754, 10), 1744 => to_unsigned(235, 10), 1745 => to_unsigned(238, 10), 1746 => to_unsigned(564, 10), 1747 => to_unsigned(180, 10), 1748 => to_unsigned(433, 10), 1749 => to_unsigned(727, 10), 1750 => to_unsigned(105, 10), 1751 => to_unsigned(732, 10), 1752 => to_unsigned(77, 10), 1753 => to_unsigned(342, 10), 1754 => to_unsigned(503, 10), 1755 => to_unsigned(750, 10), 1756 => to_unsigned(482, 10), 1757 => to_unsigned(874, 10), 1758 => to_unsigned(355, 10), 1759 => to_unsigned(87, 10), 1760 => to_unsigned(718, 10), 1761 => to_unsigned(919, 10), 1762 => to_unsigned(880, 10), 1763 => to_unsigned(37, 10), 1764 => to_unsigned(286, 10), 1765 => to_unsigned(174, 10), 1766 => to_unsigned(223, 10), 1767 => to_unsigned(931, 10), 1768 => to_unsigned(683, 10), 1769 => to_unsigned(647, 10), 1770 => to_unsigned(530, 10), 1771 => to_unsigned(799, 10), 1772 => to_unsigned(134, 10), 1773 => to_unsigned(335, 10), 1774 => to_unsigned(99, 10), 1775 => to_unsigned(441, 10), 1776 => to_unsigned(997, 10), 1777 => to_unsigned(383, 10), 1778 => to_unsigned(822, 10), 1779 => to_unsigned(272, 10), 1780 => to_unsigned(246, 10), 1781 => to_unsigned(701, 10), 1782 => to_unsigned(171, 10), 1783 => to_unsigned(193, 10), 1784 => to_unsigned(934, 10), 1785 => to_unsigned(713, 10), 1786 => to_unsigned(889, 10), 1787 => to_unsigned(67, 10), 1788 => to_unsigned(471, 10), 1789 => to_unsigned(581, 10), 1790 => to_unsigned(320, 10), 1791 => to_unsigned(838, 10), 1792 => to_unsigned(322, 10), 1793 => to_unsigned(199, 10), 1794 => to_unsigned(631, 10), 1795 => to_unsigned(1009, 10), 1796 => to_unsigned(791, 10), 1797 => to_unsigned(752, 10), 1798 => to_unsigned(352, 10), 1799 => to_unsigned(100, 10), 1800 => to_unsigned(575, 10), 1801 => to_unsigned(122, 10), 1802 => to_unsigned(807, 10), 1803 => to_unsigned(582, 10), 1804 => to_unsigned(776, 10), 1805 => to_unsigned(82, 10), 1806 => to_unsigned(248, 10), 1807 => to_unsigned(134, 10), 1808 => to_unsigned(32, 10), 1809 => to_unsigned(239, 10), 1810 => to_unsigned(819, 10), 1811 => to_unsigned(127, 10), 1812 => to_unsigned(14, 10), 1813 => to_unsigned(362, 10), 1814 => to_unsigned(287, 10), 1815 => to_unsigned(483, 10), 1816 => to_unsigned(1018, 10), 1817 => to_unsigned(729, 10), 1818 => to_unsigned(243, 10), 1819 => to_unsigned(908, 10), 1820 => to_unsigned(408, 10), 1821 => to_unsigned(52, 10), 1822 => to_unsigned(1007, 10), 1823 => to_unsigned(445, 10), 1824 => to_unsigned(306, 10), 1825 => to_unsigned(78, 10), 1826 => to_unsigned(393, 10), 1827 => to_unsigned(662, 10), 1828 => to_unsigned(332, 10), 1829 => to_unsigned(37, 10), 1830 => to_unsigned(97, 10), 1831 => to_unsigned(452, 10), 1832 => to_unsigned(382, 10), 1833 => to_unsigned(941, 10), 1834 => to_unsigned(814, 10), 1835 => to_unsigned(19, 10), 1836 => to_unsigned(40, 10), 1837 => to_unsigned(836, 10), 1838 => to_unsigned(650, 10), 1839 => to_unsigned(267, 10), 1840 => to_unsigned(628, 10), 1841 => to_unsigned(439, 10), 1842 => to_unsigned(395, 10), 1843 => to_unsigned(241, 10), 1844 => to_unsigned(257, 10), 1845 => to_unsigned(997, 10), 1846 => to_unsigned(836, 10), 1847 => to_unsigned(329, 10), 1848 => to_unsigned(878, 10), 1849 => to_unsigned(114, 10), 1850 => to_unsigned(91, 10), 1851 => to_unsigned(495, 10), 1852 => to_unsigned(735, 10), 1853 => to_unsigned(308, 10), 1854 => to_unsigned(302, 10), 1855 => to_unsigned(884, 10), 1856 => to_unsigned(852, 10), 1857 => to_unsigned(787, 10), 1858 => to_unsigned(421, 10), 1859 => to_unsigned(411, 10), 1860 => to_unsigned(822, 10), 1861 => to_unsigned(790, 10), 1862 => to_unsigned(543, 10), 1863 => to_unsigned(795, 10), 1864 => to_unsigned(898, 10), 1865 => to_unsigned(53, 10), 1866 => to_unsigned(625, 10), 1867 => to_unsigned(290, 10), 1868 => to_unsigned(592, 10), 1869 => to_unsigned(914, 10), 1870 => to_unsigned(169, 10), 1871 => to_unsigned(934, 10), 1872 => to_unsigned(707, 10), 1873 => to_unsigned(929, 10), 1874 => to_unsigned(583, 10), 1875 => to_unsigned(658, 10), 1876 => to_unsigned(755, 10), 1877 => to_unsigned(755, 10), 1878 => to_unsigned(326, 10), 1879 => to_unsigned(262, 10), 1880 => to_unsigned(302, 10), 1881 => to_unsigned(983, 10), 1882 => to_unsigned(216, 10), 1883 => to_unsigned(704, 10), 1884 => to_unsigned(100, 10), 1885 => to_unsigned(163, 10), 1886 => to_unsigned(898, 10), 1887 => to_unsigned(636, 10), 1888 => to_unsigned(828, 10), 1889 => to_unsigned(945, 10), 1890 => to_unsigned(917, 10), 1891 => to_unsigned(830, 10), 1892 => to_unsigned(1012, 10), 1893 => to_unsigned(942, 10), 1894 => to_unsigned(841, 10), 1895 => to_unsigned(661, 10), 1896 => to_unsigned(576, 10), 1897 => to_unsigned(827, 10), 1898 => to_unsigned(640, 10), 1899 => to_unsigned(297, 10), 1900 => to_unsigned(1003, 10), 1901 => to_unsigned(830, 10), 1902 => to_unsigned(35, 10), 1903 => to_unsigned(755, 10), 1904 => to_unsigned(885, 10), 1905 => to_unsigned(415, 10), 1906 => to_unsigned(452, 10), 1907 => to_unsigned(328, 10), 1908 => to_unsigned(240, 10), 1909 => to_unsigned(424, 10), 1910 => to_unsigned(710, 10), 1911 => to_unsigned(719, 10), 1912 => to_unsigned(628, 10), 1913 => to_unsigned(252, 10), 1914 => to_unsigned(996, 10), 1915 => to_unsigned(662, 10), 1916 => to_unsigned(341, 10), 1917 => to_unsigned(941, 10), 1918 => to_unsigned(403, 10), 1919 => to_unsigned(56, 10), 1920 => to_unsigned(150, 10), 1921 => to_unsigned(583, 10), 1922 => to_unsigned(971, 10), 1923 => to_unsigned(246, 10), 1924 => to_unsigned(783, 10), 1925 => to_unsigned(715, 10), 1926 => to_unsigned(174, 10), 1927 => to_unsigned(561, 10), 1928 => to_unsigned(521, 10), 1929 => to_unsigned(992, 10), 1930 => to_unsigned(803, 10), 1931 => to_unsigned(689, 10), 1932 => to_unsigned(674, 10), 1933 => to_unsigned(4, 10), 1934 => to_unsigned(458, 10), 1935 => to_unsigned(48, 10), 1936 => to_unsigned(434, 10), 1937 => to_unsigned(53, 10), 1938 => to_unsigned(19, 10), 1939 => to_unsigned(550, 10), 1940 => to_unsigned(88, 10), 1941 => to_unsigned(349, 10), 1942 => to_unsigned(629, 10), 1943 => to_unsigned(137, 10), 1944 => to_unsigned(881, 10), 1945 => to_unsigned(318, 10), 1946 => to_unsigned(951, 10), 1947 => to_unsigned(520, 10), 1948 => to_unsigned(695, 10), 1949 => to_unsigned(212, 10), 1950 => to_unsigned(373, 10), 1951 => to_unsigned(650, 10), 1952 => to_unsigned(297, 10), 1953 => to_unsigned(878, 10), 1954 => to_unsigned(837, 10), 1955 => to_unsigned(590, 10), 1956 => to_unsigned(601, 10), 1957 => to_unsigned(806, 10), 1958 => to_unsigned(629, 10), 1959 => to_unsigned(430, 10), 1960 => to_unsigned(4, 10), 1961 => to_unsigned(338, 10), 1962 => to_unsigned(970, 10), 1963 => to_unsigned(375, 10), 1964 => to_unsigned(102, 10), 1965 => to_unsigned(928, 10), 1966 => to_unsigned(432, 10), 1967 => to_unsigned(417, 10), 1968 => to_unsigned(862, 10), 1969 => to_unsigned(465, 10), 1970 => to_unsigned(261, 10), 1971 => to_unsigned(645, 10), 1972 => to_unsigned(563, 10), 1973 => to_unsigned(622, 10), 1974 => to_unsigned(840, 10), 1975 => to_unsigned(423, 10), 1976 => to_unsigned(655, 10), 1977 => to_unsigned(671, 10), 1978 => to_unsigned(182, 10), 1979 => to_unsigned(984, 10), 1980 => to_unsigned(995, 10), 1981 => to_unsigned(676, 10), 1982 => to_unsigned(548, 10), 1983 => to_unsigned(243, 10), 1984 => to_unsigned(762, 10), 1985 => to_unsigned(839, 10), 1986 => to_unsigned(720, 10), 1987 => to_unsigned(578, 10), 1988 => to_unsigned(306, 10), 1989 => to_unsigned(324, 10), 1990 => to_unsigned(377, 10), 1991 => to_unsigned(626, 10), 1992 => to_unsigned(737, 10), 1993 => to_unsigned(900, 10), 1994 => to_unsigned(223, 10), 1995 => to_unsigned(648, 10), 1996 => to_unsigned(11, 10), 1997 => to_unsigned(953, 10), 1998 => to_unsigned(263, 10), 1999 => to_unsigned(541, 10), 2000 => to_unsigned(975, 10), 2001 => to_unsigned(821, 10), 2002 => to_unsigned(160, 10), 2003 => to_unsigned(913, 10), 2004 => to_unsigned(397, 10), 2005 => to_unsigned(516, 10), 2006 => to_unsigned(680, 10), 2007 => to_unsigned(421, 10), 2008 => to_unsigned(608, 10), 2009 => to_unsigned(712, 10), 2010 => to_unsigned(211, 10), 2011 => to_unsigned(450, 10), 2012 => to_unsigned(582, 10), 2013 => to_unsigned(431, 10), 2014 => to_unsigned(240, 10), 2015 => to_unsigned(831, 10), 2016 => to_unsigned(432, 10), 2017 => to_unsigned(713, 10), 2018 => to_unsigned(575, 10), 2019 => to_unsigned(564, 10), 2020 => to_unsigned(765, 10), 2021 => to_unsigned(595, 10), 2022 => to_unsigned(22, 10), 2023 => to_unsigned(746, 10), 2024 => to_unsigned(582, 10), 2025 => to_unsigned(272, 10), 2026 => to_unsigned(107, 10), 2027 => to_unsigned(525, 10), 2028 => to_unsigned(367, 10), 2029 => to_unsigned(528, 10), 2030 => to_unsigned(835, 10), 2031 => to_unsigned(848, 10), 2032 => to_unsigned(834, 10), 2033 => to_unsigned(438, 10), 2034 => to_unsigned(49, 10), 2035 => to_unsigned(11, 10), 2036 => to_unsigned(624, 10), 2037 => to_unsigned(397, 10), 2038 => to_unsigned(657, 10), 2039 => to_unsigned(426, 10), 2040 => to_unsigned(647, 10), 2041 => to_unsigned(957, 10), 2042 => to_unsigned(895, 10), 2043 => to_unsigned(567, 10), 2044 => to_unsigned(433, 10), 2045 => to_unsigned(463, 10), 2046 => to_unsigned(726, 10), 2047 => to_unsigned(186, 10)),
            2 => (0 => to_unsigned(65, 10), 1 => to_unsigned(57, 10), 2 => to_unsigned(971, 10), 3 => to_unsigned(415, 10), 4 => to_unsigned(418, 10), 5 => to_unsigned(385, 10), 6 => to_unsigned(616, 10), 7 => to_unsigned(84, 10), 8 => to_unsigned(917, 10), 9 => to_unsigned(113, 10), 10 => to_unsigned(388, 10), 11 => to_unsigned(690, 10), 12 => to_unsigned(407, 10), 13 => to_unsigned(726, 10), 14 => to_unsigned(738, 10), 15 => to_unsigned(256, 10), 16 => to_unsigned(515, 10), 17 => to_unsigned(317, 10), 18 => to_unsigned(703, 10), 19 => to_unsigned(723, 10), 20 => to_unsigned(59, 10), 21 => to_unsigned(803, 10), 22 => to_unsigned(459, 10), 23 => to_unsigned(806, 10), 24 => to_unsigned(475, 10), 25 => to_unsigned(382, 10), 26 => to_unsigned(947, 10), 27 => to_unsigned(82, 10), 28 => to_unsigned(472, 10), 29 => to_unsigned(330, 10), 30 => to_unsigned(801, 10), 31 => to_unsigned(785, 10), 32 => to_unsigned(723, 10), 33 => to_unsigned(47, 10), 34 => to_unsigned(611, 10), 35 => to_unsigned(818, 10), 36 => to_unsigned(181, 10), 37 => to_unsigned(435, 10), 38 => to_unsigned(991, 10), 39 => to_unsigned(711, 10), 40 => to_unsigned(999, 10), 41 => to_unsigned(103, 10), 42 => to_unsigned(587, 10), 43 => to_unsigned(998, 10), 44 => to_unsigned(451, 10), 45 => to_unsigned(58, 10), 46 => to_unsigned(273, 10), 47 => to_unsigned(814, 10), 48 => to_unsigned(545, 10), 49 => to_unsigned(321, 10), 50 => to_unsigned(990, 10), 51 => to_unsigned(988, 10), 52 => to_unsigned(231, 10), 53 => to_unsigned(756, 10), 54 => to_unsigned(502, 10), 55 => to_unsigned(886, 10), 56 => to_unsigned(496, 10), 57 => to_unsigned(193, 10), 58 => to_unsigned(188, 10), 59 => to_unsigned(489, 10), 60 => to_unsigned(935, 10), 61 => to_unsigned(747, 10), 62 => to_unsigned(299, 10), 63 => to_unsigned(751, 10), 64 => to_unsigned(293, 10), 65 => to_unsigned(258, 10), 66 => to_unsigned(966, 10), 67 => to_unsigned(40, 10), 68 => to_unsigned(412, 10), 69 => to_unsigned(664, 10), 70 => to_unsigned(275, 10), 71 => to_unsigned(552, 10), 72 => to_unsigned(143, 10), 73 => to_unsigned(154, 10), 74 => to_unsigned(691, 10), 75 => to_unsigned(539, 10), 76 => to_unsigned(234, 10), 77 => to_unsigned(572, 10), 78 => to_unsigned(441, 10), 79 => to_unsigned(625, 10), 80 => to_unsigned(960, 10), 81 => to_unsigned(874, 10), 82 => to_unsigned(155, 10), 83 => to_unsigned(425, 10), 84 => to_unsigned(544, 10), 85 => to_unsigned(890, 10), 86 => to_unsigned(732, 10), 87 => to_unsigned(200, 10), 88 => to_unsigned(361, 10), 89 => to_unsigned(395, 10), 90 => to_unsigned(307, 10), 91 => to_unsigned(583, 10), 92 => to_unsigned(48, 10), 93 => to_unsigned(764, 10), 94 => to_unsigned(494, 10), 95 => to_unsigned(785, 10), 96 => to_unsigned(610, 10), 97 => to_unsigned(455, 10), 98 => to_unsigned(984, 10), 99 => to_unsigned(396, 10), 100 => to_unsigned(976, 10), 101 => to_unsigned(919, 10), 102 => to_unsigned(149, 10), 103 => to_unsigned(715, 10), 104 => to_unsigned(106, 10), 105 => to_unsigned(95, 10), 106 => to_unsigned(77, 10), 107 => to_unsigned(923, 10), 108 => to_unsigned(420, 10), 109 => to_unsigned(181, 10), 110 => to_unsigned(765, 10), 111 => to_unsigned(462, 10), 112 => to_unsigned(322, 10), 113 => to_unsigned(650, 10), 114 => to_unsigned(420, 10), 115 => to_unsigned(86, 10), 116 => to_unsigned(424, 10), 117 => to_unsigned(955, 10), 118 => to_unsigned(200, 10), 119 => to_unsigned(679, 10), 120 => to_unsigned(234, 10), 121 => to_unsigned(733, 10), 122 => to_unsigned(604, 10), 123 => to_unsigned(787, 10), 124 => to_unsigned(20, 10), 125 => to_unsigned(988, 10), 126 => to_unsigned(389, 10), 127 => to_unsigned(172, 10), 128 => to_unsigned(345, 10), 129 => to_unsigned(49, 10), 130 => to_unsigned(844, 10), 131 => to_unsigned(437, 10), 132 => to_unsigned(361, 10), 133 => to_unsigned(725, 10), 134 => to_unsigned(480, 10), 135 => to_unsigned(637, 10), 136 => to_unsigned(691, 10), 137 => to_unsigned(131, 10), 138 => to_unsigned(50, 10), 139 => to_unsigned(859, 10), 140 => to_unsigned(761, 10), 141 => to_unsigned(861, 10), 142 => to_unsigned(627, 10), 143 => to_unsigned(137, 10), 144 => to_unsigned(929, 10), 145 => to_unsigned(71, 10), 146 => to_unsigned(816, 10), 147 => to_unsigned(1020, 10), 148 => to_unsigned(899, 10), 149 => to_unsigned(795, 10), 150 => to_unsigned(1021, 10), 151 => to_unsigned(513, 10), 152 => to_unsigned(342, 10), 153 => to_unsigned(926, 10), 154 => to_unsigned(26, 10), 155 => to_unsigned(769, 10), 156 => to_unsigned(27, 10), 157 => to_unsigned(567, 10), 158 => to_unsigned(996, 10), 159 => to_unsigned(63, 10), 160 => to_unsigned(585, 10), 161 => to_unsigned(456, 10), 162 => to_unsigned(631, 10), 163 => to_unsigned(309, 10), 164 => to_unsigned(799, 10), 165 => to_unsigned(29, 10), 166 => to_unsigned(23, 10), 167 => to_unsigned(74, 10), 168 => to_unsigned(789, 10), 169 => to_unsigned(66, 10), 170 => to_unsigned(642, 10), 171 => to_unsigned(205, 10), 172 => to_unsigned(410, 10), 173 => to_unsigned(721, 10), 174 => to_unsigned(446, 10), 175 => to_unsigned(482, 10), 176 => to_unsigned(884, 10), 177 => to_unsigned(746, 10), 178 => to_unsigned(780, 10), 179 => to_unsigned(700, 10), 180 => to_unsigned(569, 10), 181 => to_unsigned(113, 10), 182 => to_unsigned(1010, 10), 183 => to_unsigned(158, 10), 184 => to_unsigned(43, 10), 185 => to_unsigned(517, 10), 186 => to_unsigned(14, 10), 187 => to_unsigned(917, 10), 188 => to_unsigned(541, 10), 189 => to_unsigned(447, 10), 190 => to_unsigned(949, 10), 191 => to_unsigned(141, 10), 192 => to_unsigned(733, 10), 193 => to_unsigned(561, 10), 194 => to_unsigned(195, 10), 195 => to_unsigned(745, 10), 196 => to_unsigned(315, 10), 197 => to_unsigned(740, 10), 198 => to_unsigned(1016, 10), 199 => to_unsigned(791, 10), 200 => to_unsigned(25, 10), 201 => to_unsigned(487, 10), 202 => to_unsigned(672, 10), 203 => to_unsigned(614, 10), 204 => to_unsigned(385, 10), 205 => to_unsigned(819, 10), 206 => to_unsigned(784, 10), 207 => to_unsigned(78, 10), 208 => to_unsigned(644, 10), 209 => to_unsigned(736, 10), 210 => to_unsigned(8, 10), 211 => to_unsigned(726, 10), 212 => to_unsigned(5, 10), 213 => to_unsigned(64, 10), 214 => to_unsigned(1002, 10), 215 => to_unsigned(725, 10), 216 => to_unsigned(697, 10), 217 => to_unsigned(269, 10), 218 => to_unsigned(63, 10), 219 => to_unsigned(611, 10), 220 => to_unsigned(190, 10), 221 => to_unsigned(248, 10), 222 => to_unsigned(227, 10), 223 => to_unsigned(928, 10), 224 => to_unsigned(754, 10), 225 => to_unsigned(507, 10), 226 => to_unsigned(215, 10), 227 => to_unsigned(692, 10), 228 => to_unsigned(342, 10), 229 => to_unsigned(924, 10), 230 => to_unsigned(639, 10), 231 => to_unsigned(140, 10), 232 => to_unsigned(138, 10), 233 => to_unsigned(39, 10), 234 => to_unsigned(147, 10), 235 => to_unsigned(715, 10), 236 => to_unsigned(747, 10), 237 => to_unsigned(737, 10), 238 => to_unsigned(497, 10), 239 => to_unsigned(149, 10), 240 => to_unsigned(412, 10), 241 => to_unsigned(662, 10), 242 => to_unsigned(159, 10), 243 => to_unsigned(518, 10), 244 => to_unsigned(261, 10), 245 => to_unsigned(794, 10), 246 => to_unsigned(441, 10), 247 => to_unsigned(477, 10), 248 => to_unsigned(531, 10), 249 => to_unsigned(85, 10), 250 => to_unsigned(171, 10), 251 => to_unsigned(781, 10), 252 => to_unsigned(116, 10), 253 => to_unsigned(607, 10), 254 => to_unsigned(14, 10), 255 => to_unsigned(523, 10), 256 => to_unsigned(503, 10), 257 => to_unsigned(878, 10), 258 => to_unsigned(712, 10), 259 => to_unsigned(933, 10), 260 => to_unsigned(241, 10), 261 => to_unsigned(873, 10), 262 => to_unsigned(980, 10), 263 => to_unsigned(529, 10), 264 => to_unsigned(146, 10), 265 => to_unsigned(180, 10), 266 => to_unsigned(353, 10), 267 => to_unsigned(656, 10), 268 => to_unsigned(559, 10), 269 => to_unsigned(488, 10), 270 => to_unsigned(507, 10), 271 => to_unsigned(92, 10), 272 => to_unsigned(211, 10), 273 => to_unsigned(119, 10), 274 => to_unsigned(223, 10), 275 => to_unsigned(497, 10), 276 => to_unsigned(670, 10), 277 => to_unsigned(705, 10), 278 => to_unsigned(786, 10), 279 => to_unsigned(304, 10), 280 => to_unsigned(567, 10), 281 => to_unsigned(700, 10), 282 => to_unsigned(803, 10), 283 => to_unsigned(497, 10), 284 => to_unsigned(1022, 10), 285 => to_unsigned(536, 10), 286 => to_unsigned(209, 10), 287 => to_unsigned(87, 10), 288 => to_unsigned(583, 10), 289 => to_unsigned(247, 10), 290 => to_unsigned(846, 10), 291 => to_unsigned(780, 10), 292 => to_unsigned(585, 10), 293 => to_unsigned(532, 10), 294 => to_unsigned(1004, 10), 295 => to_unsigned(688, 10), 296 => to_unsigned(390, 10), 297 => to_unsigned(976, 10), 298 => to_unsigned(628, 10), 299 => to_unsigned(366, 10), 300 => to_unsigned(19, 10), 301 => to_unsigned(481, 10), 302 => to_unsigned(527, 10), 303 => to_unsigned(17, 10), 304 => to_unsigned(371, 10), 305 => to_unsigned(749, 10), 306 => to_unsigned(113, 10), 307 => to_unsigned(872, 10), 308 => to_unsigned(98, 10), 309 => to_unsigned(605, 10), 310 => to_unsigned(702, 10), 311 => to_unsigned(442, 10), 312 => to_unsigned(888, 10), 313 => to_unsigned(855, 10), 314 => to_unsigned(355, 10), 315 => to_unsigned(268, 10), 316 => to_unsigned(946, 10), 317 => to_unsigned(7, 10), 318 => to_unsigned(279, 10), 319 => to_unsigned(148, 10), 320 => to_unsigned(451, 10), 321 => to_unsigned(56, 10), 322 => to_unsigned(38, 10), 323 => to_unsigned(879, 10), 324 => to_unsigned(901, 10), 325 => to_unsigned(383, 10), 326 => to_unsigned(752, 10), 327 => to_unsigned(813, 10), 328 => to_unsigned(808, 10), 329 => to_unsigned(256, 10), 330 => to_unsigned(429, 10), 331 => to_unsigned(409, 10), 332 => to_unsigned(685, 10), 333 => to_unsigned(701, 10), 334 => to_unsigned(251, 10), 335 => to_unsigned(949, 10), 336 => to_unsigned(675, 10), 337 => to_unsigned(752, 10), 338 => to_unsigned(907, 10), 339 => to_unsigned(973, 10), 340 => to_unsigned(782, 10), 341 => to_unsigned(931, 10), 342 => to_unsigned(631, 10), 343 => to_unsigned(280, 10), 344 => to_unsigned(36, 10), 345 => to_unsigned(151, 10), 346 => to_unsigned(1017, 10), 347 => to_unsigned(786, 10), 348 => to_unsigned(986, 10), 349 => to_unsigned(917, 10), 350 => to_unsigned(269, 10), 351 => to_unsigned(321, 10), 352 => to_unsigned(738, 10), 353 => to_unsigned(1007, 10), 354 => to_unsigned(87, 10), 355 => to_unsigned(125, 10), 356 => to_unsigned(44, 10), 357 => to_unsigned(598, 10), 358 => to_unsigned(525, 10), 359 => to_unsigned(942, 10), 360 => to_unsigned(1013, 10), 361 => to_unsigned(1006, 10), 362 => to_unsigned(510, 10), 363 => to_unsigned(192, 10), 364 => to_unsigned(94, 10), 365 => to_unsigned(786, 10), 366 => to_unsigned(698, 10), 367 => to_unsigned(296, 10), 368 => to_unsigned(698, 10), 369 => to_unsigned(775, 10), 370 => to_unsigned(806, 10), 371 => to_unsigned(473, 10), 372 => to_unsigned(266, 10), 373 => to_unsigned(866, 10), 374 => to_unsigned(951, 10), 375 => to_unsigned(105, 10), 376 => to_unsigned(858, 10), 377 => to_unsigned(947, 10), 378 => to_unsigned(427, 10), 379 => to_unsigned(922, 10), 380 => to_unsigned(199, 10), 381 => to_unsigned(414, 10), 382 => to_unsigned(105, 10), 383 => to_unsigned(686, 10), 384 => to_unsigned(311, 10), 385 => to_unsigned(79, 10), 386 => to_unsigned(553, 10), 387 => to_unsigned(739, 10), 388 => to_unsigned(852, 10), 389 => to_unsigned(608, 10), 390 => to_unsigned(24, 10), 391 => to_unsigned(367, 10), 392 => to_unsigned(674, 10), 393 => to_unsigned(59, 10), 394 => to_unsigned(810, 10), 395 => to_unsigned(263, 10), 396 => to_unsigned(352, 10), 397 => to_unsigned(122, 10), 398 => to_unsigned(24, 10), 399 => to_unsigned(783, 10), 400 => to_unsigned(573, 10), 401 => to_unsigned(1004, 10), 402 => to_unsigned(171, 10), 403 => to_unsigned(935, 10), 404 => to_unsigned(274, 10), 405 => to_unsigned(208, 10), 406 => to_unsigned(191, 10), 407 => to_unsigned(429, 10), 408 => to_unsigned(804, 10), 409 => to_unsigned(625, 10), 410 => to_unsigned(355, 10), 411 => to_unsigned(119, 10), 412 => to_unsigned(970, 10), 413 => to_unsigned(734, 10), 414 => to_unsigned(316, 10), 415 => to_unsigned(893, 10), 416 => to_unsigned(166, 10), 417 => to_unsigned(594, 10), 418 => to_unsigned(459, 10), 419 => to_unsigned(415, 10), 420 => to_unsigned(148, 10), 421 => to_unsigned(270, 10), 422 => to_unsigned(423, 10), 423 => to_unsigned(325, 10), 424 => to_unsigned(790, 10), 425 => to_unsigned(780, 10), 426 => to_unsigned(757, 10), 427 => to_unsigned(981, 10), 428 => to_unsigned(338, 10), 429 => to_unsigned(833, 10), 430 => to_unsigned(884, 10), 431 => to_unsigned(422, 10), 432 => to_unsigned(663, 10), 433 => to_unsigned(18, 10), 434 => to_unsigned(155, 10), 435 => to_unsigned(304, 10), 436 => to_unsigned(820, 10), 437 => to_unsigned(820, 10), 438 => to_unsigned(497, 10), 439 => to_unsigned(29, 10), 440 => to_unsigned(663, 10), 441 => to_unsigned(452, 10), 442 => to_unsigned(404, 10), 443 => to_unsigned(431, 10), 444 => to_unsigned(744, 10), 445 => to_unsigned(203, 10), 446 => to_unsigned(190, 10), 447 => to_unsigned(901, 10), 448 => to_unsigned(175, 10), 449 => to_unsigned(2, 10), 450 => to_unsigned(981, 10), 451 => to_unsigned(787, 10), 452 => to_unsigned(890, 10), 453 => to_unsigned(491, 10), 454 => to_unsigned(285, 10), 455 => to_unsigned(992, 10), 456 => to_unsigned(273, 10), 457 => to_unsigned(507, 10), 458 => to_unsigned(305, 10), 459 => to_unsigned(376, 10), 460 => to_unsigned(441, 10), 461 => to_unsigned(510, 10), 462 => to_unsigned(846, 10), 463 => to_unsigned(225, 10), 464 => to_unsigned(574, 10), 465 => to_unsigned(725, 10), 466 => to_unsigned(138, 10), 467 => to_unsigned(915, 10), 468 => to_unsigned(464, 10), 469 => to_unsigned(190, 10), 470 => to_unsigned(156, 10), 471 => to_unsigned(166, 10), 472 => to_unsigned(656, 10), 473 => to_unsigned(168, 10), 474 => to_unsigned(386, 10), 475 => to_unsigned(396, 10), 476 => to_unsigned(578, 10), 477 => to_unsigned(912, 10), 478 => to_unsigned(997, 10), 479 => to_unsigned(981, 10), 480 => to_unsigned(358, 10), 481 => to_unsigned(423, 10), 482 => to_unsigned(767, 10), 483 => to_unsigned(137, 10), 484 => to_unsigned(281, 10), 485 => to_unsigned(688, 10), 486 => to_unsigned(974, 10), 487 => to_unsigned(333, 10), 488 => to_unsigned(115, 10), 489 => to_unsigned(946, 10), 490 => to_unsigned(302, 10), 491 => to_unsigned(751, 10), 492 => to_unsigned(649, 10), 493 => to_unsigned(190, 10), 494 => to_unsigned(474, 10), 495 => to_unsigned(368, 10), 496 => to_unsigned(628, 10), 497 => to_unsigned(83, 10), 498 => to_unsigned(744, 10), 499 => to_unsigned(903, 10), 500 => to_unsigned(205, 10), 501 => to_unsigned(397, 10), 502 => to_unsigned(154, 10), 503 => to_unsigned(578, 10), 504 => to_unsigned(844, 10), 505 => to_unsigned(906, 10), 506 => to_unsigned(1019, 10), 507 => to_unsigned(951, 10), 508 => to_unsigned(641, 10), 509 => to_unsigned(583, 10), 510 => to_unsigned(127, 10), 511 => to_unsigned(49, 10), 512 => to_unsigned(525, 10), 513 => to_unsigned(980, 10), 514 => to_unsigned(205, 10), 515 => to_unsigned(427, 10), 516 => to_unsigned(244, 10), 517 => to_unsigned(865, 10), 518 => to_unsigned(599, 10), 519 => to_unsigned(366, 10), 520 => to_unsigned(946, 10), 521 => to_unsigned(860, 10), 522 => to_unsigned(291, 10), 523 => to_unsigned(1007, 10), 524 => to_unsigned(746, 10), 525 => to_unsigned(55, 10), 526 => to_unsigned(948, 10), 527 => to_unsigned(1006, 10), 528 => to_unsigned(355, 10), 529 => to_unsigned(510, 10), 530 => to_unsigned(922, 10), 531 => to_unsigned(655, 10), 532 => to_unsigned(937, 10), 533 => to_unsigned(561, 10), 534 => to_unsigned(893, 10), 535 => to_unsigned(242, 10), 536 => to_unsigned(107, 10), 537 => to_unsigned(281, 10), 538 => to_unsigned(620, 10), 539 => to_unsigned(864, 10), 540 => to_unsigned(732, 10), 541 => to_unsigned(9, 10), 542 => to_unsigned(427, 10), 543 => to_unsigned(65, 10), 544 => to_unsigned(104, 10), 545 => to_unsigned(681, 10), 546 => to_unsigned(636, 10), 547 => to_unsigned(145, 10), 548 => to_unsigned(164, 10), 549 => to_unsigned(415, 10), 550 => to_unsigned(359, 10), 551 => to_unsigned(904, 10), 552 => to_unsigned(331, 10), 553 => to_unsigned(715, 10), 554 => to_unsigned(943, 10), 555 => to_unsigned(721, 10), 556 => to_unsigned(364, 10), 557 => to_unsigned(503, 10), 558 => to_unsigned(485, 10), 559 => to_unsigned(627, 10), 560 => to_unsigned(116, 10), 561 => to_unsigned(701, 10), 562 => to_unsigned(51, 10), 563 => to_unsigned(69, 10), 564 => to_unsigned(833, 10), 565 => to_unsigned(206, 10), 566 => to_unsigned(776, 10), 567 => to_unsigned(130, 10), 568 => to_unsigned(720, 10), 569 => to_unsigned(915, 10), 570 => to_unsigned(312, 10), 571 => to_unsigned(533, 10), 572 => to_unsigned(943, 10), 573 => to_unsigned(560, 10), 574 => to_unsigned(863, 10), 575 => to_unsigned(73, 10), 576 => to_unsigned(454, 10), 577 => to_unsigned(893, 10), 578 => to_unsigned(800, 10), 579 => to_unsigned(65, 10), 580 => to_unsigned(171, 10), 581 => to_unsigned(51, 10), 582 => to_unsigned(93, 10), 583 => to_unsigned(924, 10), 584 => to_unsigned(94, 10), 585 => to_unsigned(710, 10), 586 => to_unsigned(225, 10), 587 => to_unsigned(998, 10), 588 => to_unsigned(960, 10), 589 => to_unsigned(825, 10), 590 => to_unsigned(181, 10), 591 => to_unsigned(532, 10), 592 => to_unsigned(621, 10), 593 => to_unsigned(189, 10), 594 => to_unsigned(506, 10), 595 => to_unsigned(993, 10), 596 => to_unsigned(961, 10), 597 => to_unsigned(358, 10), 598 => to_unsigned(82, 10), 599 => to_unsigned(463, 10), 600 => to_unsigned(697, 10), 601 => to_unsigned(658, 10), 602 => to_unsigned(161, 10), 603 => to_unsigned(194, 10), 604 => to_unsigned(614, 10), 605 => to_unsigned(385, 10), 606 => to_unsigned(874, 10), 607 => to_unsigned(859, 10), 608 => to_unsigned(207, 10), 609 => to_unsigned(260, 10), 610 => to_unsigned(35, 10), 611 => to_unsigned(971, 10), 612 => to_unsigned(387, 10), 613 => to_unsigned(523, 10), 614 => to_unsigned(242, 10), 615 => to_unsigned(987, 10), 616 => to_unsigned(108, 10), 617 => to_unsigned(990, 10), 618 => to_unsigned(181, 10), 619 => to_unsigned(553, 10), 620 => to_unsigned(242, 10), 621 => to_unsigned(286, 10), 622 => to_unsigned(751, 10), 623 => to_unsigned(1006, 10), 624 => to_unsigned(654, 10), 625 => to_unsigned(229, 10), 626 => to_unsigned(654, 10), 627 => to_unsigned(560, 10), 628 => to_unsigned(903, 10), 629 => to_unsigned(730, 10), 630 => to_unsigned(849, 10), 631 => to_unsigned(480, 10), 632 => to_unsigned(988, 10), 633 => to_unsigned(874, 10), 634 => to_unsigned(870, 10), 635 => to_unsigned(822, 10), 636 => to_unsigned(479, 10), 637 => to_unsigned(97, 10), 638 => to_unsigned(578, 10), 639 => to_unsigned(524, 10), 640 => to_unsigned(310, 10), 641 => to_unsigned(812, 10), 642 => to_unsigned(814, 10), 643 => to_unsigned(196, 10), 644 => to_unsigned(1004, 10), 645 => to_unsigned(27, 10), 646 => to_unsigned(466, 10), 647 => to_unsigned(726, 10), 648 => to_unsigned(894, 10), 649 => to_unsigned(287, 10), 650 => to_unsigned(428, 10), 651 => to_unsigned(604, 10), 652 => to_unsigned(384, 10), 653 => to_unsigned(394, 10), 654 => to_unsigned(329, 10), 655 => to_unsigned(406, 10), 656 => to_unsigned(996, 10), 657 => to_unsigned(185, 10), 658 => to_unsigned(390, 10), 659 => to_unsigned(592, 10), 660 => to_unsigned(692, 10), 661 => to_unsigned(378, 10), 662 => to_unsigned(370, 10), 663 => to_unsigned(1004, 10), 664 => to_unsigned(508, 10), 665 => to_unsigned(210, 10), 666 => to_unsigned(164, 10), 667 => to_unsigned(71, 10), 668 => to_unsigned(636, 10), 669 => to_unsigned(332, 10), 670 => to_unsigned(299, 10), 671 => to_unsigned(741, 10), 672 => to_unsigned(2, 10), 673 => to_unsigned(389, 10), 674 => to_unsigned(118, 10), 675 => to_unsigned(424, 10), 676 => to_unsigned(353, 10), 677 => to_unsigned(49, 10), 678 => to_unsigned(11, 10), 679 => to_unsigned(191, 10), 680 => to_unsigned(509, 10), 681 => to_unsigned(380, 10), 682 => to_unsigned(10, 10), 683 => to_unsigned(778, 10), 684 => to_unsigned(936, 10), 685 => to_unsigned(419, 10), 686 => to_unsigned(884, 10), 687 => to_unsigned(369, 10), 688 => to_unsigned(12, 10), 689 => to_unsigned(937, 10), 690 => to_unsigned(510, 10), 691 => to_unsigned(439, 10), 692 => to_unsigned(419, 10), 693 => to_unsigned(503, 10), 694 => to_unsigned(971, 10), 695 => to_unsigned(859, 10), 696 => to_unsigned(144, 10), 697 => to_unsigned(384, 10), 698 => to_unsigned(668, 10), 699 => to_unsigned(368, 10), 700 => to_unsigned(432, 10), 701 => to_unsigned(879, 10), 702 => to_unsigned(506, 10), 703 => to_unsigned(332, 10), 704 => to_unsigned(885, 10), 705 => to_unsigned(381, 10), 706 => to_unsigned(741, 10), 707 => to_unsigned(919, 10), 708 => to_unsigned(294, 10), 709 => to_unsigned(802, 10), 710 => to_unsigned(897, 10), 711 => to_unsigned(886, 10), 712 => to_unsigned(954, 10), 713 => to_unsigned(184, 10), 714 => to_unsigned(46, 10), 715 => to_unsigned(387, 10), 716 => to_unsigned(424, 10), 717 => to_unsigned(908, 10), 718 => to_unsigned(405, 10), 719 => to_unsigned(320, 10), 720 => to_unsigned(827, 10), 721 => to_unsigned(787, 10), 722 => to_unsigned(628, 10), 723 => to_unsigned(992, 10), 724 => to_unsigned(685, 10), 725 => to_unsigned(512, 10), 726 => to_unsigned(786, 10), 727 => to_unsigned(703, 10), 728 => to_unsigned(439, 10), 729 => to_unsigned(465, 10), 730 => to_unsigned(153, 10), 731 => to_unsigned(689, 10), 732 => to_unsigned(645, 10), 733 => to_unsigned(904, 10), 734 => to_unsigned(578, 10), 735 => to_unsigned(102, 10), 736 => to_unsigned(711, 10), 737 => to_unsigned(58, 10), 738 => to_unsigned(545, 10), 739 => to_unsigned(752, 10), 740 => to_unsigned(278, 10), 741 => to_unsigned(905, 10), 742 => to_unsigned(869, 10), 743 => to_unsigned(339, 10), 744 => to_unsigned(694, 10), 745 => to_unsigned(98, 10), 746 => to_unsigned(380, 10), 747 => to_unsigned(978, 10), 748 => to_unsigned(325, 10), 749 => to_unsigned(327, 10), 750 => to_unsigned(210, 10), 751 => to_unsigned(137, 10), 752 => to_unsigned(464, 10), 753 => to_unsigned(641, 10), 754 => to_unsigned(990, 10), 755 => to_unsigned(857, 10), 756 => to_unsigned(37, 10), 757 => to_unsigned(312, 10), 758 => to_unsigned(701, 10), 759 => to_unsigned(182, 10), 760 => to_unsigned(333, 10), 761 => to_unsigned(217, 10), 762 => to_unsigned(159, 10), 763 => to_unsigned(580, 10), 764 => to_unsigned(994, 10), 765 => to_unsigned(1012, 10), 766 => to_unsigned(254, 10), 767 => to_unsigned(584, 10), 768 => to_unsigned(128, 10), 769 => to_unsigned(395, 10), 770 => to_unsigned(17, 10), 771 => to_unsigned(553, 10), 772 => to_unsigned(807, 10), 773 => to_unsigned(379, 10), 774 => to_unsigned(693, 10), 775 => to_unsigned(111, 10), 776 => to_unsigned(267, 10), 777 => to_unsigned(477, 10), 778 => to_unsigned(801, 10), 779 => to_unsigned(829, 10), 780 => to_unsigned(549, 10), 781 => to_unsigned(1023, 10), 782 => to_unsigned(741, 10), 783 => to_unsigned(629, 10), 784 => to_unsigned(303, 10), 785 => to_unsigned(657, 10), 786 => to_unsigned(934, 10), 787 => to_unsigned(985, 10), 788 => to_unsigned(582, 10), 789 => to_unsigned(42, 10), 790 => to_unsigned(936, 10), 791 => to_unsigned(598, 10), 792 => to_unsigned(386, 10), 793 => to_unsigned(164, 10), 794 => to_unsigned(274, 10), 795 => to_unsigned(348, 10), 796 => to_unsigned(66, 10), 797 => to_unsigned(257, 10), 798 => to_unsigned(850, 10), 799 => to_unsigned(914, 10), 800 => to_unsigned(876, 10), 801 => to_unsigned(386, 10), 802 => to_unsigned(148, 10), 803 => to_unsigned(500, 10), 804 => to_unsigned(719, 10), 805 => to_unsigned(539, 10), 806 => to_unsigned(504, 10), 807 => to_unsigned(954, 10), 808 => to_unsigned(343, 10), 809 => to_unsigned(201, 10), 810 => to_unsigned(563, 10), 811 => to_unsigned(468, 10), 812 => to_unsigned(584, 10), 813 => to_unsigned(410, 10), 814 => to_unsigned(375, 10), 815 => to_unsigned(196, 10), 816 => to_unsigned(1003, 10), 817 => to_unsigned(895, 10), 818 => to_unsigned(291, 10), 819 => to_unsigned(393, 10), 820 => to_unsigned(394, 10), 821 => to_unsigned(24, 10), 822 => to_unsigned(553, 10), 823 => to_unsigned(722, 10), 824 => to_unsigned(81, 10), 825 => to_unsigned(538, 10), 826 => to_unsigned(547, 10), 827 => to_unsigned(404, 10), 828 => to_unsigned(856, 10), 829 => to_unsigned(809, 10), 830 => to_unsigned(358, 10), 831 => to_unsigned(835, 10), 832 => to_unsigned(1014, 10), 833 => to_unsigned(671, 10), 834 => to_unsigned(505, 10), 835 => to_unsigned(30, 10), 836 => to_unsigned(697, 10), 837 => to_unsigned(325, 10), 838 => to_unsigned(881, 10), 839 => to_unsigned(870, 10), 840 => to_unsigned(918, 10), 841 => to_unsigned(491, 10), 842 => to_unsigned(605, 10), 843 => to_unsigned(438, 10), 844 => to_unsigned(1002, 10), 845 => to_unsigned(1007, 10), 846 => to_unsigned(637, 10), 847 => to_unsigned(1007, 10), 848 => to_unsigned(312, 10), 849 => to_unsigned(633, 10), 850 => to_unsigned(745, 10), 851 => to_unsigned(221, 10), 852 => to_unsigned(695, 10), 853 => to_unsigned(5, 10), 854 => to_unsigned(124, 10), 855 => to_unsigned(55, 10), 856 => to_unsigned(45, 10), 857 => to_unsigned(44, 10), 858 => to_unsigned(204, 10), 859 => to_unsigned(944, 10), 860 => to_unsigned(428, 10), 861 => to_unsigned(72, 10), 862 => to_unsigned(846, 10), 863 => to_unsigned(360, 10), 864 => to_unsigned(308, 10), 865 => to_unsigned(530, 10), 866 => to_unsigned(733, 10), 867 => to_unsigned(490, 10), 868 => to_unsigned(806, 10), 869 => to_unsigned(538, 10), 870 => to_unsigned(594, 10), 871 => to_unsigned(138, 10), 872 => to_unsigned(217, 10), 873 => to_unsigned(642, 10), 874 => to_unsigned(823, 10), 875 => to_unsigned(222, 10), 876 => to_unsigned(738, 10), 877 => to_unsigned(281, 10), 878 => to_unsigned(374, 10), 879 => to_unsigned(6, 10), 880 => to_unsigned(615, 10), 881 => to_unsigned(239, 10), 882 => to_unsigned(290, 10), 883 => to_unsigned(579, 10), 884 => to_unsigned(12, 10), 885 => to_unsigned(528, 10), 886 => to_unsigned(916, 10), 887 => to_unsigned(417, 10), 888 => to_unsigned(459, 10), 889 => to_unsigned(625, 10), 890 => to_unsigned(796, 10), 891 => to_unsigned(729, 10), 892 => to_unsigned(103, 10), 893 => to_unsigned(787, 10), 894 => to_unsigned(230, 10), 895 => to_unsigned(988, 10), 896 => to_unsigned(554, 10), 897 => to_unsigned(694, 10), 898 => to_unsigned(414, 10), 899 => to_unsigned(52, 10), 900 => to_unsigned(203, 10), 901 => to_unsigned(332, 10), 902 => to_unsigned(492, 10), 903 => to_unsigned(890, 10), 904 => to_unsigned(544, 10), 905 => to_unsigned(539, 10), 906 => to_unsigned(300, 10), 907 => to_unsigned(303, 10), 908 => to_unsigned(238, 10), 909 => to_unsigned(46, 10), 910 => to_unsigned(209, 10), 911 => to_unsigned(846, 10), 912 => to_unsigned(367, 10), 913 => to_unsigned(323, 10), 914 => to_unsigned(113, 10), 915 => to_unsigned(56, 10), 916 => to_unsigned(763, 10), 917 => to_unsigned(65, 10), 918 => to_unsigned(590, 10), 919 => to_unsigned(165, 10), 920 => to_unsigned(835, 10), 921 => to_unsigned(1021, 10), 922 => to_unsigned(154, 10), 923 => to_unsigned(37, 10), 924 => to_unsigned(976, 10), 925 => to_unsigned(377, 10), 926 => to_unsigned(24, 10), 927 => to_unsigned(583, 10), 928 => to_unsigned(1008, 10), 929 => to_unsigned(74, 10), 930 => to_unsigned(886, 10), 931 => to_unsigned(489, 10), 932 => to_unsigned(829, 10), 933 => to_unsigned(219, 10), 934 => to_unsigned(895, 10), 935 => to_unsigned(338, 10), 936 => to_unsigned(583, 10), 937 => to_unsigned(974, 10), 938 => to_unsigned(779, 10), 939 => to_unsigned(865, 10), 940 => to_unsigned(168, 10), 941 => to_unsigned(715, 10), 942 => to_unsigned(719, 10), 943 => to_unsigned(13, 10), 944 => to_unsigned(270, 10), 945 => to_unsigned(514, 10), 946 => to_unsigned(614, 10), 947 => to_unsigned(655, 10), 948 => to_unsigned(525, 10), 949 => to_unsigned(1000, 10), 950 => to_unsigned(425, 10), 951 => to_unsigned(650, 10), 952 => to_unsigned(928, 10), 953 => to_unsigned(750, 10), 954 => to_unsigned(39, 10), 955 => to_unsigned(39, 10), 956 => to_unsigned(21, 10), 957 => to_unsigned(430, 10), 958 => to_unsigned(629, 10), 959 => to_unsigned(149, 10), 960 => to_unsigned(981, 10), 961 => to_unsigned(821, 10), 962 => to_unsigned(1000, 10), 963 => to_unsigned(103, 10), 964 => to_unsigned(212, 10), 965 => to_unsigned(241, 10), 966 => to_unsigned(332, 10), 967 => to_unsigned(368, 10), 968 => to_unsigned(719, 10), 969 => to_unsigned(490, 10), 970 => to_unsigned(999, 10), 971 => to_unsigned(747, 10), 972 => to_unsigned(572, 10), 973 => to_unsigned(67, 10), 974 => to_unsigned(844, 10), 975 => to_unsigned(5, 10), 976 => to_unsigned(938, 10), 977 => to_unsigned(166, 10), 978 => to_unsigned(111, 10), 979 => to_unsigned(152, 10), 980 => to_unsigned(255, 10), 981 => to_unsigned(867, 10), 982 => to_unsigned(543, 10), 983 => to_unsigned(851, 10), 984 => to_unsigned(627, 10), 985 => to_unsigned(987, 10), 986 => to_unsigned(528, 10), 987 => to_unsigned(715, 10), 988 => to_unsigned(104, 10), 989 => to_unsigned(765, 10), 990 => to_unsigned(895, 10), 991 => to_unsigned(536, 10), 992 => to_unsigned(752, 10), 993 => to_unsigned(1004, 10), 994 => to_unsigned(107, 10), 995 => to_unsigned(83, 10), 996 => to_unsigned(814, 10), 997 => to_unsigned(660, 10), 998 => to_unsigned(40, 10), 999 => to_unsigned(261, 10), 1000 => to_unsigned(906, 10), 1001 => to_unsigned(115, 10), 1002 => to_unsigned(22, 10), 1003 => to_unsigned(30, 10), 1004 => to_unsigned(227, 10), 1005 => to_unsigned(39, 10), 1006 => to_unsigned(426, 10), 1007 => to_unsigned(849, 10), 1008 => to_unsigned(387, 10), 1009 => to_unsigned(432, 10), 1010 => to_unsigned(933, 10), 1011 => to_unsigned(419, 10), 1012 => to_unsigned(578, 10), 1013 => to_unsigned(1008, 10), 1014 => to_unsigned(132, 10), 1015 => to_unsigned(184, 10), 1016 => to_unsigned(484, 10), 1017 => to_unsigned(148, 10), 1018 => to_unsigned(49, 10), 1019 => to_unsigned(317, 10), 1020 => to_unsigned(532, 10), 1021 => to_unsigned(349, 10), 1022 => to_unsigned(504, 10), 1023 => to_unsigned(207, 10), 1024 => to_unsigned(428, 10), 1025 => to_unsigned(466, 10), 1026 => to_unsigned(44, 10), 1027 => to_unsigned(548, 10), 1028 => to_unsigned(65, 10), 1029 => to_unsigned(995, 10), 1030 => to_unsigned(524, 10), 1031 => to_unsigned(832, 10), 1032 => to_unsigned(777, 10), 1033 => to_unsigned(398, 10), 1034 => to_unsigned(318, 10), 1035 => to_unsigned(610, 10), 1036 => to_unsigned(974, 10), 1037 => to_unsigned(815, 10), 1038 => to_unsigned(502, 10), 1039 => to_unsigned(571, 10), 1040 => to_unsigned(904, 10), 1041 => to_unsigned(181, 10), 1042 => to_unsigned(517, 10), 1043 => to_unsigned(554, 10), 1044 => to_unsigned(929, 10), 1045 => to_unsigned(261, 10), 1046 => to_unsigned(618, 10), 1047 => to_unsigned(163, 10), 1048 => to_unsigned(519, 10), 1049 => to_unsigned(36, 10), 1050 => to_unsigned(315, 10), 1051 => to_unsigned(147, 10), 1052 => to_unsigned(98, 10), 1053 => to_unsigned(335, 10), 1054 => to_unsigned(413, 10), 1055 => to_unsigned(816, 10), 1056 => to_unsigned(599, 10), 1057 => to_unsigned(247, 10), 1058 => to_unsigned(691, 10), 1059 => to_unsigned(349, 10), 1060 => to_unsigned(858, 10), 1061 => to_unsigned(839, 10), 1062 => to_unsigned(86, 10), 1063 => to_unsigned(306, 10), 1064 => to_unsigned(725, 10), 1065 => to_unsigned(741, 10), 1066 => to_unsigned(389, 10), 1067 => to_unsigned(541, 10), 1068 => to_unsigned(412, 10), 1069 => to_unsigned(342, 10), 1070 => to_unsigned(513, 10), 1071 => to_unsigned(125, 10), 1072 => to_unsigned(452, 10), 1073 => to_unsigned(887, 10), 1074 => to_unsigned(50, 10), 1075 => to_unsigned(726, 10), 1076 => to_unsigned(708, 10), 1077 => to_unsigned(878, 10), 1078 => to_unsigned(268, 10), 1079 => to_unsigned(715, 10), 1080 => to_unsigned(39, 10), 1081 => to_unsigned(222, 10), 1082 => to_unsigned(876, 10), 1083 => to_unsigned(23, 10), 1084 => to_unsigned(142, 10), 1085 => to_unsigned(114, 10), 1086 => to_unsigned(669, 10), 1087 => to_unsigned(446, 10), 1088 => to_unsigned(302, 10), 1089 => to_unsigned(859, 10), 1090 => to_unsigned(955, 10), 1091 => to_unsigned(9, 10), 1092 => to_unsigned(606, 10), 1093 => to_unsigned(71, 10), 1094 => to_unsigned(108, 10), 1095 => to_unsigned(717, 10), 1096 => to_unsigned(632, 10), 1097 => to_unsigned(798, 10), 1098 => to_unsigned(785, 10), 1099 => to_unsigned(707, 10), 1100 => to_unsigned(718, 10), 1101 => to_unsigned(446, 10), 1102 => to_unsigned(366, 10), 1103 => to_unsigned(344, 10), 1104 => to_unsigned(400, 10), 1105 => to_unsigned(753, 10), 1106 => to_unsigned(159, 10), 1107 => to_unsigned(512, 10), 1108 => to_unsigned(676, 10), 1109 => to_unsigned(249, 10), 1110 => to_unsigned(677, 10), 1111 => to_unsigned(646, 10), 1112 => to_unsigned(883, 10), 1113 => to_unsigned(906, 10), 1114 => to_unsigned(708, 10), 1115 => to_unsigned(381, 10), 1116 => to_unsigned(733, 10), 1117 => to_unsigned(747, 10), 1118 => to_unsigned(1021, 10), 1119 => to_unsigned(561, 10), 1120 => to_unsigned(108, 10), 1121 => to_unsigned(727, 10), 1122 => to_unsigned(896, 10), 1123 => to_unsigned(952, 10), 1124 => to_unsigned(348, 10), 1125 => to_unsigned(732, 10), 1126 => to_unsigned(745, 10), 1127 => to_unsigned(266, 10), 1128 => to_unsigned(567, 10), 1129 => to_unsigned(245, 10), 1130 => to_unsigned(632, 10), 1131 => to_unsigned(2, 10), 1132 => to_unsigned(668, 10), 1133 => to_unsigned(492, 10), 1134 => to_unsigned(852, 10), 1135 => to_unsigned(865, 10), 1136 => to_unsigned(965, 10), 1137 => to_unsigned(267, 10), 1138 => to_unsigned(956, 10), 1139 => to_unsigned(785, 10), 1140 => to_unsigned(191, 10), 1141 => to_unsigned(378, 10), 1142 => to_unsigned(947, 10), 1143 => to_unsigned(331, 10), 1144 => to_unsigned(306, 10), 1145 => to_unsigned(87, 10), 1146 => to_unsigned(210, 10), 1147 => to_unsigned(613, 10), 1148 => to_unsigned(399, 10), 1149 => to_unsigned(424, 10), 1150 => to_unsigned(380, 10), 1151 => to_unsigned(133, 10), 1152 => to_unsigned(612, 10), 1153 => to_unsigned(482, 10), 1154 => to_unsigned(274, 10), 1155 => to_unsigned(61, 10), 1156 => to_unsigned(694, 10), 1157 => to_unsigned(324, 10), 1158 => to_unsigned(916, 10), 1159 => to_unsigned(258, 10), 1160 => to_unsigned(621, 10), 1161 => to_unsigned(275, 10), 1162 => to_unsigned(898, 10), 1163 => to_unsigned(364, 10), 1164 => to_unsigned(241, 10), 1165 => to_unsigned(687, 10), 1166 => to_unsigned(1017, 10), 1167 => to_unsigned(350, 10), 1168 => to_unsigned(353, 10), 1169 => to_unsigned(959, 10), 1170 => to_unsigned(905, 10), 1171 => to_unsigned(523, 10), 1172 => to_unsigned(902, 10), 1173 => to_unsigned(563, 10), 1174 => to_unsigned(462, 10), 1175 => to_unsigned(530, 10), 1176 => to_unsigned(325, 10), 1177 => to_unsigned(860, 10), 1178 => to_unsigned(892, 10), 1179 => to_unsigned(444, 10), 1180 => to_unsigned(608, 10), 1181 => to_unsigned(879, 10), 1182 => to_unsigned(2, 10), 1183 => to_unsigned(748, 10), 1184 => to_unsigned(805, 10), 1185 => to_unsigned(675, 10), 1186 => to_unsigned(67, 10), 1187 => to_unsigned(970, 10), 1188 => to_unsigned(91, 10), 1189 => to_unsigned(861, 10), 1190 => to_unsigned(579, 10), 1191 => to_unsigned(63, 10), 1192 => to_unsigned(349, 10), 1193 => to_unsigned(836, 10), 1194 => to_unsigned(673, 10), 1195 => to_unsigned(377, 10), 1196 => to_unsigned(92, 10), 1197 => to_unsigned(839, 10), 1198 => to_unsigned(960, 10), 1199 => to_unsigned(233, 10), 1200 => to_unsigned(171, 10), 1201 => to_unsigned(11, 10), 1202 => to_unsigned(497, 10), 1203 => to_unsigned(179, 10), 1204 => to_unsigned(779, 10), 1205 => to_unsigned(598, 10), 1206 => to_unsigned(952, 10), 1207 => to_unsigned(292, 10), 1208 => to_unsigned(267, 10), 1209 => to_unsigned(595, 10), 1210 => to_unsigned(142, 10), 1211 => to_unsigned(484, 10), 1212 => to_unsigned(663, 10), 1213 => to_unsigned(494, 10), 1214 => to_unsigned(229, 10), 1215 => to_unsigned(978, 10), 1216 => to_unsigned(542, 10), 1217 => to_unsigned(994, 10), 1218 => to_unsigned(255, 10), 1219 => to_unsigned(1, 10), 1220 => to_unsigned(933, 10), 1221 => to_unsigned(79, 10), 1222 => to_unsigned(682, 10), 1223 => to_unsigned(358, 10), 1224 => to_unsigned(882, 10), 1225 => to_unsigned(299, 10), 1226 => to_unsigned(185, 10), 1227 => to_unsigned(32, 10), 1228 => to_unsigned(493, 10), 1229 => to_unsigned(927, 10), 1230 => to_unsigned(851, 10), 1231 => to_unsigned(975, 10), 1232 => to_unsigned(874, 10), 1233 => to_unsigned(9, 10), 1234 => to_unsigned(263, 10), 1235 => to_unsigned(253, 10), 1236 => to_unsigned(552, 10), 1237 => to_unsigned(219, 10), 1238 => to_unsigned(899, 10), 1239 => to_unsigned(956, 10), 1240 => to_unsigned(347, 10), 1241 => to_unsigned(787, 10), 1242 => to_unsigned(117, 10), 1243 => to_unsigned(919, 10), 1244 => to_unsigned(41, 10), 1245 => to_unsigned(1003, 10), 1246 => to_unsigned(819, 10), 1247 => to_unsigned(195, 10), 1248 => to_unsigned(653, 10), 1249 => to_unsigned(900, 10), 1250 => to_unsigned(657, 10), 1251 => to_unsigned(776, 10), 1252 => to_unsigned(186, 10), 1253 => to_unsigned(509, 10), 1254 => to_unsigned(150, 10), 1255 => to_unsigned(900, 10), 1256 => to_unsigned(324, 10), 1257 => to_unsigned(932, 10), 1258 => to_unsigned(49, 10), 1259 => to_unsigned(447, 10), 1260 => to_unsigned(599, 10), 1261 => to_unsigned(121, 10), 1262 => to_unsigned(213, 10), 1263 => to_unsigned(252, 10), 1264 => to_unsigned(25, 10), 1265 => to_unsigned(27, 10), 1266 => to_unsigned(549, 10), 1267 => to_unsigned(457, 10), 1268 => to_unsigned(364, 10), 1269 => to_unsigned(310, 10), 1270 => to_unsigned(57, 10), 1271 => to_unsigned(683, 10), 1272 => to_unsigned(128, 10), 1273 => to_unsigned(282, 10), 1274 => to_unsigned(711, 10), 1275 => to_unsigned(107, 10), 1276 => to_unsigned(788, 10), 1277 => to_unsigned(0, 10), 1278 => to_unsigned(538, 10), 1279 => to_unsigned(339, 10), 1280 => to_unsigned(276, 10), 1281 => to_unsigned(645, 10), 1282 => to_unsigned(227, 10), 1283 => to_unsigned(69, 10), 1284 => to_unsigned(876, 10), 1285 => to_unsigned(994, 10), 1286 => to_unsigned(486, 10), 1287 => to_unsigned(788, 10), 1288 => to_unsigned(917, 10), 1289 => to_unsigned(988, 10), 1290 => to_unsigned(276, 10), 1291 => to_unsigned(685, 10), 1292 => to_unsigned(504, 10), 1293 => to_unsigned(300, 10), 1294 => to_unsigned(365, 10), 1295 => to_unsigned(900, 10), 1296 => to_unsigned(861, 10), 1297 => to_unsigned(576, 10), 1298 => to_unsigned(566, 10), 1299 => to_unsigned(638, 10), 1300 => to_unsigned(36, 10), 1301 => to_unsigned(455, 10), 1302 => to_unsigned(920, 10), 1303 => to_unsigned(98, 10), 1304 => to_unsigned(849, 10), 1305 => to_unsigned(929, 10), 1306 => to_unsigned(195, 10), 1307 => to_unsigned(192, 10), 1308 => to_unsigned(116, 10), 1309 => to_unsigned(680, 10), 1310 => to_unsigned(846, 10), 1311 => to_unsigned(774, 10), 1312 => to_unsigned(790, 10), 1313 => to_unsigned(453, 10), 1314 => to_unsigned(708, 10), 1315 => to_unsigned(755, 10), 1316 => to_unsigned(286, 10), 1317 => to_unsigned(83, 10), 1318 => to_unsigned(103, 10), 1319 => to_unsigned(655, 10), 1320 => to_unsigned(381, 10), 1321 => to_unsigned(314, 10), 1322 => to_unsigned(345, 10), 1323 => to_unsigned(225, 10), 1324 => to_unsigned(1007, 10), 1325 => to_unsigned(149, 10), 1326 => to_unsigned(299, 10), 1327 => to_unsigned(318, 10), 1328 => to_unsigned(846, 10), 1329 => to_unsigned(178, 10), 1330 => to_unsigned(1005, 10), 1331 => to_unsigned(577, 10), 1332 => to_unsigned(744, 10), 1333 => to_unsigned(626, 10), 1334 => to_unsigned(64, 10), 1335 => to_unsigned(827, 10), 1336 => to_unsigned(524, 10), 1337 => to_unsigned(949, 10), 1338 => to_unsigned(232, 10), 1339 => to_unsigned(452, 10), 1340 => to_unsigned(48, 10), 1341 => to_unsigned(122, 10), 1342 => to_unsigned(326, 10), 1343 => to_unsigned(505, 10), 1344 => to_unsigned(940, 10), 1345 => to_unsigned(205, 10), 1346 => to_unsigned(632, 10), 1347 => to_unsigned(633, 10), 1348 => to_unsigned(183, 10), 1349 => to_unsigned(479, 10), 1350 => to_unsigned(926, 10), 1351 => to_unsigned(1001, 10), 1352 => to_unsigned(583, 10), 1353 => to_unsigned(356, 10), 1354 => to_unsigned(571, 10), 1355 => to_unsigned(790, 10), 1356 => to_unsigned(274, 10), 1357 => to_unsigned(623, 10), 1358 => to_unsigned(457, 10), 1359 => to_unsigned(740, 10), 1360 => to_unsigned(795, 10), 1361 => to_unsigned(274, 10), 1362 => to_unsigned(483, 10), 1363 => to_unsigned(22, 10), 1364 => to_unsigned(338, 10), 1365 => to_unsigned(556, 10), 1366 => to_unsigned(817, 10), 1367 => to_unsigned(746, 10), 1368 => to_unsigned(742, 10), 1369 => to_unsigned(517, 10), 1370 => to_unsigned(947, 10), 1371 => to_unsigned(48, 10), 1372 => to_unsigned(114, 10), 1373 => to_unsigned(283, 10), 1374 => to_unsigned(642, 10), 1375 => to_unsigned(78, 10), 1376 => to_unsigned(304, 10), 1377 => to_unsigned(89, 10), 1378 => to_unsigned(705, 10), 1379 => to_unsigned(159, 10), 1380 => to_unsigned(739, 10), 1381 => to_unsigned(886, 10), 1382 => to_unsigned(533, 10), 1383 => to_unsigned(864, 10), 1384 => to_unsigned(199, 10), 1385 => to_unsigned(558, 10), 1386 => to_unsigned(569, 10), 1387 => to_unsigned(842, 10), 1388 => to_unsigned(777, 10), 1389 => to_unsigned(688, 10), 1390 => to_unsigned(310, 10), 1391 => to_unsigned(539, 10), 1392 => to_unsigned(891, 10), 1393 => to_unsigned(416, 10), 1394 => to_unsigned(398, 10), 1395 => to_unsigned(993, 10), 1396 => to_unsigned(519, 10), 1397 => to_unsigned(997, 10), 1398 => to_unsigned(126, 10), 1399 => to_unsigned(165, 10), 1400 => to_unsigned(399, 10), 1401 => to_unsigned(355, 10), 1402 => to_unsigned(594, 10), 1403 => to_unsigned(589, 10), 1404 => to_unsigned(98, 10), 1405 => to_unsigned(655, 10), 1406 => to_unsigned(236, 10), 1407 => to_unsigned(983, 10), 1408 => to_unsigned(415, 10), 1409 => to_unsigned(426, 10), 1410 => to_unsigned(179, 10), 1411 => to_unsigned(766, 10), 1412 => to_unsigned(911, 10), 1413 => to_unsigned(186, 10), 1414 => to_unsigned(294, 10), 1415 => to_unsigned(163, 10), 1416 => to_unsigned(394, 10), 1417 => to_unsigned(41, 10), 1418 => to_unsigned(599, 10), 1419 => to_unsigned(579, 10), 1420 => to_unsigned(378, 10), 1421 => to_unsigned(941, 10), 1422 => to_unsigned(483, 10), 1423 => to_unsigned(890, 10), 1424 => to_unsigned(425, 10), 1425 => to_unsigned(242, 10), 1426 => to_unsigned(770, 10), 1427 => to_unsigned(828, 10), 1428 => to_unsigned(530, 10), 1429 => to_unsigned(101, 10), 1430 => to_unsigned(227, 10), 1431 => to_unsigned(845, 10), 1432 => to_unsigned(155, 10), 1433 => to_unsigned(1023, 10), 1434 => to_unsigned(704, 10), 1435 => to_unsigned(407, 10), 1436 => to_unsigned(278, 10), 1437 => to_unsigned(847, 10), 1438 => to_unsigned(790, 10), 1439 => to_unsigned(189, 10), 1440 => to_unsigned(252, 10), 1441 => to_unsigned(235, 10), 1442 => to_unsigned(653, 10), 1443 => to_unsigned(594, 10), 1444 => to_unsigned(107, 10), 1445 => to_unsigned(664, 10), 1446 => to_unsigned(480, 10), 1447 => to_unsigned(549, 10), 1448 => to_unsigned(733, 10), 1449 => to_unsigned(732, 10), 1450 => to_unsigned(473, 10), 1451 => to_unsigned(453, 10), 1452 => to_unsigned(679, 10), 1453 => to_unsigned(572, 10), 1454 => to_unsigned(958, 10), 1455 => to_unsigned(229, 10), 1456 => to_unsigned(107, 10), 1457 => to_unsigned(175, 10), 1458 => to_unsigned(1019, 10), 1459 => to_unsigned(720, 10), 1460 => to_unsigned(163, 10), 1461 => to_unsigned(105, 10), 1462 => to_unsigned(92, 10), 1463 => to_unsigned(135, 10), 1464 => to_unsigned(386, 10), 1465 => to_unsigned(88, 10), 1466 => to_unsigned(607, 10), 1467 => to_unsigned(137, 10), 1468 => to_unsigned(251, 10), 1469 => to_unsigned(427, 10), 1470 => to_unsigned(122, 10), 1471 => to_unsigned(817, 10), 1472 => to_unsigned(680, 10), 1473 => to_unsigned(440, 10), 1474 => to_unsigned(597, 10), 1475 => to_unsigned(52, 10), 1476 => to_unsigned(578, 10), 1477 => to_unsigned(605, 10), 1478 => to_unsigned(532, 10), 1479 => to_unsigned(179, 10), 1480 => to_unsigned(366, 10), 1481 => to_unsigned(830, 10), 1482 => to_unsigned(482, 10), 1483 => to_unsigned(334, 10), 1484 => to_unsigned(812, 10), 1485 => to_unsigned(772, 10), 1486 => to_unsigned(156, 10), 1487 => to_unsigned(739, 10), 1488 => to_unsigned(930, 10), 1489 => to_unsigned(247, 10), 1490 => to_unsigned(435, 10), 1491 => to_unsigned(836, 10), 1492 => to_unsigned(277, 10), 1493 => to_unsigned(289, 10), 1494 => to_unsigned(719, 10), 1495 => to_unsigned(209, 10), 1496 => to_unsigned(802, 10), 1497 => to_unsigned(802, 10), 1498 => to_unsigned(630, 10), 1499 => to_unsigned(484, 10), 1500 => to_unsigned(726, 10), 1501 => to_unsigned(460, 10), 1502 => to_unsigned(346, 10), 1503 => to_unsigned(880, 10), 1504 => to_unsigned(160, 10), 1505 => to_unsigned(898, 10), 1506 => to_unsigned(928, 10), 1507 => to_unsigned(161, 10), 1508 => to_unsigned(521, 10), 1509 => to_unsigned(199, 10), 1510 => to_unsigned(407, 10), 1511 => to_unsigned(455, 10), 1512 => to_unsigned(139, 10), 1513 => to_unsigned(726, 10), 1514 => to_unsigned(163, 10), 1515 => to_unsigned(152, 10), 1516 => to_unsigned(201, 10), 1517 => to_unsigned(981, 10), 1518 => to_unsigned(46, 10), 1519 => to_unsigned(791, 10), 1520 => to_unsigned(683, 10), 1521 => to_unsigned(23, 10), 1522 => to_unsigned(344, 10), 1523 => to_unsigned(134, 10), 1524 => to_unsigned(916, 10), 1525 => to_unsigned(484, 10), 1526 => to_unsigned(302, 10), 1527 => to_unsigned(416, 10), 1528 => to_unsigned(298, 10), 1529 => to_unsigned(915, 10), 1530 => to_unsigned(576, 10), 1531 => to_unsigned(446, 10), 1532 => to_unsigned(772, 10), 1533 => to_unsigned(85, 10), 1534 => to_unsigned(184, 10), 1535 => to_unsigned(671, 10), 1536 => to_unsigned(688, 10), 1537 => to_unsigned(711, 10), 1538 => to_unsigned(177, 10), 1539 => to_unsigned(1008, 10), 1540 => to_unsigned(112, 10), 1541 => to_unsigned(524, 10), 1542 => to_unsigned(657, 10), 1543 => to_unsigned(925, 10), 1544 => to_unsigned(1016, 10), 1545 => to_unsigned(179, 10), 1546 => to_unsigned(387, 10), 1547 => to_unsigned(158, 10), 1548 => to_unsigned(90, 10), 1549 => to_unsigned(557, 10), 1550 => to_unsigned(663, 10), 1551 => to_unsigned(377, 10), 1552 => to_unsigned(481, 10), 1553 => to_unsigned(721, 10), 1554 => to_unsigned(274, 10), 1555 => to_unsigned(733, 10), 1556 => to_unsigned(450, 10), 1557 => to_unsigned(916, 10), 1558 => to_unsigned(48, 10), 1559 => to_unsigned(533, 10), 1560 => to_unsigned(190, 10), 1561 => to_unsigned(740, 10), 1562 => to_unsigned(285, 10), 1563 => to_unsigned(324, 10), 1564 => to_unsigned(169, 10), 1565 => to_unsigned(445, 10), 1566 => to_unsigned(286, 10), 1567 => to_unsigned(114, 10), 1568 => to_unsigned(363, 10), 1569 => to_unsigned(490, 10), 1570 => to_unsigned(642, 10), 1571 => to_unsigned(520, 10), 1572 => to_unsigned(251, 10), 1573 => to_unsigned(972, 10), 1574 => to_unsigned(249, 10), 1575 => to_unsigned(902, 10), 1576 => to_unsigned(682, 10), 1577 => to_unsigned(941, 10), 1578 => to_unsigned(819, 10), 1579 => to_unsigned(601, 10), 1580 => to_unsigned(932, 10), 1581 => to_unsigned(407, 10), 1582 => to_unsigned(128, 10), 1583 => to_unsigned(368, 10), 1584 => to_unsigned(513, 10), 1585 => to_unsigned(170, 10), 1586 => to_unsigned(794, 10), 1587 => to_unsigned(688, 10), 1588 => to_unsigned(176, 10), 1589 => to_unsigned(456, 10), 1590 => to_unsigned(402, 10), 1591 => to_unsigned(18, 10), 1592 => to_unsigned(269, 10), 1593 => to_unsigned(135, 10), 1594 => to_unsigned(364, 10), 1595 => to_unsigned(741, 10), 1596 => to_unsigned(387, 10), 1597 => to_unsigned(404, 10), 1598 => to_unsigned(950, 10), 1599 => to_unsigned(234, 10), 1600 => to_unsigned(690, 10), 1601 => to_unsigned(578, 10), 1602 => to_unsigned(568, 10), 1603 => to_unsigned(618, 10), 1604 => to_unsigned(250, 10), 1605 => to_unsigned(336, 10), 1606 => to_unsigned(634, 10), 1607 => to_unsigned(974, 10), 1608 => to_unsigned(235, 10), 1609 => to_unsigned(1007, 10), 1610 => to_unsigned(953, 10), 1611 => to_unsigned(756, 10), 1612 => to_unsigned(396, 10), 1613 => to_unsigned(168, 10), 1614 => to_unsigned(755, 10), 1615 => to_unsigned(489, 10), 1616 => to_unsigned(825, 10), 1617 => to_unsigned(338, 10), 1618 => to_unsigned(915, 10), 1619 => to_unsigned(194, 10), 1620 => to_unsigned(324, 10), 1621 => to_unsigned(983, 10), 1622 => to_unsigned(406, 10), 1623 => to_unsigned(41, 10), 1624 => to_unsigned(105, 10), 1625 => to_unsigned(188, 10), 1626 => to_unsigned(140, 10), 1627 => to_unsigned(511, 10), 1628 => to_unsigned(873, 10), 1629 => to_unsigned(615, 10), 1630 => to_unsigned(833, 10), 1631 => to_unsigned(18, 10), 1632 => to_unsigned(722, 10), 1633 => to_unsigned(131, 10), 1634 => to_unsigned(575, 10), 1635 => to_unsigned(661, 10), 1636 => to_unsigned(423, 10), 1637 => to_unsigned(520, 10), 1638 => to_unsigned(833, 10), 1639 => to_unsigned(373, 10), 1640 => to_unsigned(741, 10), 1641 => to_unsigned(553, 10), 1642 => to_unsigned(160, 10), 1643 => to_unsigned(950, 10), 1644 => to_unsigned(560, 10), 1645 => to_unsigned(402, 10), 1646 => to_unsigned(799, 10), 1647 => to_unsigned(610, 10), 1648 => to_unsigned(868, 10), 1649 => to_unsigned(887, 10), 1650 => to_unsigned(435, 10), 1651 => to_unsigned(503, 10), 1652 => to_unsigned(700, 10), 1653 => to_unsigned(866, 10), 1654 => to_unsigned(783, 10), 1655 => to_unsigned(276, 10), 1656 => to_unsigned(145, 10), 1657 => to_unsigned(679, 10), 1658 => to_unsigned(322, 10), 1659 => to_unsigned(973, 10), 1660 => to_unsigned(62, 10), 1661 => to_unsigned(612, 10), 1662 => to_unsigned(12, 10), 1663 => to_unsigned(943, 10), 1664 => to_unsigned(878, 10), 1665 => to_unsigned(930, 10), 1666 => to_unsigned(369, 10), 1667 => to_unsigned(605, 10), 1668 => to_unsigned(887, 10), 1669 => to_unsigned(403, 10), 1670 => to_unsigned(304, 10), 1671 => to_unsigned(265, 10), 1672 => to_unsigned(923, 10), 1673 => to_unsigned(325, 10), 1674 => to_unsigned(421, 10), 1675 => to_unsigned(599, 10), 1676 => to_unsigned(574, 10), 1677 => to_unsigned(510, 10), 1678 => to_unsigned(755, 10), 1679 => to_unsigned(536, 10), 1680 => to_unsigned(57, 10), 1681 => to_unsigned(522, 10), 1682 => to_unsigned(1016, 10), 1683 => to_unsigned(586, 10), 1684 => to_unsigned(392, 10), 1685 => to_unsigned(771, 10), 1686 => to_unsigned(720, 10), 1687 => to_unsigned(28, 10), 1688 => to_unsigned(565, 10), 1689 => to_unsigned(1004, 10), 1690 => to_unsigned(107, 10), 1691 => to_unsigned(806, 10), 1692 => to_unsigned(409, 10), 1693 => to_unsigned(420, 10), 1694 => to_unsigned(8, 10), 1695 => to_unsigned(124, 10), 1696 => to_unsigned(312, 10), 1697 => to_unsigned(350, 10), 1698 => to_unsigned(758, 10), 1699 => to_unsigned(10, 10), 1700 => to_unsigned(932, 10), 1701 => to_unsigned(341, 10), 1702 => to_unsigned(807, 10), 1703 => to_unsigned(412, 10), 1704 => to_unsigned(365, 10), 1705 => to_unsigned(817, 10), 1706 => to_unsigned(99, 10), 1707 => to_unsigned(161, 10), 1708 => to_unsigned(624, 10), 1709 => to_unsigned(1019, 10), 1710 => to_unsigned(939, 10), 1711 => to_unsigned(603, 10), 1712 => to_unsigned(639, 10), 1713 => to_unsigned(28, 10), 1714 => to_unsigned(833, 10), 1715 => to_unsigned(350, 10), 1716 => to_unsigned(942, 10), 1717 => to_unsigned(542, 10), 1718 => to_unsigned(240, 10), 1719 => to_unsigned(974, 10), 1720 => to_unsigned(705, 10), 1721 => to_unsigned(499, 10), 1722 => to_unsigned(928, 10), 1723 => to_unsigned(494, 10), 1724 => to_unsigned(522, 10), 1725 => to_unsigned(121, 10), 1726 => to_unsigned(602, 10), 1727 => to_unsigned(872, 10), 1728 => to_unsigned(653, 10), 1729 => to_unsigned(138, 10), 1730 => to_unsigned(700, 10), 1731 => to_unsigned(957, 10), 1732 => to_unsigned(405, 10), 1733 => to_unsigned(432, 10), 1734 => to_unsigned(343, 10), 1735 => to_unsigned(76, 10), 1736 => to_unsigned(291, 10), 1737 => to_unsigned(365, 10), 1738 => to_unsigned(989, 10), 1739 => to_unsigned(16, 10), 1740 => to_unsigned(245, 10), 1741 => to_unsigned(107, 10), 1742 => to_unsigned(777, 10), 1743 => to_unsigned(1021, 10), 1744 => to_unsigned(1004, 10), 1745 => to_unsigned(652, 10), 1746 => to_unsigned(127, 10), 1747 => to_unsigned(782, 10), 1748 => to_unsigned(556, 10), 1749 => to_unsigned(397, 10), 1750 => to_unsigned(348, 10), 1751 => to_unsigned(906, 10), 1752 => to_unsigned(410, 10), 1753 => to_unsigned(988, 10), 1754 => to_unsigned(830, 10), 1755 => to_unsigned(256, 10), 1756 => to_unsigned(114, 10), 1757 => to_unsigned(219, 10), 1758 => to_unsigned(883, 10), 1759 => to_unsigned(711, 10), 1760 => to_unsigned(173, 10), 1761 => to_unsigned(819, 10), 1762 => to_unsigned(52, 10), 1763 => to_unsigned(247, 10), 1764 => to_unsigned(197, 10), 1765 => to_unsigned(395, 10), 1766 => to_unsigned(833, 10), 1767 => to_unsigned(306, 10), 1768 => to_unsigned(340, 10), 1769 => to_unsigned(223, 10), 1770 => to_unsigned(797, 10), 1771 => to_unsigned(445, 10), 1772 => to_unsigned(136, 10), 1773 => to_unsigned(608, 10), 1774 => to_unsigned(283, 10), 1775 => to_unsigned(125, 10), 1776 => to_unsigned(761, 10), 1777 => to_unsigned(32, 10), 1778 => to_unsigned(557, 10), 1779 => to_unsigned(174, 10), 1780 => to_unsigned(734, 10), 1781 => to_unsigned(565, 10), 1782 => to_unsigned(714, 10), 1783 => to_unsigned(948, 10), 1784 => to_unsigned(347, 10), 1785 => to_unsigned(47, 10), 1786 => to_unsigned(68, 10), 1787 => to_unsigned(394, 10), 1788 => to_unsigned(752, 10), 1789 => to_unsigned(728, 10), 1790 => to_unsigned(43, 10), 1791 => to_unsigned(612, 10), 1792 => to_unsigned(384, 10), 1793 => to_unsigned(181, 10), 1794 => to_unsigned(537, 10), 1795 => to_unsigned(132, 10), 1796 => to_unsigned(390, 10), 1797 => to_unsigned(26, 10), 1798 => to_unsigned(517, 10), 1799 => to_unsigned(479, 10), 1800 => to_unsigned(1001, 10), 1801 => to_unsigned(944, 10), 1802 => to_unsigned(180, 10), 1803 => to_unsigned(554, 10), 1804 => to_unsigned(442, 10), 1805 => to_unsigned(912, 10), 1806 => to_unsigned(954, 10), 1807 => to_unsigned(914, 10), 1808 => to_unsigned(191, 10), 1809 => to_unsigned(830, 10), 1810 => to_unsigned(777, 10), 1811 => to_unsigned(616, 10), 1812 => to_unsigned(809, 10), 1813 => to_unsigned(604, 10), 1814 => to_unsigned(2, 10), 1815 => to_unsigned(94, 10), 1816 => to_unsigned(90, 10), 1817 => to_unsigned(456, 10), 1818 => to_unsigned(149, 10), 1819 => to_unsigned(858, 10), 1820 => to_unsigned(795, 10), 1821 => to_unsigned(679, 10), 1822 => to_unsigned(940, 10), 1823 => to_unsigned(377, 10), 1824 => to_unsigned(382, 10), 1825 => to_unsigned(255, 10), 1826 => to_unsigned(391, 10), 1827 => to_unsigned(365, 10), 1828 => to_unsigned(446, 10), 1829 => to_unsigned(361, 10), 1830 => to_unsigned(963, 10), 1831 => to_unsigned(237, 10), 1832 => to_unsigned(740, 10), 1833 => to_unsigned(35, 10), 1834 => to_unsigned(24, 10), 1835 => to_unsigned(913, 10), 1836 => to_unsigned(425, 10), 1837 => to_unsigned(537, 10), 1838 => to_unsigned(986, 10), 1839 => to_unsigned(761, 10), 1840 => to_unsigned(995, 10), 1841 => to_unsigned(470, 10), 1842 => to_unsigned(272, 10), 1843 => to_unsigned(779, 10), 1844 => to_unsigned(215, 10), 1845 => to_unsigned(180, 10), 1846 => to_unsigned(0, 10), 1847 => to_unsigned(690, 10), 1848 => to_unsigned(86, 10), 1849 => to_unsigned(77, 10), 1850 => to_unsigned(816, 10), 1851 => to_unsigned(770, 10), 1852 => to_unsigned(419, 10), 1853 => to_unsigned(321, 10), 1854 => to_unsigned(128, 10), 1855 => to_unsigned(941, 10), 1856 => to_unsigned(533, 10), 1857 => to_unsigned(10, 10), 1858 => to_unsigned(70, 10), 1859 => to_unsigned(478, 10), 1860 => to_unsigned(692, 10), 1861 => to_unsigned(228, 10), 1862 => to_unsigned(119, 10), 1863 => to_unsigned(865, 10), 1864 => to_unsigned(811, 10), 1865 => to_unsigned(69, 10), 1866 => to_unsigned(847, 10), 1867 => to_unsigned(162, 10), 1868 => to_unsigned(1008, 10), 1869 => to_unsigned(905, 10), 1870 => to_unsigned(748, 10), 1871 => to_unsigned(874, 10), 1872 => to_unsigned(156, 10), 1873 => to_unsigned(747, 10), 1874 => to_unsigned(1006, 10), 1875 => to_unsigned(425, 10), 1876 => to_unsigned(613, 10), 1877 => to_unsigned(854, 10), 1878 => to_unsigned(771, 10), 1879 => to_unsigned(130, 10), 1880 => to_unsigned(344, 10), 1881 => to_unsigned(70, 10), 1882 => to_unsigned(773, 10), 1883 => to_unsigned(311, 10), 1884 => to_unsigned(173, 10), 1885 => to_unsigned(123, 10), 1886 => to_unsigned(365, 10), 1887 => to_unsigned(66, 10), 1888 => to_unsigned(462, 10), 1889 => to_unsigned(646, 10), 1890 => to_unsigned(68, 10), 1891 => to_unsigned(653, 10), 1892 => to_unsigned(914, 10), 1893 => to_unsigned(674, 10), 1894 => to_unsigned(240, 10), 1895 => to_unsigned(180, 10), 1896 => to_unsigned(171, 10), 1897 => to_unsigned(171, 10), 1898 => to_unsigned(854, 10), 1899 => to_unsigned(617, 10), 1900 => to_unsigned(223, 10), 1901 => to_unsigned(996, 10), 1902 => to_unsigned(29, 10), 1903 => to_unsigned(188, 10), 1904 => to_unsigned(773, 10), 1905 => to_unsigned(480, 10), 1906 => to_unsigned(539, 10), 1907 => to_unsigned(550, 10), 1908 => to_unsigned(38, 10), 1909 => to_unsigned(277, 10), 1910 => to_unsigned(573, 10), 1911 => to_unsigned(923, 10), 1912 => to_unsigned(538, 10), 1913 => to_unsigned(923, 10), 1914 => to_unsigned(796, 10), 1915 => to_unsigned(629, 10), 1916 => to_unsigned(790, 10), 1917 => to_unsigned(620, 10), 1918 => to_unsigned(985, 10), 1919 => to_unsigned(891, 10), 1920 => to_unsigned(993, 10), 1921 => to_unsigned(501, 10), 1922 => to_unsigned(966, 10), 1923 => to_unsigned(476, 10), 1924 => to_unsigned(334, 10), 1925 => to_unsigned(370, 10), 1926 => to_unsigned(8, 10), 1927 => to_unsigned(551, 10), 1928 => to_unsigned(694, 10), 1929 => to_unsigned(309, 10), 1930 => to_unsigned(462, 10), 1931 => to_unsigned(119, 10), 1932 => to_unsigned(522, 10), 1933 => to_unsigned(419, 10), 1934 => to_unsigned(403, 10), 1935 => to_unsigned(929, 10), 1936 => to_unsigned(655, 10), 1937 => to_unsigned(1022, 10), 1938 => to_unsigned(720, 10), 1939 => to_unsigned(565, 10), 1940 => to_unsigned(105, 10), 1941 => to_unsigned(838, 10), 1942 => to_unsigned(684, 10), 1943 => to_unsigned(272, 10), 1944 => to_unsigned(145, 10), 1945 => to_unsigned(876, 10), 1946 => to_unsigned(954, 10), 1947 => to_unsigned(605, 10), 1948 => to_unsigned(408, 10), 1949 => to_unsigned(159, 10), 1950 => to_unsigned(227, 10), 1951 => to_unsigned(484, 10), 1952 => to_unsigned(240, 10), 1953 => to_unsigned(14, 10), 1954 => to_unsigned(330, 10), 1955 => to_unsigned(412, 10), 1956 => to_unsigned(263, 10), 1957 => to_unsigned(952, 10), 1958 => to_unsigned(346, 10), 1959 => to_unsigned(318, 10), 1960 => to_unsigned(935, 10), 1961 => to_unsigned(541, 10), 1962 => to_unsigned(908, 10), 1963 => to_unsigned(356, 10), 1964 => to_unsigned(204, 10), 1965 => to_unsigned(868, 10), 1966 => to_unsigned(745, 10), 1967 => to_unsigned(193, 10), 1968 => to_unsigned(529, 10), 1969 => to_unsigned(995, 10), 1970 => to_unsigned(877, 10), 1971 => to_unsigned(801, 10), 1972 => to_unsigned(860, 10), 1973 => to_unsigned(372, 10), 1974 => to_unsigned(541, 10), 1975 => to_unsigned(569, 10), 1976 => to_unsigned(378, 10), 1977 => to_unsigned(216, 10), 1978 => to_unsigned(986, 10), 1979 => to_unsigned(929, 10), 1980 => to_unsigned(253, 10), 1981 => to_unsigned(241, 10), 1982 => to_unsigned(456, 10), 1983 => to_unsigned(937, 10), 1984 => to_unsigned(312, 10), 1985 => to_unsigned(597, 10), 1986 => to_unsigned(146, 10), 1987 => to_unsigned(55, 10), 1988 => to_unsigned(840, 10), 1989 => to_unsigned(819, 10), 1990 => to_unsigned(913, 10), 1991 => to_unsigned(531, 10), 1992 => to_unsigned(706, 10), 1993 => to_unsigned(551, 10), 1994 => to_unsigned(571, 10), 1995 => to_unsigned(19, 10), 1996 => to_unsigned(933, 10), 1997 => to_unsigned(180, 10), 1998 => to_unsigned(653, 10), 1999 => to_unsigned(539, 10), 2000 => to_unsigned(633, 10), 2001 => to_unsigned(254, 10), 2002 => to_unsigned(848, 10), 2003 => to_unsigned(785, 10), 2004 => to_unsigned(78, 10), 2005 => to_unsigned(1021, 10), 2006 => to_unsigned(663, 10), 2007 => to_unsigned(922, 10), 2008 => to_unsigned(988, 10), 2009 => to_unsigned(407, 10), 2010 => to_unsigned(356, 10), 2011 => to_unsigned(513, 10), 2012 => to_unsigned(956, 10), 2013 => to_unsigned(471, 10), 2014 => to_unsigned(845, 10), 2015 => to_unsigned(103, 10), 2016 => to_unsigned(971, 10), 2017 => to_unsigned(14, 10), 2018 => to_unsigned(513, 10), 2019 => to_unsigned(689, 10), 2020 => to_unsigned(17, 10), 2021 => to_unsigned(298, 10), 2022 => to_unsigned(137, 10), 2023 => to_unsigned(272, 10), 2024 => to_unsigned(907, 10), 2025 => to_unsigned(331, 10), 2026 => to_unsigned(678, 10), 2027 => to_unsigned(646, 10), 2028 => to_unsigned(453, 10), 2029 => to_unsigned(824, 10), 2030 => to_unsigned(796, 10), 2031 => to_unsigned(490, 10), 2032 => to_unsigned(457, 10), 2033 => to_unsigned(814, 10), 2034 => to_unsigned(938, 10), 2035 => to_unsigned(313, 10), 2036 => to_unsigned(121, 10), 2037 => to_unsigned(167, 10), 2038 => to_unsigned(110, 10), 2039 => to_unsigned(1019, 10), 2040 => to_unsigned(619, 10), 2041 => to_unsigned(932, 10), 2042 => to_unsigned(393, 10), 2043 => to_unsigned(516, 10), 2044 => to_unsigned(983, 10), 2045 => to_unsigned(871, 10), 2046 => to_unsigned(365, 10), 2047 => to_unsigned(736, 10)),
            3 => (0 => to_unsigned(245, 10), 1 => to_unsigned(909, 10), 2 => to_unsigned(239, 10), 3 => to_unsigned(288, 10), 4 => to_unsigned(67, 10), 5 => to_unsigned(497, 10), 6 => to_unsigned(175, 10), 7 => to_unsigned(861, 10), 8 => to_unsigned(977, 10), 9 => to_unsigned(920, 10), 10 => to_unsigned(72, 10), 11 => to_unsigned(644, 10), 12 => to_unsigned(263, 10), 13 => to_unsigned(478, 10), 14 => to_unsigned(19, 10), 15 => to_unsigned(459, 10), 16 => to_unsigned(260, 10), 17 => to_unsigned(707, 10), 18 => to_unsigned(949, 10), 19 => to_unsigned(617, 10), 20 => to_unsigned(706, 10), 21 => to_unsigned(9, 10), 22 => to_unsigned(721, 10), 23 => to_unsigned(668, 10), 24 => to_unsigned(1007, 10), 25 => to_unsigned(736, 10), 26 => to_unsigned(94, 10), 27 => to_unsigned(547, 10), 28 => to_unsigned(452, 10), 29 => to_unsigned(276, 10), 30 => to_unsigned(509, 10), 31 => to_unsigned(175, 10), 32 => to_unsigned(996, 10), 33 => to_unsigned(862, 10), 34 => to_unsigned(234, 10), 35 => to_unsigned(925, 10), 36 => to_unsigned(548, 10), 37 => to_unsigned(187, 10), 38 => to_unsigned(932, 10), 39 => to_unsigned(88, 10), 40 => to_unsigned(905, 10), 41 => to_unsigned(206, 10), 42 => to_unsigned(51, 10), 43 => to_unsigned(388, 10), 44 => to_unsigned(463, 10), 45 => to_unsigned(760, 10), 46 => to_unsigned(137, 10), 47 => to_unsigned(479, 10), 48 => to_unsigned(181, 10), 49 => to_unsigned(751, 10), 50 => to_unsigned(859, 10), 51 => to_unsigned(787, 10), 52 => to_unsigned(293, 10), 53 => to_unsigned(875, 10), 54 => to_unsigned(467, 10), 55 => to_unsigned(17, 10), 56 => to_unsigned(138, 10), 57 => to_unsigned(745, 10), 58 => to_unsigned(315, 10), 59 => to_unsigned(398, 10), 60 => to_unsigned(60, 10), 61 => to_unsigned(816, 10), 62 => to_unsigned(255, 10), 63 => to_unsigned(27, 10), 64 => to_unsigned(466, 10), 65 => to_unsigned(261, 10), 66 => to_unsigned(173, 10), 67 => to_unsigned(132, 10), 68 => to_unsigned(936, 10), 69 => to_unsigned(482, 10), 70 => to_unsigned(453, 10), 71 => to_unsigned(393, 10), 72 => to_unsigned(33, 10), 73 => to_unsigned(84, 10), 74 => to_unsigned(296, 10), 75 => to_unsigned(343, 10), 76 => to_unsigned(427, 10), 77 => to_unsigned(436, 10), 78 => to_unsigned(719, 10), 79 => to_unsigned(519, 10), 80 => to_unsigned(373, 10), 81 => to_unsigned(685, 10), 82 => to_unsigned(166, 10), 83 => to_unsigned(816, 10), 84 => to_unsigned(920, 10), 85 => to_unsigned(215, 10), 86 => to_unsigned(965, 10), 87 => to_unsigned(381, 10), 88 => to_unsigned(588, 10), 89 => to_unsigned(212, 10), 90 => to_unsigned(766, 10), 91 => to_unsigned(780, 10), 92 => to_unsigned(348, 10), 93 => to_unsigned(547, 10), 94 => to_unsigned(469, 10), 95 => to_unsigned(901, 10), 96 => to_unsigned(294, 10), 97 => to_unsigned(948, 10), 98 => to_unsigned(81, 10), 99 => to_unsigned(183, 10), 100 => to_unsigned(252, 10), 101 => to_unsigned(500, 10), 102 => to_unsigned(321, 10), 103 => to_unsigned(179, 10), 104 => to_unsigned(780, 10), 105 => to_unsigned(8, 10), 106 => to_unsigned(707, 10), 107 => to_unsigned(573, 10), 108 => to_unsigned(676, 10), 109 => to_unsigned(141, 10), 110 => to_unsigned(727, 10), 111 => to_unsigned(327, 10), 112 => to_unsigned(423, 10), 113 => to_unsigned(53, 10), 114 => to_unsigned(606, 10), 115 => to_unsigned(804, 10), 116 => to_unsigned(942, 10), 117 => to_unsigned(968, 10), 118 => to_unsigned(842, 10), 119 => to_unsigned(517, 10), 120 => to_unsigned(39, 10), 121 => to_unsigned(642, 10), 122 => to_unsigned(275, 10), 123 => to_unsigned(569, 10), 124 => to_unsigned(515, 10), 125 => to_unsigned(506, 10), 126 => to_unsigned(951, 10), 127 => to_unsigned(600, 10), 128 => to_unsigned(330, 10), 129 => to_unsigned(342, 10), 130 => to_unsigned(513, 10), 131 => to_unsigned(403, 10), 132 => to_unsigned(284, 10), 133 => to_unsigned(379, 10), 134 => to_unsigned(882, 10), 135 => to_unsigned(157, 10), 136 => to_unsigned(865, 10), 137 => to_unsigned(22, 10), 138 => to_unsigned(903, 10), 139 => to_unsigned(136, 10), 140 => to_unsigned(878, 10), 141 => to_unsigned(624, 10), 142 => to_unsigned(681, 10), 143 => to_unsigned(989, 10), 144 => to_unsigned(723, 10), 145 => to_unsigned(22, 10), 146 => to_unsigned(745, 10), 147 => to_unsigned(840, 10), 148 => to_unsigned(689, 10), 149 => to_unsigned(583, 10), 150 => to_unsigned(64, 10), 151 => to_unsigned(28, 10), 152 => to_unsigned(197, 10), 153 => to_unsigned(403, 10), 154 => to_unsigned(241, 10), 155 => to_unsigned(263, 10), 156 => to_unsigned(572, 10), 157 => to_unsigned(699, 10), 158 => to_unsigned(806, 10), 159 => to_unsigned(360, 10), 160 => to_unsigned(985, 10), 161 => to_unsigned(645, 10), 162 => to_unsigned(803, 10), 163 => to_unsigned(216, 10), 164 => to_unsigned(118, 10), 165 => to_unsigned(522, 10), 166 => to_unsigned(828, 10), 167 => to_unsigned(107, 10), 168 => to_unsigned(201, 10), 169 => to_unsigned(932, 10), 170 => to_unsigned(698, 10), 171 => to_unsigned(789, 10), 172 => to_unsigned(272, 10), 173 => to_unsigned(45, 10), 174 => to_unsigned(627, 10), 175 => to_unsigned(996, 10), 176 => to_unsigned(208, 10), 177 => to_unsigned(362, 10), 178 => to_unsigned(902, 10), 179 => to_unsigned(437, 10), 180 => to_unsigned(681, 10), 181 => to_unsigned(793, 10), 182 => to_unsigned(244, 10), 183 => to_unsigned(418, 10), 184 => to_unsigned(67, 10), 185 => to_unsigned(251, 10), 186 => to_unsigned(662, 10), 187 => to_unsigned(93, 10), 188 => to_unsigned(692, 10), 189 => to_unsigned(408, 10), 190 => to_unsigned(945, 10), 191 => to_unsigned(801, 10), 192 => to_unsigned(995, 10), 193 => to_unsigned(344, 10), 194 => to_unsigned(294, 10), 195 => to_unsigned(75, 10), 196 => to_unsigned(702, 10), 197 => to_unsigned(618, 10), 198 => to_unsigned(931, 10), 199 => to_unsigned(728, 10), 200 => to_unsigned(953, 10), 201 => to_unsigned(753, 10), 202 => to_unsigned(519, 10), 203 => to_unsigned(100, 10), 204 => to_unsigned(651, 10), 205 => to_unsigned(128, 10), 206 => to_unsigned(420, 10), 207 => to_unsigned(5, 10), 208 => to_unsigned(9, 10), 209 => to_unsigned(889, 10), 210 => to_unsigned(581, 10), 211 => to_unsigned(682, 10), 212 => to_unsigned(270, 10), 213 => to_unsigned(86, 10), 214 => to_unsigned(294, 10), 215 => to_unsigned(289, 10), 216 => to_unsigned(35, 10), 217 => to_unsigned(648, 10), 218 => to_unsigned(479, 10), 219 => to_unsigned(2, 10), 220 => to_unsigned(951, 10), 221 => to_unsigned(36, 10), 222 => to_unsigned(956, 10), 223 => to_unsigned(20, 10), 224 => to_unsigned(915, 10), 225 => to_unsigned(109, 10), 226 => to_unsigned(670, 10), 227 => to_unsigned(329, 10), 228 => to_unsigned(916, 10), 229 => to_unsigned(161, 10), 230 => to_unsigned(871, 10), 231 => to_unsigned(994, 10), 232 => to_unsigned(986, 10), 233 => to_unsigned(594, 10), 234 => to_unsigned(740, 10), 235 => to_unsigned(178, 10), 236 => to_unsigned(291, 10), 237 => to_unsigned(190, 10), 238 => to_unsigned(745, 10), 239 => to_unsigned(714, 10), 240 => to_unsigned(587, 10), 241 => to_unsigned(581, 10), 242 => to_unsigned(826, 10), 243 => to_unsigned(760, 10), 244 => to_unsigned(732, 10), 245 => to_unsigned(356, 10), 246 => to_unsigned(459, 10), 247 => to_unsigned(870, 10), 248 => to_unsigned(438, 10), 249 => to_unsigned(464, 10), 250 => to_unsigned(675, 10), 251 => to_unsigned(340, 10), 252 => to_unsigned(866, 10), 253 => to_unsigned(844, 10), 254 => to_unsigned(387, 10), 255 => to_unsigned(701, 10), 256 => to_unsigned(253, 10), 257 => to_unsigned(166, 10), 258 => to_unsigned(1001, 10), 259 => to_unsigned(636, 10), 260 => to_unsigned(583, 10), 261 => to_unsigned(495, 10), 262 => to_unsigned(779, 10), 263 => to_unsigned(213, 10), 264 => to_unsigned(885, 10), 265 => to_unsigned(597, 10), 266 => to_unsigned(718, 10), 267 => to_unsigned(139, 10), 268 => to_unsigned(257, 10), 269 => to_unsigned(652, 10), 270 => to_unsigned(554, 10), 271 => to_unsigned(791, 10), 272 => to_unsigned(197, 10), 273 => to_unsigned(944, 10), 274 => to_unsigned(879, 10), 275 => to_unsigned(549, 10), 276 => to_unsigned(140, 10), 277 => to_unsigned(563, 10), 278 => to_unsigned(338, 10), 279 => to_unsigned(536, 10), 280 => to_unsigned(20, 10), 281 => to_unsigned(528, 10), 282 => to_unsigned(15, 10), 283 => to_unsigned(654, 10), 284 => to_unsigned(869, 10), 285 => to_unsigned(164, 10), 286 => to_unsigned(380, 10), 287 => to_unsigned(343, 10), 288 => to_unsigned(675, 10), 289 => to_unsigned(660, 10), 290 => to_unsigned(310, 10), 291 => to_unsigned(106, 10), 292 => to_unsigned(255, 10), 293 => to_unsigned(247, 10), 294 => to_unsigned(906, 10), 295 => to_unsigned(199, 10), 296 => to_unsigned(189, 10), 297 => to_unsigned(116, 10), 298 => to_unsigned(935, 10), 299 => to_unsigned(405, 10), 300 => to_unsigned(449, 10), 301 => to_unsigned(884, 10), 302 => to_unsigned(266, 10), 303 => to_unsigned(605, 10), 304 => to_unsigned(155, 10), 305 => to_unsigned(436, 10), 306 => to_unsigned(611, 10), 307 => to_unsigned(365, 10), 308 => to_unsigned(544, 10), 309 => to_unsigned(135, 10), 310 => to_unsigned(422, 10), 311 => to_unsigned(633, 10), 312 => to_unsigned(174, 10), 313 => to_unsigned(566, 10), 314 => to_unsigned(406, 10), 315 => to_unsigned(232, 10), 316 => to_unsigned(788, 10), 317 => to_unsigned(68, 10), 318 => to_unsigned(766, 10), 319 => to_unsigned(982, 10), 320 => to_unsigned(868, 10), 321 => to_unsigned(160, 10), 322 => to_unsigned(576, 10), 323 => to_unsigned(851, 10), 324 => to_unsigned(656, 10), 325 => to_unsigned(299, 10), 326 => to_unsigned(457, 10), 327 => to_unsigned(323, 10), 328 => to_unsigned(80, 10), 329 => to_unsigned(497, 10), 330 => to_unsigned(502, 10), 331 => to_unsigned(719, 10), 332 => to_unsigned(721, 10), 333 => to_unsigned(844, 10), 334 => to_unsigned(546, 10), 335 => to_unsigned(811, 10), 336 => to_unsigned(312, 10), 337 => to_unsigned(920, 10), 338 => to_unsigned(832, 10), 339 => to_unsigned(688, 10), 340 => to_unsigned(928, 10), 341 => to_unsigned(392, 10), 342 => to_unsigned(611, 10), 343 => to_unsigned(143, 10), 344 => to_unsigned(1008, 10), 345 => to_unsigned(930, 10), 346 => to_unsigned(506, 10), 347 => to_unsigned(485, 10), 348 => to_unsigned(759, 10), 349 => to_unsigned(792, 10), 350 => to_unsigned(596, 10), 351 => to_unsigned(428, 10), 352 => to_unsigned(599, 10), 353 => to_unsigned(559, 10), 354 => to_unsigned(978, 10), 355 => to_unsigned(261, 10), 356 => to_unsigned(244, 10), 357 => to_unsigned(309, 10), 358 => to_unsigned(66, 10), 359 => to_unsigned(1004, 10), 360 => to_unsigned(112, 10), 361 => to_unsigned(692, 10), 362 => to_unsigned(917, 10), 363 => to_unsigned(740, 10), 364 => to_unsigned(859, 10), 365 => to_unsigned(843, 10), 366 => to_unsigned(588, 10), 367 => to_unsigned(879, 10), 368 => to_unsigned(887, 10), 369 => to_unsigned(633, 10), 370 => to_unsigned(702, 10), 371 => to_unsigned(488, 10), 372 => to_unsigned(174, 10), 373 => to_unsigned(781, 10), 374 => to_unsigned(538, 10), 375 => to_unsigned(299, 10), 376 => to_unsigned(481, 10), 377 => to_unsigned(681, 10), 378 => to_unsigned(140, 10), 379 => to_unsigned(38, 10), 380 => to_unsigned(18, 10), 381 => to_unsigned(169, 10), 382 => to_unsigned(667, 10), 383 => to_unsigned(389, 10), 384 => to_unsigned(828, 10), 385 => to_unsigned(10, 10), 386 => to_unsigned(223, 10), 387 => to_unsigned(961, 10), 388 => to_unsigned(282, 10), 389 => to_unsigned(661, 10), 390 => to_unsigned(151, 10), 391 => to_unsigned(437, 10), 392 => to_unsigned(85, 10), 393 => to_unsigned(1023, 10), 394 => to_unsigned(463, 10), 395 => to_unsigned(48, 10), 396 => to_unsigned(932, 10), 397 => to_unsigned(129, 10), 398 => to_unsigned(823, 10), 399 => to_unsigned(342, 10), 400 => to_unsigned(967, 10), 401 => to_unsigned(701, 10), 402 => to_unsigned(686, 10), 403 => to_unsigned(497, 10), 404 => to_unsigned(585, 10), 405 => to_unsigned(712, 10), 406 => to_unsigned(12, 10), 407 => to_unsigned(956, 10), 408 => to_unsigned(603, 10), 409 => to_unsigned(259, 10), 410 => to_unsigned(917, 10), 411 => to_unsigned(77, 10), 412 => to_unsigned(181, 10), 413 => to_unsigned(422, 10), 414 => to_unsigned(228, 10), 415 => to_unsigned(570, 10), 416 => to_unsigned(692, 10), 417 => to_unsigned(739, 10), 418 => to_unsigned(65, 10), 419 => to_unsigned(107, 10), 420 => to_unsigned(948, 10), 421 => to_unsigned(336, 10), 422 => to_unsigned(714, 10), 423 => to_unsigned(13, 10), 424 => to_unsigned(520, 10), 425 => to_unsigned(370, 10), 426 => to_unsigned(837, 10), 427 => to_unsigned(232, 10), 428 => to_unsigned(54, 10), 429 => to_unsigned(467, 10), 430 => to_unsigned(1009, 10), 431 => to_unsigned(751, 10), 432 => to_unsigned(891, 10), 433 => to_unsigned(178, 10), 434 => to_unsigned(930, 10), 435 => to_unsigned(735, 10), 436 => to_unsigned(294, 10), 437 => to_unsigned(850, 10), 438 => to_unsigned(966, 10), 439 => to_unsigned(875, 10), 440 => to_unsigned(654, 10), 441 => to_unsigned(159, 10), 442 => to_unsigned(758, 10), 443 => to_unsigned(368, 10), 444 => to_unsigned(428, 10), 445 => to_unsigned(160, 10), 446 => to_unsigned(31, 10), 447 => to_unsigned(593, 10), 448 => to_unsigned(832, 10), 449 => to_unsigned(379, 10), 450 => to_unsigned(660, 10), 451 => to_unsigned(266, 10), 452 => to_unsigned(338, 10), 453 => to_unsigned(931, 10), 454 => to_unsigned(223, 10), 455 => to_unsigned(950, 10), 456 => to_unsigned(116, 10), 457 => to_unsigned(541, 10), 458 => to_unsigned(736, 10), 459 => to_unsigned(940, 10), 460 => to_unsigned(142, 10), 461 => to_unsigned(464, 10), 462 => to_unsigned(160, 10), 463 => to_unsigned(476, 10), 464 => to_unsigned(950, 10), 465 => to_unsigned(241, 10), 466 => to_unsigned(206, 10), 467 => to_unsigned(935, 10), 468 => to_unsigned(244, 10), 469 => to_unsigned(691, 10), 470 => to_unsigned(57, 10), 471 => to_unsigned(920, 10), 472 => to_unsigned(623, 10), 473 => to_unsigned(400, 10), 474 => to_unsigned(757, 10), 475 => to_unsigned(362, 10), 476 => to_unsigned(405, 10), 477 => to_unsigned(1005, 10), 478 => to_unsigned(779, 10), 479 => to_unsigned(37, 10), 480 => to_unsigned(162, 10), 481 => to_unsigned(545, 10), 482 => to_unsigned(278, 10), 483 => to_unsigned(102, 10), 484 => to_unsigned(528, 10), 485 => to_unsigned(629, 10), 486 => to_unsigned(292, 10), 487 => to_unsigned(704, 10), 488 => to_unsigned(410, 10), 489 => to_unsigned(77, 10), 490 => to_unsigned(857, 10), 491 => to_unsigned(766, 10), 492 => to_unsigned(590, 10), 493 => to_unsigned(927, 10), 494 => to_unsigned(800, 10), 495 => to_unsigned(537, 10), 496 => to_unsigned(496, 10), 497 => to_unsigned(756, 10), 498 => to_unsigned(135, 10), 499 => to_unsigned(575, 10), 500 => to_unsigned(460, 10), 501 => to_unsigned(144, 10), 502 => to_unsigned(296, 10), 503 => to_unsigned(517, 10), 504 => to_unsigned(627, 10), 505 => to_unsigned(169, 10), 506 => to_unsigned(685, 10), 507 => to_unsigned(469, 10), 508 => to_unsigned(282, 10), 509 => to_unsigned(329, 10), 510 => to_unsigned(765, 10), 511 => to_unsigned(694, 10), 512 => to_unsigned(840, 10), 513 => to_unsigned(837, 10), 514 => to_unsigned(732, 10), 515 => to_unsigned(530, 10), 516 => to_unsigned(668, 10), 517 => to_unsigned(292, 10), 518 => to_unsigned(555, 10), 519 => to_unsigned(602, 10), 520 => to_unsigned(4, 10), 521 => to_unsigned(357, 10), 522 => to_unsigned(324, 10), 523 => to_unsigned(711, 10), 524 => to_unsigned(312, 10), 525 => to_unsigned(1012, 10), 526 => to_unsigned(706, 10), 527 => to_unsigned(906, 10), 528 => to_unsigned(617, 10), 529 => to_unsigned(231, 10), 530 => to_unsigned(93, 10), 531 => to_unsigned(698, 10), 532 => to_unsigned(648, 10), 533 => to_unsigned(1006, 10), 534 => to_unsigned(793, 10), 535 => to_unsigned(422, 10), 536 => to_unsigned(656, 10), 537 => to_unsigned(783, 10), 538 => to_unsigned(298, 10), 539 => to_unsigned(643, 10), 540 => to_unsigned(438, 10), 541 => to_unsigned(20, 10), 542 => to_unsigned(286, 10), 543 => to_unsigned(346, 10), 544 => to_unsigned(618, 10), 545 => to_unsigned(691, 10), 546 => to_unsigned(402, 10), 547 => to_unsigned(199, 10), 548 => to_unsigned(924, 10), 549 => to_unsigned(103, 10), 550 => to_unsigned(244, 10), 551 => to_unsigned(851, 10), 552 => to_unsigned(374, 10), 553 => to_unsigned(542, 10), 554 => to_unsigned(371, 10), 555 => to_unsigned(577, 10), 556 => to_unsigned(981, 10), 557 => to_unsigned(866, 10), 558 => to_unsigned(709, 10), 559 => to_unsigned(196, 10), 560 => to_unsigned(290, 10), 561 => to_unsigned(54, 10), 562 => to_unsigned(602, 10), 563 => to_unsigned(1004, 10), 564 => to_unsigned(489, 10), 565 => to_unsigned(433, 10), 566 => to_unsigned(23, 10), 567 => to_unsigned(871, 10), 568 => to_unsigned(389, 10), 569 => to_unsigned(286, 10), 570 => to_unsigned(750, 10), 571 => to_unsigned(664, 10), 572 => to_unsigned(289, 10), 573 => to_unsigned(745, 10), 574 => to_unsigned(156, 10), 575 => to_unsigned(264, 10), 576 => to_unsigned(883, 10), 577 => to_unsigned(187, 10), 578 => to_unsigned(352, 10), 579 => to_unsigned(366, 10), 580 => to_unsigned(857, 10), 581 => to_unsigned(648, 10), 582 => to_unsigned(9, 10), 583 => to_unsigned(538, 10), 584 => to_unsigned(710, 10), 585 => to_unsigned(620, 10), 586 => to_unsigned(243, 10), 587 => to_unsigned(118, 10), 588 => to_unsigned(87, 10), 589 => to_unsigned(170, 10), 590 => to_unsigned(927, 10), 591 => to_unsigned(156, 10), 592 => to_unsigned(463, 10), 593 => to_unsigned(324, 10), 594 => to_unsigned(863, 10), 595 => to_unsigned(1016, 10), 596 => to_unsigned(725, 10), 597 => to_unsigned(77, 10), 598 => to_unsigned(664, 10), 599 => to_unsigned(958, 10), 600 => to_unsigned(60, 10), 601 => to_unsigned(608, 10), 602 => to_unsigned(984, 10), 603 => to_unsigned(196, 10), 604 => to_unsigned(410, 10), 605 => to_unsigned(612, 10), 606 => to_unsigned(53, 10), 607 => to_unsigned(761, 10), 608 => to_unsigned(757, 10), 609 => to_unsigned(403, 10), 610 => to_unsigned(834, 10), 611 => to_unsigned(496, 10), 612 => to_unsigned(597, 10), 613 => to_unsigned(709, 10), 614 => to_unsigned(926, 10), 615 => to_unsigned(900, 10), 616 => to_unsigned(538, 10), 617 => to_unsigned(734, 10), 618 => to_unsigned(911, 10), 619 => to_unsigned(267, 10), 620 => to_unsigned(729, 10), 621 => to_unsigned(678, 10), 622 => to_unsigned(437, 10), 623 => to_unsigned(494, 10), 624 => to_unsigned(362, 10), 625 => to_unsigned(634, 10), 626 => to_unsigned(73, 10), 627 => to_unsigned(280, 10), 628 => to_unsigned(857, 10), 629 => to_unsigned(822, 10), 630 => to_unsigned(195, 10), 631 => to_unsigned(489, 10), 632 => to_unsigned(694, 10), 633 => to_unsigned(346, 10), 634 => to_unsigned(930, 10), 635 => to_unsigned(791, 10), 636 => to_unsigned(95, 10), 637 => to_unsigned(962, 10), 638 => to_unsigned(968, 10), 639 => to_unsigned(75, 10), 640 => to_unsigned(749, 10), 641 => to_unsigned(482, 10), 642 => to_unsigned(739, 10), 643 => to_unsigned(585, 10), 644 => to_unsigned(825, 10), 645 => to_unsigned(954, 10), 646 => to_unsigned(205, 10), 647 => to_unsigned(553, 10), 648 => to_unsigned(999, 10), 649 => to_unsigned(959, 10), 650 => to_unsigned(491, 10), 651 => to_unsigned(142, 10), 652 => to_unsigned(135, 10), 653 => to_unsigned(975, 10), 654 => to_unsigned(163, 10), 655 => to_unsigned(54, 10), 656 => to_unsigned(413, 10), 657 => to_unsigned(379, 10), 658 => to_unsigned(301, 10), 659 => to_unsigned(66, 10), 660 => to_unsigned(824, 10), 661 => to_unsigned(274, 10), 662 => to_unsigned(745, 10), 663 => to_unsigned(224, 10), 664 => to_unsigned(203, 10), 665 => to_unsigned(160, 10), 666 => to_unsigned(61, 10), 667 => to_unsigned(308, 10), 668 => to_unsigned(262, 10), 669 => to_unsigned(626, 10), 670 => to_unsigned(489, 10), 671 => to_unsigned(649, 10), 672 => to_unsigned(1002, 10), 673 => to_unsigned(486, 10), 674 => to_unsigned(684, 10), 675 => to_unsigned(523, 10), 676 => to_unsigned(484, 10), 677 => to_unsigned(366, 10), 678 => to_unsigned(937, 10), 679 => to_unsigned(992, 10), 680 => to_unsigned(725, 10), 681 => to_unsigned(595, 10), 682 => to_unsigned(26, 10), 683 => to_unsigned(364, 10), 684 => to_unsigned(473, 10), 685 => to_unsigned(241, 10), 686 => to_unsigned(872, 10), 687 => to_unsigned(831, 10), 688 => to_unsigned(807, 10), 689 => to_unsigned(937, 10), 690 => to_unsigned(574, 10), 691 => to_unsigned(288, 10), 692 => to_unsigned(510, 10), 693 => to_unsigned(57, 10), 694 => to_unsigned(5, 10), 695 => to_unsigned(90, 10), 696 => to_unsigned(793, 10), 697 => to_unsigned(160, 10), 698 => to_unsigned(748, 10), 699 => to_unsigned(209, 10), 700 => to_unsigned(260, 10), 701 => to_unsigned(581, 10), 702 => to_unsigned(100, 10), 703 => to_unsigned(947, 10), 704 => to_unsigned(17, 10), 705 => to_unsigned(50, 10), 706 => to_unsigned(767, 10), 707 => to_unsigned(1011, 10), 708 => to_unsigned(268, 10), 709 => to_unsigned(12, 10), 710 => to_unsigned(641, 10), 711 => to_unsigned(818, 10), 712 => to_unsigned(741, 10), 713 => to_unsigned(312, 10), 714 => to_unsigned(370, 10), 715 => to_unsigned(384, 10), 716 => to_unsigned(727, 10), 717 => to_unsigned(774, 10), 718 => to_unsigned(778, 10), 719 => to_unsigned(1007, 10), 720 => to_unsigned(201, 10), 721 => to_unsigned(944, 10), 722 => to_unsigned(725, 10), 723 => to_unsigned(760, 10), 724 => to_unsigned(859, 10), 725 => to_unsigned(567, 10), 726 => to_unsigned(886, 10), 727 => to_unsigned(336, 10), 728 => to_unsigned(230, 10), 729 => to_unsigned(347, 10), 730 => to_unsigned(377, 10), 731 => to_unsigned(381, 10), 732 => to_unsigned(934, 10), 733 => to_unsigned(974, 10), 734 => to_unsigned(427, 10), 735 => to_unsigned(556, 10), 736 => to_unsigned(586, 10), 737 => to_unsigned(1010, 10), 738 => to_unsigned(885, 10), 739 => to_unsigned(29, 10), 740 => to_unsigned(741, 10), 741 => to_unsigned(27, 10), 742 => to_unsigned(284, 10), 743 => to_unsigned(982, 10), 744 => to_unsigned(999, 10), 745 => to_unsigned(852, 10), 746 => to_unsigned(608, 10), 747 => to_unsigned(117, 10), 748 => to_unsigned(716, 10), 749 => to_unsigned(953, 10), 750 => to_unsigned(1012, 10), 751 => to_unsigned(413, 10), 752 => to_unsigned(122, 10), 753 => to_unsigned(561, 10), 754 => to_unsigned(579, 10), 755 => to_unsigned(431, 10), 756 => to_unsigned(843, 10), 757 => to_unsigned(278, 10), 758 => to_unsigned(329, 10), 759 => to_unsigned(311, 10), 760 => to_unsigned(476, 10), 761 => to_unsigned(1004, 10), 762 => to_unsigned(529, 10), 763 => to_unsigned(662, 10), 764 => to_unsigned(198, 10), 765 => to_unsigned(79, 10), 766 => to_unsigned(871, 10), 767 => to_unsigned(531, 10), 768 => to_unsigned(90, 10), 769 => to_unsigned(343, 10), 770 => to_unsigned(875, 10), 771 => to_unsigned(827, 10), 772 => to_unsigned(463, 10), 773 => to_unsigned(882, 10), 774 => to_unsigned(340, 10), 775 => to_unsigned(945, 10), 776 => to_unsigned(693, 10), 777 => to_unsigned(429, 10), 778 => to_unsigned(172, 10), 779 => to_unsigned(222, 10), 780 => to_unsigned(683, 10), 781 => to_unsigned(865, 10), 782 => to_unsigned(512, 10), 783 => to_unsigned(719, 10), 784 => to_unsigned(362, 10), 785 => to_unsigned(223, 10), 786 => to_unsigned(348, 10), 787 => to_unsigned(391, 10), 788 => to_unsigned(221, 10), 789 => to_unsigned(781, 10), 790 => to_unsigned(346, 10), 791 => to_unsigned(742, 10), 792 => to_unsigned(580, 10), 793 => to_unsigned(621, 10), 794 => to_unsigned(739, 10), 795 => to_unsigned(609, 10), 796 => to_unsigned(942, 10), 797 => to_unsigned(521, 10), 798 => to_unsigned(838, 10), 799 => to_unsigned(677, 10), 800 => to_unsigned(547, 10), 801 => to_unsigned(782, 10), 802 => to_unsigned(146, 10), 803 => to_unsigned(820, 10), 804 => to_unsigned(927, 10), 805 => to_unsigned(397, 10), 806 => to_unsigned(884, 10), 807 => to_unsigned(197, 10), 808 => to_unsigned(851, 10), 809 => to_unsigned(941, 10), 810 => to_unsigned(172, 10), 811 => to_unsigned(589, 10), 812 => to_unsigned(830, 10), 813 => to_unsigned(756, 10), 814 => to_unsigned(241, 10), 815 => to_unsigned(693, 10), 816 => to_unsigned(411, 10), 817 => to_unsigned(280, 10), 818 => to_unsigned(673, 10), 819 => to_unsigned(644, 10), 820 => to_unsigned(950, 10), 821 => to_unsigned(249, 10), 822 => to_unsigned(300, 10), 823 => to_unsigned(76, 10), 824 => to_unsigned(795, 10), 825 => to_unsigned(333, 10), 826 => to_unsigned(590, 10), 827 => to_unsigned(65, 10), 828 => to_unsigned(966, 10), 829 => to_unsigned(535, 10), 830 => to_unsigned(262, 10), 831 => to_unsigned(228, 10), 832 => to_unsigned(698, 10), 833 => to_unsigned(707, 10), 834 => to_unsigned(259, 10), 835 => to_unsigned(307, 10), 836 => to_unsigned(643, 10), 837 => to_unsigned(828, 10), 838 => to_unsigned(870, 10), 839 => to_unsigned(748, 10), 840 => to_unsigned(324, 10), 841 => to_unsigned(827, 10), 842 => to_unsigned(286, 10), 843 => to_unsigned(778, 10), 844 => to_unsigned(326, 10), 845 => to_unsigned(486, 10), 846 => to_unsigned(159, 10), 847 => to_unsigned(175, 10), 848 => to_unsigned(120, 10), 849 => to_unsigned(736, 10), 850 => to_unsigned(936, 10), 851 => to_unsigned(63, 10), 852 => to_unsigned(920, 10), 853 => to_unsigned(437, 10), 854 => to_unsigned(25, 10), 855 => to_unsigned(858, 10), 856 => to_unsigned(477, 10), 857 => to_unsigned(758, 10), 858 => to_unsigned(837, 10), 859 => to_unsigned(460, 10), 860 => to_unsigned(3, 10), 861 => to_unsigned(83, 10), 862 => to_unsigned(228, 10), 863 => to_unsigned(1, 10), 864 => to_unsigned(645, 10), 865 => to_unsigned(43, 10), 866 => to_unsigned(107, 10), 867 => to_unsigned(783, 10), 868 => to_unsigned(140, 10), 869 => to_unsigned(311, 10), 870 => to_unsigned(251, 10), 871 => to_unsigned(633, 10), 872 => to_unsigned(437, 10), 873 => to_unsigned(427, 10), 874 => to_unsigned(136, 10), 875 => to_unsigned(486, 10), 876 => to_unsigned(181, 10), 877 => to_unsigned(607, 10), 878 => to_unsigned(966, 10), 879 => to_unsigned(681, 10), 880 => to_unsigned(632, 10), 881 => to_unsigned(7, 10), 882 => to_unsigned(48, 10), 883 => to_unsigned(437, 10), 884 => to_unsigned(871, 10), 885 => to_unsigned(205, 10), 886 => to_unsigned(264, 10), 887 => to_unsigned(173, 10), 888 => to_unsigned(853, 10), 889 => to_unsigned(518, 10), 890 => to_unsigned(507, 10), 891 => to_unsigned(907, 10), 892 => to_unsigned(713, 10), 893 => to_unsigned(161, 10), 894 => to_unsigned(652, 10), 895 => to_unsigned(499, 10), 896 => to_unsigned(751, 10), 897 => to_unsigned(498, 10), 898 => to_unsigned(895, 10), 899 => to_unsigned(932, 10), 900 => to_unsigned(258, 10), 901 => to_unsigned(475, 10), 902 => to_unsigned(283, 10), 903 => to_unsigned(375, 10), 904 => to_unsigned(100, 10), 905 => to_unsigned(888, 10), 906 => to_unsigned(442, 10), 907 => to_unsigned(783, 10), 908 => to_unsigned(41, 10), 909 => to_unsigned(806, 10), 910 => to_unsigned(296, 10), 911 => to_unsigned(661, 10), 912 => to_unsigned(242, 10), 913 => to_unsigned(241, 10), 914 => to_unsigned(479, 10), 915 => to_unsigned(136, 10), 916 => to_unsigned(684, 10), 917 => to_unsigned(994, 10), 918 => to_unsigned(200, 10), 919 => to_unsigned(834, 10), 920 => to_unsigned(144, 10), 921 => to_unsigned(168, 10), 922 => to_unsigned(395, 10), 923 => to_unsigned(970, 10), 924 => to_unsigned(396, 10), 925 => to_unsigned(18, 10), 926 => to_unsigned(629, 10), 927 => to_unsigned(115, 10), 928 => to_unsigned(537, 10), 929 => to_unsigned(68, 10), 930 => to_unsigned(948, 10), 931 => to_unsigned(897, 10), 932 => to_unsigned(133, 10), 933 => to_unsigned(834, 10), 934 => to_unsigned(770, 10), 935 => to_unsigned(44, 10), 936 => to_unsigned(373, 10), 937 => to_unsigned(491, 10), 938 => to_unsigned(39, 10), 939 => to_unsigned(49, 10), 940 => to_unsigned(914, 10), 941 => to_unsigned(336, 10), 942 => to_unsigned(17, 10), 943 => to_unsigned(879, 10), 944 => to_unsigned(437, 10), 945 => to_unsigned(852, 10), 946 => to_unsigned(1004, 10), 947 => to_unsigned(206, 10), 948 => to_unsigned(852, 10), 949 => to_unsigned(289, 10), 950 => to_unsigned(969, 10), 951 => to_unsigned(648, 10), 952 => to_unsigned(241, 10), 953 => to_unsigned(728, 10), 954 => to_unsigned(153, 10), 955 => to_unsigned(418, 10), 956 => to_unsigned(479, 10), 957 => to_unsigned(611, 10), 958 => to_unsigned(18, 10), 959 => to_unsigned(251, 10), 960 => to_unsigned(1022, 10), 961 => to_unsigned(645, 10), 962 => to_unsigned(684, 10), 963 => to_unsigned(407, 10), 964 => to_unsigned(696, 10), 965 => to_unsigned(417, 10), 966 => to_unsigned(496, 10), 967 => to_unsigned(862, 10), 968 => to_unsigned(162, 10), 969 => to_unsigned(541, 10), 970 => to_unsigned(894, 10), 971 => to_unsigned(780, 10), 972 => to_unsigned(298, 10), 973 => to_unsigned(583, 10), 974 => to_unsigned(499, 10), 975 => to_unsigned(836, 10), 976 => to_unsigned(235, 10), 977 => to_unsigned(939, 10), 978 => to_unsigned(576, 10), 979 => to_unsigned(64, 10), 980 => to_unsigned(806, 10), 981 => to_unsigned(177, 10), 982 => to_unsigned(713, 10), 983 => to_unsigned(212, 10), 984 => to_unsigned(584, 10), 985 => to_unsigned(560, 10), 986 => to_unsigned(582, 10), 987 => to_unsigned(884, 10), 988 => to_unsigned(823, 10), 989 => to_unsigned(788, 10), 990 => to_unsigned(364, 10), 991 => to_unsigned(953, 10), 992 => to_unsigned(1, 10), 993 => to_unsigned(361, 10), 994 => to_unsigned(772, 10), 995 => to_unsigned(348, 10), 996 => to_unsigned(65, 10), 997 => to_unsigned(339, 10), 998 => to_unsigned(174, 10), 999 => to_unsigned(734, 10), 1000 => to_unsigned(322, 10), 1001 => to_unsigned(400, 10), 1002 => to_unsigned(559, 10), 1003 => to_unsigned(718, 10), 1004 => to_unsigned(470, 10), 1005 => to_unsigned(248, 10), 1006 => to_unsigned(272, 10), 1007 => to_unsigned(587, 10), 1008 => to_unsigned(974, 10), 1009 => to_unsigned(404, 10), 1010 => to_unsigned(927, 10), 1011 => to_unsigned(202, 10), 1012 => to_unsigned(360, 10), 1013 => to_unsigned(633, 10), 1014 => to_unsigned(142, 10), 1015 => to_unsigned(166, 10), 1016 => to_unsigned(651, 10), 1017 => to_unsigned(13, 10), 1018 => to_unsigned(558, 10), 1019 => to_unsigned(507, 10), 1020 => to_unsigned(256, 10), 1021 => to_unsigned(936, 10), 1022 => to_unsigned(7, 10), 1023 => to_unsigned(396, 10), 1024 => to_unsigned(124, 10), 1025 => to_unsigned(769, 10), 1026 => to_unsigned(146, 10), 1027 => to_unsigned(44, 10), 1028 => to_unsigned(323, 10), 1029 => to_unsigned(430, 10), 1030 => to_unsigned(322, 10), 1031 => to_unsigned(918, 10), 1032 => to_unsigned(636, 10), 1033 => to_unsigned(501, 10), 1034 => to_unsigned(922, 10), 1035 => to_unsigned(445, 10), 1036 => to_unsigned(274, 10), 1037 => to_unsigned(162, 10), 1038 => to_unsigned(457, 10), 1039 => to_unsigned(1018, 10), 1040 => to_unsigned(563, 10), 1041 => to_unsigned(491, 10), 1042 => to_unsigned(323, 10), 1043 => to_unsigned(972, 10), 1044 => to_unsigned(809, 10), 1045 => to_unsigned(806, 10), 1046 => to_unsigned(880, 10), 1047 => to_unsigned(1007, 10), 1048 => to_unsigned(285, 10), 1049 => to_unsigned(981, 10), 1050 => to_unsigned(577, 10), 1051 => to_unsigned(474, 10), 1052 => to_unsigned(52, 10), 1053 => to_unsigned(31, 10), 1054 => to_unsigned(155, 10), 1055 => to_unsigned(895, 10), 1056 => to_unsigned(520, 10), 1057 => to_unsigned(657, 10), 1058 => to_unsigned(280, 10), 1059 => to_unsigned(518, 10), 1060 => to_unsigned(622, 10), 1061 => to_unsigned(6, 10), 1062 => to_unsigned(90, 10), 1063 => to_unsigned(139, 10), 1064 => to_unsigned(444, 10), 1065 => to_unsigned(599, 10), 1066 => to_unsigned(495, 10), 1067 => to_unsigned(204, 10), 1068 => to_unsigned(95, 10), 1069 => to_unsigned(735, 10), 1070 => to_unsigned(336, 10), 1071 => to_unsigned(999, 10), 1072 => to_unsigned(29, 10), 1073 => to_unsigned(1007, 10), 1074 => to_unsigned(727, 10), 1075 => to_unsigned(109, 10), 1076 => to_unsigned(292, 10), 1077 => to_unsigned(240, 10), 1078 => to_unsigned(857, 10), 1079 => to_unsigned(473, 10), 1080 => to_unsigned(357, 10), 1081 => to_unsigned(401, 10), 1082 => to_unsigned(914, 10), 1083 => to_unsigned(685, 10), 1084 => to_unsigned(118, 10), 1085 => to_unsigned(406, 10), 1086 => to_unsigned(315, 10), 1087 => to_unsigned(2, 10), 1088 => to_unsigned(869, 10), 1089 => to_unsigned(174, 10), 1090 => to_unsigned(730, 10), 1091 => to_unsigned(521, 10), 1092 => to_unsigned(680, 10), 1093 => to_unsigned(434, 10), 1094 => to_unsigned(449, 10), 1095 => to_unsigned(155, 10), 1096 => to_unsigned(483, 10), 1097 => to_unsigned(428, 10), 1098 => to_unsigned(234, 10), 1099 => to_unsigned(941, 10), 1100 => to_unsigned(332, 10), 1101 => to_unsigned(774, 10), 1102 => to_unsigned(111, 10), 1103 => to_unsigned(208, 10), 1104 => to_unsigned(83, 10), 1105 => to_unsigned(52, 10), 1106 => to_unsigned(552, 10), 1107 => to_unsigned(175, 10), 1108 => to_unsigned(881, 10), 1109 => to_unsigned(671, 10), 1110 => to_unsigned(191, 10), 1111 => to_unsigned(450, 10), 1112 => to_unsigned(1016, 10), 1113 => to_unsigned(590, 10), 1114 => to_unsigned(780, 10), 1115 => to_unsigned(584, 10), 1116 => to_unsigned(280, 10), 1117 => to_unsigned(115, 10), 1118 => to_unsigned(13, 10), 1119 => to_unsigned(137, 10), 1120 => to_unsigned(614, 10), 1121 => to_unsigned(466, 10), 1122 => to_unsigned(585, 10), 1123 => to_unsigned(937, 10), 1124 => to_unsigned(366, 10), 1125 => to_unsigned(355, 10), 1126 => to_unsigned(834, 10), 1127 => to_unsigned(313, 10), 1128 => to_unsigned(552, 10), 1129 => to_unsigned(599, 10), 1130 => to_unsigned(694, 10), 1131 => to_unsigned(356, 10), 1132 => to_unsigned(716, 10), 1133 => to_unsigned(98, 10), 1134 => to_unsigned(476, 10), 1135 => to_unsigned(368, 10), 1136 => to_unsigned(269, 10), 1137 => to_unsigned(292, 10), 1138 => to_unsigned(1003, 10), 1139 => to_unsigned(586, 10), 1140 => to_unsigned(847, 10), 1141 => to_unsigned(298, 10), 1142 => to_unsigned(484, 10), 1143 => to_unsigned(422, 10), 1144 => to_unsigned(862, 10), 1145 => to_unsigned(427, 10), 1146 => to_unsigned(789, 10), 1147 => to_unsigned(835, 10), 1148 => to_unsigned(716, 10), 1149 => to_unsigned(530, 10), 1150 => to_unsigned(145, 10), 1151 => to_unsigned(606, 10), 1152 => to_unsigned(698, 10), 1153 => to_unsigned(678, 10), 1154 => to_unsigned(340, 10), 1155 => to_unsigned(721, 10), 1156 => to_unsigned(45, 10), 1157 => to_unsigned(945, 10), 1158 => to_unsigned(288, 10), 1159 => to_unsigned(370, 10), 1160 => to_unsigned(829, 10), 1161 => to_unsigned(260, 10), 1162 => to_unsigned(291, 10), 1163 => to_unsigned(726, 10), 1164 => to_unsigned(179, 10), 1165 => to_unsigned(643, 10), 1166 => to_unsigned(935, 10), 1167 => to_unsigned(180, 10), 1168 => to_unsigned(667, 10), 1169 => to_unsigned(661, 10), 1170 => to_unsigned(743, 10), 1171 => to_unsigned(58, 10), 1172 => to_unsigned(533, 10), 1173 => to_unsigned(530, 10), 1174 => to_unsigned(791, 10), 1175 => to_unsigned(498, 10), 1176 => to_unsigned(719, 10), 1177 => to_unsigned(383, 10), 1178 => to_unsigned(665, 10), 1179 => to_unsigned(310, 10), 1180 => to_unsigned(718, 10), 1181 => to_unsigned(32, 10), 1182 => to_unsigned(280, 10), 1183 => to_unsigned(508, 10), 1184 => to_unsigned(4, 10), 1185 => to_unsigned(126, 10), 1186 => to_unsigned(848, 10), 1187 => to_unsigned(361, 10), 1188 => to_unsigned(227, 10), 1189 => to_unsigned(978, 10), 1190 => to_unsigned(772, 10), 1191 => to_unsigned(503, 10), 1192 => to_unsigned(727, 10), 1193 => to_unsigned(502, 10), 1194 => to_unsigned(1010, 10), 1195 => to_unsigned(89, 10), 1196 => to_unsigned(40, 10), 1197 => to_unsigned(732, 10), 1198 => to_unsigned(333, 10), 1199 => to_unsigned(911, 10), 1200 => to_unsigned(50, 10), 1201 => to_unsigned(712, 10), 1202 => to_unsigned(947, 10), 1203 => to_unsigned(955, 10), 1204 => to_unsigned(92, 10), 1205 => to_unsigned(579, 10), 1206 => to_unsigned(512, 10), 1207 => to_unsigned(785, 10), 1208 => to_unsigned(749, 10), 1209 => to_unsigned(879, 10), 1210 => to_unsigned(845, 10), 1211 => to_unsigned(649, 10), 1212 => to_unsigned(652, 10), 1213 => to_unsigned(392, 10), 1214 => to_unsigned(506, 10), 1215 => to_unsigned(574, 10), 1216 => to_unsigned(467, 10), 1217 => to_unsigned(580, 10), 1218 => to_unsigned(237, 10), 1219 => to_unsigned(267, 10), 1220 => to_unsigned(541, 10), 1221 => to_unsigned(799, 10), 1222 => to_unsigned(25, 10), 1223 => to_unsigned(616, 10), 1224 => to_unsigned(416, 10), 1225 => to_unsigned(618, 10), 1226 => to_unsigned(349, 10), 1227 => to_unsigned(760, 10), 1228 => to_unsigned(389, 10), 1229 => to_unsigned(256, 10), 1230 => to_unsigned(653, 10), 1231 => to_unsigned(759, 10), 1232 => to_unsigned(842, 10), 1233 => to_unsigned(475, 10), 1234 => to_unsigned(28, 10), 1235 => to_unsigned(452, 10), 1236 => to_unsigned(175, 10), 1237 => to_unsigned(434, 10), 1238 => to_unsigned(117, 10), 1239 => to_unsigned(421, 10), 1240 => to_unsigned(543, 10), 1241 => to_unsigned(480, 10), 1242 => to_unsigned(273, 10), 1243 => to_unsigned(760, 10), 1244 => to_unsigned(553, 10), 1245 => to_unsigned(946, 10), 1246 => to_unsigned(632, 10), 1247 => to_unsigned(627, 10), 1248 => to_unsigned(304, 10), 1249 => to_unsigned(384, 10), 1250 => to_unsigned(710, 10), 1251 => to_unsigned(383, 10), 1252 => to_unsigned(617, 10), 1253 => to_unsigned(858, 10), 1254 => to_unsigned(460, 10), 1255 => to_unsigned(634, 10), 1256 => to_unsigned(43, 10), 1257 => to_unsigned(537, 10), 1258 => to_unsigned(854, 10), 1259 => to_unsigned(684, 10), 1260 => to_unsigned(866, 10), 1261 => to_unsigned(801, 10), 1262 => to_unsigned(417, 10), 1263 => to_unsigned(76, 10), 1264 => to_unsigned(86, 10), 1265 => to_unsigned(802, 10), 1266 => to_unsigned(892, 10), 1267 => to_unsigned(85, 10), 1268 => to_unsigned(266, 10), 1269 => to_unsigned(578, 10), 1270 => to_unsigned(188, 10), 1271 => to_unsigned(586, 10), 1272 => to_unsigned(801, 10), 1273 => to_unsigned(798, 10), 1274 => to_unsigned(496, 10), 1275 => to_unsigned(327, 10), 1276 => to_unsigned(879, 10), 1277 => to_unsigned(668, 10), 1278 => to_unsigned(223, 10), 1279 => to_unsigned(124, 10), 1280 => to_unsigned(266, 10), 1281 => to_unsigned(646, 10), 1282 => to_unsigned(824, 10), 1283 => to_unsigned(227, 10), 1284 => to_unsigned(599, 10), 1285 => to_unsigned(131, 10), 1286 => to_unsigned(881, 10), 1287 => to_unsigned(780, 10), 1288 => to_unsigned(348, 10), 1289 => to_unsigned(131, 10), 1290 => to_unsigned(552, 10), 1291 => to_unsigned(380, 10), 1292 => to_unsigned(983, 10), 1293 => to_unsigned(643, 10), 1294 => to_unsigned(854, 10), 1295 => to_unsigned(928, 10), 1296 => to_unsigned(663, 10), 1297 => to_unsigned(34, 10), 1298 => to_unsigned(237, 10), 1299 => to_unsigned(253, 10), 1300 => to_unsigned(889, 10), 1301 => to_unsigned(916, 10), 1302 => to_unsigned(704, 10), 1303 => to_unsigned(883, 10), 1304 => to_unsigned(231, 10), 1305 => to_unsigned(287, 10), 1306 => to_unsigned(359, 10), 1307 => to_unsigned(784, 10), 1308 => to_unsigned(572, 10), 1309 => to_unsigned(214, 10), 1310 => to_unsigned(220, 10), 1311 => to_unsigned(619, 10), 1312 => to_unsigned(814, 10), 1313 => to_unsigned(754, 10), 1314 => to_unsigned(126, 10), 1315 => to_unsigned(987, 10), 1316 => to_unsigned(73, 10), 1317 => to_unsigned(684, 10), 1318 => to_unsigned(223, 10), 1319 => to_unsigned(53, 10), 1320 => to_unsigned(271, 10), 1321 => to_unsigned(805, 10), 1322 => to_unsigned(502, 10), 1323 => to_unsigned(833, 10), 1324 => to_unsigned(228, 10), 1325 => to_unsigned(399, 10), 1326 => to_unsigned(628, 10), 1327 => to_unsigned(510, 10), 1328 => to_unsigned(407, 10), 1329 => to_unsigned(965, 10), 1330 => to_unsigned(787, 10), 1331 => to_unsigned(479, 10), 1332 => to_unsigned(641, 10), 1333 => to_unsigned(699, 10), 1334 => to_unsigned(20, 10), 1335 => to_unsigned(971, 10), 1336 => to_unsigned(1005, 10), 1337 => to_unsigned(390, 10), 1338 => to_unsigned(311, 10), 1339 => to_unsigned(904, 10), 1340 => to_unsigned(514, 10), 1341 => to_unsigned(954, 10), 1342 => to_unsigned(162, 10), 1343 => to_unsigned(622, 10), 1344 => to_unsigned(367, 10), 1345 => to_unsigned(143, 10), 1346 => to_unsigned(842, 10), 1347 => to_unsigned(432, 10), 1348 => to_unsigned(366, 10), 1349 => to_unsigned(362, 10), 1350 => to_unsigned(888, 10), 1351 => to_unsigned(591, 10), 1352 => to_unsigned(937, 10), 1353 => to_unsigned(884, 10), 1354 => to_unsigned(826, 10), 1355 => to_unsigned(422, 10), 1356 => to_unsigned(850, 10), 1357 => to_unsigned(966, 10), 1358 => to_unsigned(289, 10), 1359 => to_unsigned(607, 10), 1360 => to_unsigned(184, 10), 1361 => to_unsigned(331, 10), 1362 => to_unsigned(881, 10), 1363 => to_unsigned(27, 10), 1364 => to_unsigned(279, 10), 1365 => to_unsigned(458, 10), 1366 => to_unsigned(555, 10), 1367 => to_unsigned(1010, 10), 1368 => to_unsigned(372, 10), 1369 => to_unsigned(116, 10), 1370 => to_unsigned(822, 10), 1371 => to_unsigned(808, 10), 1372 => to_unsigned(181, 10), 1373 => to_unsigned(453, 10), 1374 => to_unsigned(46, 10), 1375 => to_unsigned(380, 10), 1376 => to_unsigned(130, 10), 1377 => to_unsigned(800, 10), 1378 => to_unsigned(621, 10), 1379 => to_unsigned(848, 10), 1380 => to_unsigned(729, 10), 1381 => to_unsigned(699, 10), 1382 => to_unsigned(574, 10), 1383 => to_unsigned(908, 10), 1384 => to_unsigned(338, 10), 1385 => to_unsigned(22, 10), 1386 => to_unsigned(431, 10), 1387 => to_unsigned(650, 10), 1388 => to_unsigned(560, 10), 1389 => to_unsigned(286, 10), 1390 => to_unsigned(67, 10), 1391 => to_unsigned(136, 10), 1392 => to_unsigned(175, 10), 1393 => to_unsigned(925, 10), 1394 => to_unsigned(1020, 10), 1395 => to_unsigned(434, 10), 1396 => to_unsigned(973, 10), 1397 => to_unsigned(921, 10), 1398 => to_unsigned(282, 10), 1399 => to_unsigned(45, 10), 1400 => to_unsigned(856, 10), 1401 => to_unsigned(844, 10), 1402 => to_unsigned(203, 10), 1403 => to_unsigned(568, 10), 1404 => to_unsigned(291, 10), 1405 => to_unsigned(422, 10), 1406 => to_unsigned(66, 10), 1407 => to_unsigned(936, 10), 1408 => to_unsigned(329, 10), 1409 => to_unsigned(812, 10), 1410 => to_unsigned(456, 10), 1411 => to_unsigned(650, 10), 1412 => to_unsigned(529, 10), 1413 => to_unsigned(425, 10), 1414 => to_unsigned(145, 10), 1415 => to_unsigned(528, 10), 1416 => to_unsigned(160, 10), 1417 => to_unsigned(101, 10), 1418 => to_unsigned(133, 10), 1419 => to_unsigned(73, 10), 1420 => to_unsigned(645, 10), 1421 => to_unsigned(271, 10), 1422 => to_unsigned(277, 10), 1423 => to_unsigned(930, 10), 1424 => to_unsigned(678, 10), 1425 => to_unsigned(638, 10), 1426 => to_unsigned(928, 10), 1427 => to_unsigned(790, 10), 1428 => to_unsigned(137, 10), 1429 => to_unsigned(783, 10), 1430 => to_unsigned(400, 10), 1431 => to_unsigned(410, 10), 1432 => to_unsigned(875, 10), 1433 => to_unsigned(659, 10), 1434 => to_unsigned(512, 10), 1435 => to_unsigned(877, 10), 1436 => to_unsigned(157, 10), 1437 => to_unsigned(1023, 10), 1438 => to_unsigned(770, 10), 1439 => to_unsigned(700, 10), 1440 => to_unsigned(594, 10), 1441 => to_unsigned(169, 10), 1442 => to_unsigned(789, 10), 1443 => to_unsigned(615, 10), 1444 => to_unsigned(434, 10), 1445 => to_unsigned(661, 10), 1446 => to_unsigned(197, 10), 1447 => to_unsigned(626, 10), 1448 => to_unsigned(320, 10), 1449 => to_unsigned(583, 10), 1450 => to_unsigned(225, 10), 1451 => to_unsigned(841, 10), 1452 => to_unsigned(851, 10), 1453 => to_unsigned(178, 10), 1454 => to_unsigned(380, 10), 1455 => to_unsigned(903, 10), 1456 => to_unsigned(952, 10), 1457 => to_unsigned(1007, 10), 1458 => to_unsigned(662, 10), 1459 => to_unsigned(328, 10), 1460 => to_unsigned(64, 10), 1461 => to_unsigned(730, 10), 1462 => to_unsigned(917, 10), 1463 => to_unsigned(48, 10), 1464 => to_unsigned(738, 10), 1465 => to_unsigned(588, 10), 1466 => to_unsigned(969, 10), 1467 => to_unsigned(147, 10), 1468 => to_unsigned(407, 10), 1469 => to_unsigned(562, 10), 1470 => to_unsigned(884, 10), 1471 => to_unsigned(353, 10), 1472 => to_unsigned(620, 10), 1473 => to_unsigned(862, 10), 1474 => to_unsigned(140, 10), 1475 => to_unsigned(291, 10), 1476 => to_unsigned(463, 10), 1477 => to_unsigned(303, 10), 1478 => to_unsigned(416, 10), 1479 => to_unsigned(739, 10), 1480 => to_unsigned(467, 10), 1481 => to_unsigned(878, 10), 1482 => to_unsigned(669, 10), 1483 => to_unsigned(745, 10), 1484 => to_unsigned(157, 10), 1485 => to_unsigned(36, 10), 1486 => to_unsigned(298, 10), 1487 => to_unsigned(952, 10), 1488 => to_unsigned(436, 10), 1489 => to_unsigned(541, 10), 1490 => to_unsigned(946, 10), 1491 => to_unsigned(582, 10), 1492 => to_unsigned(340, 10), 1493 => to_unsigned(338, 10), 1494 => to_unsigned(323, 10), 1495 => to_unsigned(725, 10), 1496 => to_unsigned(73, 10), 1497 => to_unsigned(1018, 10), 1498 => to_unsigned(75, 10), 1499 => to_unsigned(187, 10), 1500 => to_unsigned(362, 10), 1501 => to_unsigned(221, 10), 1502 => to_unsigned(268, 10), 1503 => to_unsigned(119, 10), 1504 => to_unsigned(1001, 10), 1505 => to_unsigned(720, 10), 1506 => to_unsigned(225, 10), 1507 => to_unsigned(55, 10), 1508 => to_unsigned(767, 10), 1509 => to_unsigned(41, 10), 1510 => to_unsigned(306, 10), 1511 => to_unsigned(375, 10), 1512 => to_unsigned(501, 10), 1513 => to_unsigned(154, 10), 1514 => to_unsigned(346, 10), 1515 => to_unsigned(393, 10), 1516 => to_unsigned(387, 10), 1517 => to_unsigned(912, 10), 1518 => to_unsigned(449, 10), 1519 => to_unsigned(621, 10), 1520 => to_unsigned(681, 10), 1521 => to_unsigned(160, 10), 1522 => to_unsigned(953, 10), 1523 => to_unsigned(200, 10), 1524 => to_unsigned(940, 10), 1525 => to_unsigned(627, 10), 1526 => to_unsigned(598, 10), 1527 => to_unsigned(765, 10), 1528 => to_unsigned(696, 10), 1529 => to_unsigned(363, 10), 1530 => to_unsigned(987, 10), 1531 => to_unsigned(261, 10), 1532 => to_unsigned(669, 10), 1533 => to_unsigned(502, 10), 1534 => to_unsigned(106, 10), 1535 => to_unsigned(856, 10), 1536 => to_unsigned(657, 10), 1537 => to_unsigned(803, 10), 1538 => to_unsigned(811, 10), 1539 => to_unsigned(435, 10), 1540 => to_unsigned(843, 10), 1541 => to_unsigned(989, 10), 1542 => to_unsigned(703, 10), 1543 => to_unsigned(696, 10), 1544 => to_unsigned(231, 10), 1545 => to_unsigned(403, 10), 1546 => to_unsigned(350, 10), 1547 => to_unsigned(660, 10), 1548 => to_unsigned(167, 10), 1549 => to_unsigned(912, 10), 1550 => to_unsigned(970, 10), 1551 => to_unsigned(495, 10), 1552 => to_unsigned(548, 10), 1553 => to_unsigned(485, 10), 1554 => to_unsigned(85, 10), 1555 => to_unsigned(894, 10), 1556 => to_unsigned(682, 10), 1557 => to_unsigned(64, 10), 1558 => to_unsigned(338, 10), 1559 => to_unsigned(275, 10), 1560 => to_unsigned(698, 10), 1561 => to_unsigned(524, 10), 1562 => to_unsigned(349, 10), 1563 => to_unsigned(384, 10), 1564 => to_unsigned(454, 10), 1565 => to_unsigned(490, 10), 1566 => to_unsigned(874, 10), 1567 => to_unsigned(275, 10), 1568 => to_unsigned(905, 10), 1569 => to_unsigned(400, 10), 1570 => to_unsigned(142, 10), 1571 => to_unsigned(61, 10), 1572 => to_unsigned(626, 10), 1573 => to_unsigned(705, 10), 1574 => to_unsigned(285, 10), 1575 => to_unsigned(817, 10), 1576 => to_unsigned(147, 10), 1577 => to_unsigned(21, 10), 1578 => to_unsigned(570, 10), 1579 => to_unsigned(767, 10), 1580 => to_unsigned(920, 10), 1581 => to_unsigned(620, 10), 1582 => to_unsigned(84, 10), 1583 => to_unsigned(221, 10), 1584 => to_unsigned(627, 10), 1585 => to_unsigned(550, 10), 1586 => to_unsigned(581, 10), 1587 => to_unsigned(593, 10), 1588 => to_unsigned(648, 10), 1589 => to_unsigned(174, 10), 1590 => to_unsigned(755, 10), 1591 => to_unsigned(351, 10), 1592 => to_unsigned(875, 10), 1593 => to_unsigned(606, 10), 1594 => to_unsigned(994, 10), 1595 => to_unsigned(1020, 10), 1596 => to_unsigned(597, 10), 1597 => to_unsigned(165, 10), 1598 => to_unsigned(303, 10), 1599 => to_unsigned(630, 10), 1600 => to_unsigned(472, 10), 1601 => to_unsigned(822, 10), 1602 => to_unsigned(482, 10), 1603 => to_unsigned(818, 10), 1604 => to_unsigned(1018, 10), 1605 => to_unsigned(515, 10), 1606 => to_unsigned(651, 10), 1607 => to_unsigned(383, 10), 1608 => to_unsigned(671, 10), 1609 => to_unsigned(879, 10), 1610 => to_unsigned(658, 10), 1611 => to_unsigned(538, 10), 1612 => to_unsigned(420, 10), 1613 => to_unsigned(1000, 10), 1614 => to_unsigned(122, 10), 1615 => to_unsigned(617, 10), 1616 => to_unsigned(696, 10), 1617 => to_unsigned(574, 10), 1618 => to_unsigned(277, 10), 1619 => to_unsigned(94, 10), 1620 => to_unsigned(833, 10), 1621 => to_unsigned(237, 10), 1622 => to_unsigned(437, 10), 1623 => to_unsigned(923, 10), 1624 => to_unsigned(300, 10), 1625 => to_unsigned(525, 10), 1626 => to_unsigned(914, 10), 1627 => to_unsigned(885, 10), 1628 => to_unsigned(835, 10), 1629 => to_unsigned(22, 10), 1630 => to_unsigned(1008, 10), 1631 => to_unsigned(379, 10), 1632 => to_unsigned(740, 10), 1633 => to_unsigned(111, 10), 1634 => to_unsigned(225, 10), 1635 => to_unsigned(787, 10), 1636 => to_unsigned(119, 10), 1637 => to_unsigned(478, 10), 1638 => to_unsigned(310, 10), 1639 => to_unsigned(656, 10), 1640 => to_unsigned(655, 10), 1641 => to_unsigned(943, 10), 1642 => to_unsigned(158, 10), 1643 => to_unsigned(256, 10), 1644 => to_unsigned(938, 10), 1645 => to_unsigned(635, 10), 1646 => to_unsigned(16, 10), 1647 => to_unsigned(727, 10), 1648 => to_unsigned(464, 10), 1649 => to_unsigned(204, 10), 1650 => to_unsigned(828, 10), 1651 => to_unsigned(617, 10), 1652 => to_unsigned(895, 10), 1653 => to_unsigned(686, 10), 1654 => to_unsigned(448, 10), 1655 => to_unsigned(629, 10), 1656 => to_unsigned(503, 10), 1657 => to_unsigned(618, 10), 1658 => to_unsigned(878, 10), 1659 => to_unsigned(256, 10), 1660 => to_unsigned(833, 10), 1661 => to_unsigned(667, 10), 1662 => to_unsigned(546, 10), 1663 => to_unsigned(534, 10), 1664 => to_unsigned(946, 10), 1665 => to_unsigned(864, 10), 1666 => to_unsigned(1004, 10), 1667 => to_unsigned(907, 10), 1668 => to_unsigned(711, 10), 1669 => to_unsigned(109, 10), 1670 => to_unsigned(348, 10), 1671 => to_unsigned(627, 10), 1672 => to_unsigned(160, 10), 1673 => to_unsigned(97, 10), 1674 => to_unsigned(921, 10), 1675 => to_unsigned(374, 10), 1676 => to_unsigned(538, 10), 1677 => to_unsigned(133, 10), 1678 => to_unsigned(657, 10), 1679 => to_unsigned(98, 10), 1680 => to_unsigned(184, 10), 1681 => to_unsigned(422, 10), 1682 => to_unsigned(260, 10), 1683 => to_unsigned(431, 10), 1684 => to_unsigned(1020, 10), 1685 => to_unsigned(50, 10), 1686 => to_unsigned(882, 10), 1687 => to_unsigned(428, 10), 1688 => to_unsigned(109, 10), 1689 => to_unsigned(726, 10), 1690 => to_unsigned(27, 10), 1691 => to_unsigned(954, 10), 1692 => to_unsigned(320, 10), 1693 => to_unsigned(436, 10), 1694 => to_unsigned(386, 10), 1695 => to_unsigned(578, 10), 1696 => to_unsigned(502, 10), 1697 => to_unsigned(148, 10), 1698 => to_unsigned(312, 10), 1699 => to_unsigned(979, 10), 1700 => to_unsigned(798, 10), 1701 => to_unsigned(28, 10), 1702 => to_unsigned(96, 10), 1703 => to_unsigned(795, 10), 1704 => to_unsigned(303, 10), 1705 => to_unsigned(479, 10), 1706 => to_unsigned(830, 10), 1707 => to_unsigned(868, 10), 1708 => to_unsigned(740, 10), 1709 => to_unsigned(842, 10), 1710 => to_unsigned(361, 10), 1711 => to_unsigned(172, 10), 1712 => to_unsigned(802, 10), 1713 => to_unsigned(885, 10), 1714 => to_unsigned(574, 10), 1715 => to_unsigned(1003, 10), 1716 => to_unsigned(284, 10), 1717 => to_unsigned(204, 10), 1718 => to_unsigned(446, 10), 1719 => to_unsigned(187, 10), 1720 => to_unsigned(1019, 10), 1721 => to_unsigned(714, 10), 1722 => to_unsigned(904, 10), 1723 => to_unsigned(642, 10), 1724 => to_unsigned(61, 10), 1725 => to_unsigned(670, 10), 1726 => to_unsigned(114, 10), 1727 => to_unsigned(873, 10), 1728 => to_unsigned(203, 10), 1729 => to_unsigned(785, 10), 1730 => to_unsigned(405, 10), 1731 => to_unsigned(38, 10), 1732 => to_unsigned(208, 10), 1733 => to_unsigned(440, 10), 1734 => to_unsigned(594, 10), 1735 => to_unsigned(684, 10), 1736 => to_unsigned(805, 10), 1737 => to_unsigned(875, 10), 1738 => to_unsigned(472, 10), 1739 => to_unsigned(758, 10), 1740 => to_unsigned(428, 10), 1741 => to_unsigned(108, 10), 1742 => to_unsigned(841, 10), 1743 => to_unsigned(487, 10), 1744 => to_unsigned(229, 10), 1745 => to_unsigned(47, 10), 1746 => to_unsigned(112, 10), 1747 => to_unsigned(341, 10), 1748 => to_unsigned(595, 10), 1749 => to_unsigned(830, 10), 1750 => to_unsigned(636, 10), 1751 => to_unsigned(192, 10), 1752 => to_unsigned(46, 10), 1753 => to_unsigned(972, 10), 1754 => to_unsigned(155, 10), 1755 => to_unsigned(99, 10), 1756 => to_unsigned(305, 10), 1757 => to_unsigned(456, 10), 1758 => to_unsigned(460, 10), 1759 => to_unsigned(524, 10), 1760 => to_unsigned(368, 10), 1761 => to_unsigned(22, 10), 1762 => to_unsigned(97, 10), 1763 => to_unsigned(716, 10), 1764 => to_unsigned(702, 10), 1765 => to_unsigned(518, 10), 1766 => to_unsigned(1003, 10), 1767 => to_unsigned(469, 10), 1768 => to_unsigned(652, 10), 1769 => to_unsigned(853, 10), 1770 => to_unsigned(429, 10), 1771 => to_unsigned(140, 10), 1772 => to_unsigned(379, 10), 1773 => to_unsigned(363, 10), 1774 => to_unsigned(557, 10), 1775 => to_unsigned(174, 10), 1776 => to_unsigned(80, 10), 1777 => to_unsigned(925, 10), 1778 => to_unsigned(753, 10), 1779 => to_unsigned(669, 10), 1780 => to_unsigned(897, 10), 1781 => to_unsigned(126, 10), 1782 => to_unsigned(571, 10), 1783 => to_unsigned(994, 10), 1784 => to_unsigned(284, 10), 1785 => to_unsigned(182, 10), 1786 => to_unsigned(361, 10), 1787 => to_unsigned(677, 10), 1788 => to_unsigned(18, 10), 1789 => to_unsigned(92, 10), 1790 => to_unsigned(558, 10), 1791 => to_unsigned(464, 10), 1792 => to_unsigned(752, 10), 1793 => to_unsigned(356, 10), 1794 => to_unsigned(137, 10), 1795 => to_unsigned(921, 10), 1796 => to_unsigned(225, 10), 1797 => to_unsigned(536, 10), 1798 => to_unsigned(215, 10), 1799 => to_unsigned(637, 10), 1800 => to_unsigned(193, 10), 1801 => to_unsigned(108, 10), 1802 => to_unsigned(492, 10), 1803 => to_unsigned(456, 10), 1804 => to_unsigned(340, 10), 1805 => to_unsigned(734, 10), 1806 => to_unsigned(445, 10), 1807 => to_unsigned(283, 10), 1808 => to_unsigned(539, 10), 1809 => to_unsigned(555, 10), 1810 => to_unsigned(496, 10), 1811 => to_unsigned(460, 10), 1812 => to_unsigned(993, 10), 1813 => to_unsigned(689, 10), 1814 => to_unsigned(766, 10), 1815 => to_unsigned(329, 10), 1816 => to_unsigned(26, 10), 1817 => to_unsigned(173, 10), 1818 => to_unsigned(646, 10), 1819 => to_unsigned(462, 10), 1820 => to_unsigned(599, 10), 1821 => to_unsigned(201, 10), 1822 => to_unsigned(514, 10), 1823 => to_unsigned(369, 10), 1824 => to_unsigned(820, 10), 1825 => to_unsigned(868, 10), 1826 => to_unsigned(754, 10), 1827 => to_unsigned(996, 10), 1828 => to_unsigned(678, 10), 1829 => to_unsigned(814, 10), 1830 => to_unsigned(595, 10), 1831 => to_unsigned(702, 10), 1832 => to_unsigned(829, 10), 1833 => to_unsigned(924, 10), 1834 => to_unsigned(850, 10), 1835 => to_unsigned(948, 10), 1836 => to_unsigned(212, 10), 1837 => to_unsigned(254, 10), 1838 => to_unsigned(642, 10), 1839 => to_unsigned(64, 10), 1840 => to_unsigned(602, 10), 1841 => to_unsigned(476, 10), 1842 => to_unsigned(925, 10), 1843 => to_unsigned(126, 10), 1844 => to_unsigned(702, 10), 1845 => to_unsigned(296, 10), 1846 => to_unsigned(317, 10), 1847 => to_unsigned(706, 10), 1848 => to_unsigned(825, 10), 1849 => to_unsigned(11, 10), 1850 => to_unsigned(538, 10), 1851 => to_unsigned(300, 10), 1852 => to_unsigned(960, 10), 1853 => to_unsigned(414, 10), 1854 => to_unsigned(400, 10), 1855 => to_unsigned(565, 10), 1856 => to_unsigned(149, 10), 1857 => to_unsigned(712, 10), 1858 => to_unsigned(824, 10), 1859 => to_unsigned(1000, 10), 1860 => to_unsigned(395, 10), 1861 => to_unsigned(152, 10), 1862 => to_unsigned(122, 10), 1863 => to_unsigned(559, 10), 1864 => to_unsigned(819, 10), 1865 => to_unsigned(337, 10), 1866 => to_unsigned(932, 10), 1867 => to_unsigned(879, 10), 1868 => to_unsigned(184, 10), 1869 => to_unsigned(483, 10), 1870 => to_unsigned(524, 10), 1871 => to_unsigned(656, 10), 1872 => to_unsigned(148, 10), 1873 => to_unsigned(974, 10), 1874 => to_unsigned(415, 10), 1875 => to_unsigned(294, 10), 1876 => to_unsigned(866, 10), 1877 => to_unsigned(374, 10), 1878 => to_unsigned(484, 10), 1879 => to_unsigned(853, 10), 1880 => to_unsigned(978, 10), 1881 => to_unsigned(690, 10), 1882 => to_unsigned(929, 10), 1883 => to_unsigned(174, 10), 1884 => to_unsigned(576, 10), 1885 => to_unsigned(783, 10), 1886 => to_unsigned(895, 10), 1887 => to_unsigned(245, 10), 1888 => to_unsigned(989, 10), 1889 => to_unsigned(820, 10), 1890 => to_unsigned(856, 10), 1891 => to_unsigned(623, 10), 1892 => to_unsigned(314, 10), 1893 => to_unsigned(656, 10), 1894 => to_unsigned(498, 10), 1895 => to_unsigned(0, 10), 1896 => to_unsigned(499, 10), 1897 => to_unsigned(874, 10), 1898 => to_unsigned(920, 10), 1899 => to_unsigned(214, 10), 1900 => to_unsigned(985, 10), 1901 => to_unsigned(937, 10), 1902 => to_unsigned(235, 10), 1903 => to_unsigned(71, 10), 1904 => to_unsigned(769, 10), 1905 => to_unsigned(1011, 10), 1906 => to_unsigned(656, 10), 1907 => to_unsigned(718, 10), 1908 => to_unsigned(23, 10), 1909 => to_unsigned(125, 10), 1910 => to_unsigned(140, 10), 1911 => to_unsigned(565, 10), 1912 => to_unsigned(658, 10), 1913 => to_unsigned(105, 10), 1914 => to_unsigned(373, 10), 1915 => to_unsigned(594, 10), 1916 => to_unsigned(676, 10), 1917 => to_unsigned(212, 10), 1918 => to_unsigned(835, 10), 1919 => to_unsigned(612, 10), 1920 => to_unsigned(693, 10), 1921 => to_unsigned(183, 10), 1922 => to_unsigned(871, 10), 1923 => to_unsigned(145, 10), 1924 => to_unsigned(382, 10), 1925 => to_unsigned(371, 10), 1926 => to_unsigned(854, 10), 1927 => to_unsigned(210, 10), 1928 => to_unsigned(291, 10), 1929 => to_unsigned(996, 10), 1930 => to_unsigned(34, 10), 1931 => to_unsigned(1017, 10), 1932 => to_unsigned(516, 10), 1933 => to_unsigned(350, 10), 1934 => to_unsigned(554, 10), 1935 => to_unsigned(53, 10), 1936 => to_unsigned(353, 10), 1937 => to_unsigned(119, 10), 1938 => to_unsigned(487, 10), 1939 => to_unsigned(527, 10), 1940 => to_unsigned(283, 10), 1941 => to_unsigned(69, 10), 1942 => to_unsigned(343, 10), 1943 => to_unsigned(467, 10), 1944 => to_unsigned(633, 10), 1945 => to_unsigned(269, 10), 1946 => to_unsigned(119, 10), 1947 => to_unsigned(569, 10), 1948 => to_unsigned(788, 10), 1949 => to_unsigned(410, 10), 1950 => to_unsigned(351, 10), 1951 => to_unsigned(655, 10), 1952 => to_unsigned(465, 10), 1953 => to_unsigned(934, 10), 1954 => to_unsigned(338, 10), 1955 => to_unsigned(873, 10), 1956 => to_unsigned(934, 10), 1957 => to_unsigned(16, 10), 1958 => to_unsigned(217, 10), 1959 => to_unsigned(938, 10), 1960 => to_unsigned(269, 10), 1961 => to_unsigned(750, 10), 1962 => to_unsigned(303, 10), 1963 => to_unsigned(139, 10), 1964 => to_unsigned(555, 10), 1965 => to_unsigned(402, 10), 1966 => to_unsigned(657, 10), 1967 => to_unsigned(990, 10), 1968 => to_unsigned(356, 10), 1969 => to_unsigned(217, 10), 1970 => to_unsigned(5, 10), 1971 => to_unsigned(180, 10), 1972 => to_unsigned(88, 10), 1973 => to_unsigned(101, 10), 1974 => to_unsigned(437, 10), 1975 => to_unsigned(932, 10), 1976 => to_unsigned(515, 10), 1977 => to_unsigned(642, 10), 1978 => to_unsigned(988, 10), 1979 => to_unsigned(769, 10), 1980 => to_unsigned(787, 10), 1981 => to_unsigned(242, 10), 1982 => to_unsigned(797, 10), 1983 => to_unsigned(246, 10), 1984 => to_unsigned(553, 10), 1985 => to_unsigned(612, 10), 1986 => to_unsigned(562, 10), 1987 => to_unsigned(94, 10), 1988 => to_unsigned(940, 10), 1989 => to_unsigned(832, 10), 1990 => to_unsigned(95, 10), 1991 => to_unsigned(830, 10), 1992 => to_unsigned(894, 10), 1993 => to_unsigned(85, 10), 1994 => to_unsigned(475, 10), 1995 => to_unsigned(852, 10), 1996 => to_unsigned(496, 10), 1997 => to_unsigned(754, 10), 1998 => to_unsigned(323, 10), 1999 => to_unsigned(768, 10), 2000 => to_unsigned(748, 10), 2001 => to_unsigned(862, 10), 2002 => to_unsigned(303, 10), 2003 => to_unsigned(278, 10), 2004 => to_unsigned(200, 10), 2005 => to_unsigned(73, 10), 2006 => to_unsigned(102, 10), 2007 => to_unsigned(501, 10), 2008 => to_unsigned(220, 10), 2009 => to_unsigned(121, 10), 2010 => to_unsigned(135, 10), 2011 => to_unsigned(354, 10), 2012 => to_unsigned(172, 10), 2013 => to_unsigned(612, 10), 2014 => to_unsigned(875, 10), 2015 => to_unsigned(1021, 10), 2016 => to_unsigned(973, 10), 2017 => to_unsigned(730, 10), 2018 => to_unsigned(186, 10), 2019 => to_unsigned(656, 10), 2020 => to_unsigned(956, 10), 2021 => to_unsigned(371, 10), 2022 => to_unsigned(261, 10), 2023 => to_unsigned(302, 10), 2024 => to_unsigned(237, 10), 2025 => to_unsigned(1021, 10), 2026 => to_unsigned(109, 10), 2027 => to_unsigned(70, 10), 2028 => to_unsigned(682, 10), 2029 => to_unsigned(428, 10), 2030 => to_unsigned(717, 10), 2031 => to_unsigned(345, 10), 2032 => to_unsigned(406, 10), 2033 => to_unsigned(187, 10), 2034 => to_unsigned(844, 10), 2035 => to_unsigned(567, 10), 2036 => to_unsigned(152, 10), 2037 => to_unsigned(125, 10), 2038 => to_unsigned(772, 10), 2039 => to_unsigned(16, 10), 2040 => to_unsigned(444, 10), 2041 => to_unsigned(71, 10), 2042 => to_unsigned(548, 10), 2043 => to_unsigned(986, 10), 2044 => to_unsigned(473, 10), 2045 => to_unsigned(758, 10), 2046 => to_unsigned(189, 10), 2047 => to_unsigned(894, 10)),
            4 => (0 => to_unsigned(409, 10), 1 => to_unsigned(607, 10), 2 => to_unsigned(602, 10), 3 => to_unsigned(128, 10), 4 => to_unsigned(560, 10), 5 => to_unsigned(881, 10), 6 => to_unsigned(510, 10), 7 => to_unsigned(38, 10), 8 => to_unsigned(735, 10), 9 => to_unsigned(650, 10), 10 => to_unsigned(422, 10), 11 => to_unsigned(770, 10), 12 => to_unsigned(273, 10), 13 => to_unsigned(260, 10), 14 => to_unsigned(827, 10), 15 => to_unsigned(820, 10), 16 => to_unsigned(993, 10), 17 => to_unsigned(515, 10), 18 => to_unsigned(511, 10), 19 => to_unsigned(437, 10), 20 => to_unsigned(466, 10), 21 => to_unsigned(971, 10), 22 => to_unsigned(515, 10), 23 => to_unsigned(519, 10), 24 => to_unsigned(738, 10), 25 => to_unsigned(126, 10), 26 => to_unsigned(459, 10), 27 => to_unsigned(302, 10), 28 => to_unsigned(958, 10), 29 => to_unsigned(612, 10), 30 => to_unsigned(290, 10), 31 => to_unsigned(816, 10), 32 => to_unsigned(375, 10), 33 => to_unsigned(306, 10), 34 => to_unsigned(757, 10), 35 => to_unsigned(696, 10), 36 => to_unsigned(307, 10), 37 => to_unsigned(788, 10), 38 => to_unsigned(141, 10), 39 => to_unsigned(716, 10), 40 => to_unsigned(559, 10), 41 => to_unsigned(503, 10), 42 => to_unsigned(155, 10), 43 => to_unsigned(776, 10), 44 => to_unsigned(857, 10), 45 => to_unsigned(180, 10), 46 => to_unsigned(461, 10), 47 => to_unsigned(641, 10), 48 => to_unsigned(543, 10), 49 => to_unsigned(755, 10), 50 => to_unsigned(142, 10), 51 => to_unsigned(800, 10), 52 => to_unsigned(949, 10), 53 => to_unsigned(511, 10), 54 => to_unsigned(506, 10), 55 => to_unsigned(933, 10), 56 => to_unsigned(858, 10), 57 => to_unsigned(664, 10), 58 => to_unsigned(724, 10), 59 => to_unsigned(183, 10), 60 => to_unsigned(273, 10), 61 => to_unsigned(123, 10), 62 => to_unsigned(954, 10), 63 => to_unsigned(218, 10), 64 => to_unsigned(972, 10), 65 => to_unsigned(301, 10), 66 => to_unsigned(513, 10), 67 => to_unsigned(130, 10), 68 => to_unsigned(211, 10), 69 => to_unsigned(410, 10), 70 => to_unsigned(699, 10), 71 => to_unsigned(37, 10), 72 => to_unsigned(711, 10), 73 => to_unsigned(406, 10), 74 => to_unsigned(196, 10), 75 => to_unsigned(373, 10), 76 => to_unsigned(218, 10), 77 => to_unsigned(743, 10), 78 => to_unsigned(298, 10), 79 => to_unsigned(141, 10), 80 => to_unsigned(324, 10), 81 => to_unsigned(854, 10), 82 => to_unsigned(436, 10), 83 => to_unsigned(548, 10), 84 => to_unsigned(331, 10), 85 => to_unsigned(651, 10), 86 => to_unsigned(456, 10), 87 => to_unsigned(1015, 10), 88 => to_unsigned(942, 10), 89 => to_unsigned(43, 10), 90 => to_unsigned(819, 10), 91 => to_unsigned(102, 10), 92 => to_unsigned(616, 10), 93 => to_unsigned(360, 10), 94 => to_unsigned(123, 10), 95 => to_unsigned(732, 10), 96 => to_unsigned(606, 10), 97 => to_unsigned(215, 10), 98 => to_unsigned(270, 10), 99 => to_unsigned(250, 10), 100 => to_unsigned(319, 10), 101 => to_unsigned(159, 10), 102 => to_unsigned(702, 10), 103 => to_unsigned(214, 10), 104 => to_unsigned(362, 10), 105 => to_unsigned(657, 10), 106 => to_unsigned(244, 10), 107 => to_unsigned(110, 10), 108 => to_unsigned(719, 10), 109 => to_unsigned(628, 10), 110 => to_unsigned(306, 10), 111 => to_unsigned(804, 10), 112 => to_unsigned(333, 10), 113 => to_unsigned(961, 10), 114 => to_unsigned(264, 10), 115 => to_unsigned(445, 10), 116 => to_unsigned(254, 10), 117 => to_unsigned(525, 10), 118 => to_unsigned(720, 10), 119 => to_unsigned(529, 10), 120 => to_unsigned(845, 10), 121 => to_unsigned(764, 10), 122 => to_unsigned(826, 10), 123 => to_unsigned(530, 10), 124 => to_unsigned(1002, 10), 125 => to_unsigned(285, 10), 126 => to_unsigned(38, 10), 127 => to_unsigned(1005, 10), 128 => to_unsigned(910, 10), 129 => to_unsigned(431, 10), 130 => to_unsigned(357, 10), 131 => to_unsigned(820, 10), 132 => to_unsigned(495, 10), 133 => to_unsigned(423, 10), 134 => to_unsigned(1014, 10), 135 => to_unsigned(393, 10), 136 => to_unsigned(319, 10), 137 => to_unsigned(1013, 10), 138 => to_unsigned(775, 10), 139 => to_unsigned(977, 10), 140 => to_unsigned(958, 10), 141 => to_unsigned(225, 10), 142 => to_unsigned(924, 10), 143 => to_unsigned(581, 10), 144 => to_unsigned(992, 10), 145 => to_unsigned(362, 10), 146 => to_unsigned(719, 10), 147 => to_unsigned(53, 10), 148 => to_unsigned(769, 10), 149 => to_unsigned(789, 10), 150 => to_unsigned(424, 10), 151 => to_unsigned(516, 10), 152 => to_unsigned(484, 10), 153 => to_unsigned(229, 10), 154 => to_unsigned(1005, 10), 155 => to_unsigned(85, 10), 156 => to_unsigned(172, 10), 157 => to_unsigned(987, 10), 158 => to_unsigned(759, 10), 159 => to_unsigned(92, 10), 160 => to_unsigned(864, 10), 161 => to_unsigned(547, 10), 162 => to_unsigned(270, 10), 163 => to_unsigned(208, 10), 164 => to_unsigned(947, 10), 165 => to_unsigned(682, 10), 166 => to_unsigned(169, 10), 167 => to_unsigned(969, 10), 168 => to_unsigned(245, 10), 169 => to_unsigned(143, 10), 170 => to_unsigned(84, 10), 171 => to_unsigned(539, 10), 172 => to_unsigned(566, 10), 173 => to_unsigned(944, 10), 174 => to_unsigned(665, 10), 175 => to_unsigned(592, 10), 176 => to_unsigned(448, 10), 177 => to_unsigned(512, 10), 178 => to_unsigned(205, 10), 179 => to_unsigned(1017, 10), 180 => to_unsigned(355, 10), 181 => to_unsigned(1021, 10), 182 => to_unsigned(390, 10), 183 => to_unsigned(747, 10), 184 => to_unsigned(184, 10), 185 => to_unsigned(743, 10), 186 => to_unsigned(383, 10), 187 => to_unsigned(664, 10), 188 => to_unsigned(32, 10), 189 => to_unsigned(241, 10), 190 => to_unsigned(256, 10), 191 => to_unsigned(552, 10), 192 => to_unsigned(184, 10), 193 => to_unsigned(1014, 10), 194 => to_unsigned(228, 10), 195 => to_unsigned(550, 10), 196 => to_unsigned(697, 10), 197 => to_unsigned(205, 10), 198 => to_unsigned(771, 10), 199 => to_unsigned(678, 10), 200 => to_unsigned(713, 10), 201 => to_unsigned(60, 10), 202 => to_unsigned(396, 10), 203 => to_unsigned(246, 10), 204 => to_unsigned(588, 10), 205 => to_unsigned(34, 10), 206 => to_unsigned(846, 10), 207 => to_unsigned(231, 10), 208 => to_unsigned(973, 10), 209 => to_unsigned(255, 10), 210 => to_unsigned(868, 10), 211 => to_unsigned(517, 10), 212 => to_unsigned(320, 10), 213 => to_unsigned(621, 10), 214 => to_unsigned(782, 10), 215 => to_unsigned(409, 10), 216 => to_unsigned(474, 10), 217 => to_unsigned(879, 10), 218 => to_unsigned(179, 10), 219 => to_unsigned(1018, 10), 220 => to_unsigned(502, 10), 221 => to_unsigned(700, 10), 222 => to_unsigned(121, 10), 223 => to_unsigned(13, 10), 224 => to_unsigned(406, 10), 225 => to_unsigned(1018, 10), 226 => to_unsigned(355, 10), 227 => to_unsigned(78, 10), 228 => to_unsigned(464, 10), 229 => to_unsigned(782, 10), 230 => to_unsigned(123, 10), 231 => to_unsigned(145, 10), 232 => to_unsigned(593, 10), 233 => to_unsigned(772, 10), 234 => to_unsigned(380, 10), 235 => to_unsigned(52, 10), 236 => to_unsigned(400, 10), 237 => to_unsigned(573, 10), 238 => to_unsigned(802, 10), 239 => to_unsigned(610, 10), 240 => to_unsigned(771, 10), 241 => to_unsigned(380, 10), 242 => to_unsigned(333, 10), 243 => to_unsigned(520, 10), 244 => to_unsigned(483, 10), 245 => to_unsigned(315, 10), 246 => to_unsigned(192, 10), 247 => to_unsigned(795, 10), 248 => to_unsigned(347, 10), 249 => to_unsigned(73, 10), 250 => to_unsigned(705, 10), 251 => to_unsigned(682, 10), 252 => to_unsigned(999, 10), 253 => to_unsigned(803, 10), 254 => to_unsigned(931, 10), 255 => to_unsigned(229, 10), 256 => to_unsigned(739, 10), 257 => to_unsigned(664, 10), 258 => to_unsigned(790, 10), 259 => to_unsigned(485, 10), 260 => to_unsigned(537, 10), 261 => to_unsigned(196, 10), 262 => to_unsigned(13, 10), 263 => to_unsigned(894, 10), 264 => to_unsigned(333, 10), 265 => to_unsigned(342, 10), 266 => to_unsigned(938, 10), 267 => to_unsigned(150, 10), 268 => to_unsigned(680, 10), 269 => to_unsigned(999, 10), 270 => to_unsigned(291, 10), 271 => to_unsigned(524, 10), 272 => to_unsigned(400, 10), 273 => to_unsigned(471, 10), 274 => to_unsigned(956, 10), 275 => to_unsigned(451, 10), 276 => to_unsigned(714, 10), 277 => to_unsigned(423, 10), 278 => to_unsigned(394, 10), 279 => to_unsigned(273, 10), 280 => to_unsigned(343, 10), 281 => to_unsigned(279, 10), 282 => to_unsigned(826, 10), 283 => to_unsigned(478, 10), 284 => to_unsigned(663, 10), 285 => to_unsigned(731, 10), 286 => to_unsigned(10, 10), 287 => to_unsigned(532, 10), 288 => to_unsigned(9, 10), 289 => to_unsigned(261, 10), 290 => to_unsigned(862, 10), 291 => to_unsigned(733, 10), 292 => to_unsigned(91, 10), 293 => to_unsigned(914, 10), 294 => to_unsigned(755, 10), 295 => to_unsigned(327, 10), 296 => to_unsigned(106, 10), 297 => to_unsigned(846, 10), 298 => to_unsigned(640, 10), 299 => to_unsigned(1011, 10), 300 => to_unsigned(128, 10), 301 => to_unsigned(510, 10), 302 => to_unsigned(138, 10), 303 => to_unsigned(503, 10), 304 => to_unsigned(16, 10), 305 => to_unsigned(83, 10), 306 => to_unsigned(688, 10), 307 => to_unsigned(206, 10), 308 => to_unsigned(304, 10), 309 => to_unsigned(298, 10), 310 => to_unsigned(232, 10), 311 => to_unsigned(258, 10), 312 => to_unsigned(303, 10), 313 => to_unsigned(896, 10), 314 => to_unsigned(517, 10), 315 => to_unsigned(562, 10), 316 => to_unsigned(341, 10), 317 => to_unsigned(633, 10), 318 => to_unsigned(88, 10), 319 => to_unsigned(173, 10), 320 => to_unsigned(382, 10), 321 => to_unsigned(356, 10), 322 => to_unsigned(63, 10), 323 => to_unsigned(300, 10), 324 => to_unsigned(297, 10), 325 => to_unsigned(37, 10), 326 => to_unsigned(905, 10), 327 => to_unsigned(989, 10), 328 => to_unsigned(93, 10), 329 => to_unsigned(336, 10), 330 => to_unsigned(986, 10), 331 => to_unsigned(374, 10), 332 => to_unsigned(835, 10), 333 => to_unsigned(954, 10), 334 => to_unsigned(791, 10), 335 => to_unsigned(901, 10), 336 => to_unsigned(427, 10), 337 => to_unsigned(476, 10), 338 => to_unsigned(715, 10), 339 => to_unsigned(755, 10), 340 => to_unsigned(818, 10), 341 => to_unsigned(155, 10), 342 => to_unsigned(663, 10), 343 => to_unsigned(710, 10), 344 => to_unsigned(220, 10), 345 => to_unsigned(8, 10), 346 => to_unsigned(204, 10), 347 => to_unsigned(627, 10), 348 => to_unsigned(918, 10), 349 => to_unsigned(468, 10), 350 => to_unsigned(549, 10), 351 => to_unsigned(991, 10), 352 => to_unsigned(1015, 10), 353 => to_unsigned(353, 10), 354 => to_unsigned(773, 10), 355 => to_unsigned(159, 10), 356 => to_unsigned(737, 10), 357 => to_unsigned(264, 10), 358 => to_unsigned(827, 10), 359 => to_unsigned(416, 10), 360 => to_unsigned(950, 10), 361 => to_unsigned(958, 10), 362 => to_unsigned(705, 10), 363 => to_unsigned(954, 10), 364 => to_unsigned(530, 10), 365 => to_unsigned(221, 10), 366 => to_unsigned(622, 10), 367 => to_unsigned(349, 10), 368 => to_unsigned(474, 10), 369 => to_unsigned(621, 10), 370 => to_unsigned(581, 10), 371 => to_unsigned(453, 10), 372 => to_unsigned(673, 10), 373 => to_unsigned(184, 10), 374 => to_unsigned(38, 10), 375 => to_unsigned(0, 10), 376 => to_unsigned(622, 10), 377 => to_unsigned(404, 10), 378 => to_unsigned(111, 10), 379 => to_unsigned(939, 10), 380 => to_unsigned(737, 10), 381 => to_unsigned(398, 10), 382 => to_unsigned(423, 10), 383 => to_unsigned(950, 10), 384 => to_unsigned(450, 10), 385 => to_unsigned(109, 10), 386 => to_unsigned(795, 10), 387 => to_unsigned(648, 10), 388 => to_unsigned(165, 10), 389 => to_unsigned(19, 10), 390 => to_unsigned(834, 10), 391 => to_unsigned(647, 10), 392 => to_unsigned(547, 10), 393 => to_unsigned(621, 10), 394 => to_unsigned(818, 10), 395 => to_unsigned(871, 10), 396 => to_unsigned(782, 10), 397 => to_unsigned(33, 10), 398 => to_unsigned(967, 10), 399 => to_unsigned(183, 10), 400 => to_unsigned(691, 10), 401 => to_unsigned(629, 10), 402 => to_unsigned(373, 10), 403 => to_unsigned(144, 10), 404 => to_unsigned(24, 10), 405 => to_unsigned(926, 10), 406 => to_unsigned(486, 10), 407 => to_unsigned(556, 10), 408 => to_unsigned(391, 10), 409 => to_unsigned(175, 10), 410 => to_unsigned(101, 10), 411 => to_unsigned(745, 10), 412 => to_unsigned(1004, 10), 413 => to_unsigned(211, 10), 414 => to_unsigned(399, 10), 415 => to_unsigned(859, 10), 416 => to_unsigned(330, 10), 417 => to_unsigned(337, 10), 418 => to_unsigned(95, 10), 419 => to_unsigned(60, 10), 420 => to_unsigned(672, 10), 421 => to_unsigned(886, 10), 422 => to_unsigned(437, 10), 423 => to_unsigned(92, 10), 424 => to_unsigned(511, 10), 425 => to_unsigned(490, 10), 426 => to_unsigned(773, 10), 427 => to_unsigned(474, 10), 428 => to_unsigned(161, 10), 429 => to_unsigned(757, 10), 430 => to_unsigned(126, 10), 431 => to_unsigned(123, 10), 432 => to_unsigned(435, 10), 433 => to_unsigned(933, 10), 434 => to_unsigned(970, 10), 435 => to_unsigned(695, 10), 436 => to_unsigned(112, 10), 437 => to_unsigned(6, 10), 438 => to_unsigned(357, 10), 439 => to_unsigned(223, 10), 440 => to_unsigned(797, 10), 441 => to_unsigned(599, 10), 442 => to_unsigned(557, 10), 443 => to_unsigned(788, 10), 444 => to_unsigned(125, 10), 445 => to_unsigned(462, 10), 446 => to_unsigned(962, 10), 447 => to_unsigned(774, 10), 448 => to_unsigned(660, 10), 449 => to_unsigned(407, 10), 450 => to_unsigned(878, 10), 451 => to_unsigned(400, 10), 452 => to_unsigned(340, 10), 453 => to_unsigned(405, 10), 454 => to_unsigned(557, 10), 455 => to_unsigned(16, 10), 456 => to_unsigned(317, 10), 457 => to_unsigned(258, 10), 458 => to_unsigned(35, 10), 459 => to_unsigned(678, 10), 460 => to_unsigned(711, 10), 461 => to_unsigned(737, 10), 462 => to_unsigned(981, 10), 463 => to_unsigned(305, 10), 464 => to_unsigned(751, 10), 465 => to_unsigned(842, 10), 466 => to_unsigned(622, 10), 467 => to_unsigned(443, 10), 468 => to_unsigned(197, 10), 469 => to_unsigned(277, 10), 470 => to_unsigned(708, 10), 471 => to_unsigned(679, 10), 472 => to_unsigned(309, 10), 473 => to_unsigned(765, 10), 474 => to_unsigned(461, 10), 475 => to_unsigned(464, 10), 476 => to_unsigned(876, 10), 477 => to_unsigned(476, 10), 478 => to_unsigned(42, 10), 479 => to_unsigned(397, 10), 480 => to_unsigned(909, 10), 481 => to_unsigned(115, 10), 482 => to_unsigned(407, 10), 483 => to_unsigned(964, 10), 484 => to_unsigned(183, 10), 485 => to_unsigned(703, 10), 486 => to_unsigned(17, 10), 487 => to_unsigned(990, 10), 488 => to_unsigned(971, 10), 489 => to_unsigned(401, 10), 490 => to_unsigned(136, 10), 491 => to_unsigned(57, 10), 492 => to_unsigned(959, 10), 493 => to_unsigned(16, 10), 494 => to_unsigned(681, 10), 495 => to_unsigned(176, 10), 496 => to_unsigned(282, 10), 497 => to_unsigned(994, 10), 498 => to_unsigned(377, 10), 499 => to_unsigned(100, 10), 500 => to_unsigned(699, 10), 501 => to_unsigned(448, 10), 502 => to_unsigned(941, 10), 503 => to_unsigned(241, 10), 504 => to_unsigned(136, 10), 505 => to_unsigned(127, 10), 506 => to_unsigned(379, 10), 507 => to_unsigned(547, 10), 508 => to_unsigned(13, 10), 509 => to_unsigned(468, 10), 510 => to_unsigned(865, 10), 511 => to_unsigned(849, 10), 512 => to_unsigned(954, 10), 513 => to_unsigned(70, 10), 514 => to_unsigned(364, 10), 515 => to_unsigned(273, 10), 516 => to_unsigned(605, 10), 517 => to_unsigned(930, 10), 518 => to_unsigned(415, 10), 519 => to_unsigned(84, 10), 520 => to_unsigned(87, 10), 521 => to_unsigned(488, 10), 522 => to_unsigned(984, 10), 523 => to_unsigned(459, 10), 524 => to_unsigned(809, 10), 525 => to_unsigned(466, 10), 526 => to_unsigned(73, 10), 527 => to_unsigned(969, 10), 528 => to_unsigned(625, 10), 529 => to_unsigned(636, 10), 530 => to_unsigned(285, 10), 531 => to_unsigned(993, 10), 532 => to_unsigned(238, 10), 533 => to_unsigned(635, 10), 534 => to_unsigned(223, 10), 535 => to_unsigned(982, 10), 536 => to_unsigned(89, 10), 537 => to_unsigned(702, 10), 538 => to_unsigned(5, 10), 539 => to_unsigned(637, 10), 540 => to_unsigned(296, 10), 541 => to_unsigned(547, 10), 542 => to_unsigned(813, 10), 543 => to_unsigned(274, 10), 544 => to_unsigned(214, 10), 545 => to_unsigned(865, 10), 546 => to_unsigned(974, 10), 547 => to_unsigned(737, 10), 548 => to_unsigned(871, 10), 549 => to_unsigned(678, 10), 550 => to_unsigned(389, 10), 551 => to_unsigned(769, 10), 552 => to_unsigned(5, 10), 553 => to_unsigned(486, 10), 554 => to_unsigned(799, 10), 555 => to_unsigned(481, 10), 556 => to_unsigned(168, 10), 557 => to_unsigned(364, 10), 558 => to_unsigned(129, 10), 559 => to_unsigned(468, 10), 560 => to_unsigned(870, 10), 561 => to_unsigned(111, 10), 562 => to_unsigned(423, 10), 563 => to_unsigned(724, 10), 564 => to_unsigned(781, 10), 565 => to_unsigned(427, 10), 566 => to_unsigned(83, 10), 567 => to_unsigned(491, 10), 568 => to_unsigned(409, 10), 569 => to_unsigned(312, 10), 570 => to_unsigned(884, 10), 571 => to_unsigned(572, 10), 572 => to_unsigned(316, 10), 573 => to_unsigned(257, 10), 574 => to_unsigned(748, 10), 575 => to_unsigned(5, 10), 576 => to_unsigned(5, 10), 577 => to_unsigned(472, 10), 578 => to_unsigned(858, 10), 579 => to_unsigned(121, 10), 580 => to_unsigned(604, 10), 581 => to_unsigned(290, 10), 582 => to_unsigned(756, 10), 583 => to_unsigned(24, 10), 584 => to_unsigned(340, 10), 585 => to_unsigned(1006, 10), 586 => to_unsigned(977, 10), 587 => to_unsigned(823, 10), 588 => to_unsigned(1008, 10), 589 => to_unsigned(571, 10), 590 => to_unsigned(640, 10), 591 => to_unsigned(290, 10), 592 => to_unsigned(478, 10), 593 => to_unsigned(755, 10), 594 => to_unsigned(902, 10), 595 => to_unsigned(952, 10), 596 => to_unsigned(238, 10), 597 => to_unsigned(68, 10), 598 => to_unsigned(264, 10), 599 => to_unsigned(275, 10), 600 => to_unsigned(323, 10), 601 => to_unsigned(416, 10), 602 => to_unsigned(383, 10), 603 => to_unsigned(579, 10), 604 => to_unsigned(615, 10), 605 => to_unsigned(61, 10), 606 => to_unsigned(922, 10), 607 => to_unsigned(147, 10), 608 => to_unsigned(204, 10), 609 => to_unsigned(896, 10), 610 => to_unsigned(981, 10), 611 => to_unsigned(980, 10), 612 => to_unsigned(817, 10), 613 => to_unsigned(379, 10), 614 => to_unsigned(106, 10), 615 => to_unsigned(578, 10), 616 => to_unsigned(256, 10), 617 => to_unsigned(401, 10), 618 => to_unsigned(544, 10), 619 => to_unsigned(176, 10), 620 => to_unsigned(802, 10), 621 => to_unsigned(105, 10), 622 => to_unsigned(901, 10), 623 => to_unsigned(422, 10), 624 => to_unsigned(306, 10), 625 => to_unsigned(530, 10), 626 => to_unsigned(696, 10), 627 => to_unsigned(850, 10), 628 => to_unsigned(224, 10), 629 => to_unsigned(166, 10), 630 => to_unsigned(728, 10), 631 => to_unsigned(960, 10), 632 => to_unsigned(392, 10), 633 => to_unsigned(353, 10), 634 => to_unsigned(899, 10), 635 => to_unsigned(684, 10), 636 => to_unsigned(428, 10), 637 => to_unsigned(434, 10), 638 => to_unsigned(571, 10), 639 => to_unsigned(252, 10), 640 => to_unsigned(459, 10), 641 => to_unsigned(568, 10), 642 => to_unsigned(513, 10), 643 => to_unsigned(553, 10), 644 => to_unsigned(26, 10), 645 => to_unsigned(856, 10), 646 => to_unsigned(1012, 10), 647 => to_unsigned(443, 10), 648 => to_unsigned(125, 10), 649 => to_unsigned(406, 10), 650 => to_unsigned(639, 10), 651 => to_unsigned(1005, 10), 652 => to_unsigned(495, 10), 653 => to_unsigned(452, 10), 654 => to_unsigned(397, 10), 655 => to_unsigned(1014, 10), 656 => to_unsigned(308, 10), 657 => to_unsigned(100, 10), 658 => to_unsigned(722, 10), 659 => to_unsigned(701, 10), 660 => to_unsigned(810, 10), 661 => to_unsigned(857, 10), 662 => to_unsigned(896, 10), 663 => to_unsigned(513, 10), 664 => to_unsigned(28, 10), 665 => to_unsigned(787, 10), 666 => to_unsigned(159, 10), 667 => to_unsigned(532, 10), 668 => to_unsigned(755, 10), 669 => to_unsigned(684, 10), 670 => to_unsigned(779, 10), 671 => to_unsigned(915, 10), 672 => to_unsigned(168, 10), 673 => to_unsigned(991, 10), 674 => to_unsigned(953, 10), 675 => to_unsigned(393, 10), 676 => to_unsigned(249, 10), 677 => to_unsigned(847, 10), 678 => to_unsigned(929, 10), 679 => to_unsigned(372, 10), 680 => to_unsigned(660, 10), 681 => to_unsigned(776, 10), 682 => to_unsigned(453, 10), 683 => to_unsigned(207, 10), 684 => to_unsigned(722, 10), 685 => to_unsigned(777, 10), 686 => to_unsigned(700, 10), 687 => to_unsigned(6, 10), 688 => to_unsigned(435, 10), 689 => to_unsigned(130, 10), 690 => to_unsigned(781, 10), 691 => to_unsigned(534, 10), 692 => to_unsigned(895, 10), 693 => to_unsigned(950, 10), 694 => to_unsigned(898, 10), 695 => to_unsigned(567, 10), 696 => to_unsigned(377, 10), 697 => to_unsigned(344, 10), 698 => to_unsigned(303, 10), 699 => to_unsigned(177, 10), 700 => to_unsigned(476, 10), 701 => to_unsigned(809, 10), 702 => to_unsigned(425, 10), 703 => to_unsigned(438, 10), 704 => to_unsigned(28, 10), 705 => to_unsigned(468, 10), 706 => to_unsigned(856, 10), 707 => to_unsigned(199, 10), 708 => to_unsigned(269, 10), 709 => to_unsigned(877, 10), 710 => to_unsigned(242, 10), 711 => to_unsigned(111, 10), 712 => to_unsigned(570, 10), 713 => to_unsigned(243, 10), 714 => to_unsigned(1013, 10), 715 => to_unsigned(342, 10), 716 => to_unsigned(622, 10), 717 => to_unsigned(726, 10), 718 => to_unsigned(805, 10), 719 => to_unsigned(209, 10), 720 => to_unsigned(255, 10), 721 => to_unsigned(149, 10), 722 => to_unsigned(532, 10), 723 => to_unsigned(950, 10), 724 => to_unsigned(66, 10), 725 => to_unsigned(621, 10), 726 => to_unsigned(333, 10), 727 => to_unsigned(47, 10), 728 => to_unsigned(778, 10), 729 => to_unsigned(770, 10), 730 => to_unsigned(763, 10), 731 => to_unsigned(646, 10), 732 => to_unsigned(335, 10), 733 => to_unsigned(325, 10), 734 => to_unsigned(144, 10), 735 => to_unsigned(718, 10), 736 => to_unsigned(554, 10), 737 => to_unsigned(795, 10), 738 => to_unsigned(904, 10), 739 => to_unsigned(109, 10), 740 => to_unsigned(940, 10), 741 => to_unsigned(69, 10), 742 => to_unsigned(956, 10), 743 => to_unsigned(329, 10), 744 => to_unsigned(383, 10), 745 => to_unsigned(307, 10), 746 => to_unsigned(931, 10), 747 => to_unsigned(712, 10), 748 => to_unsigned(549, 10), 749 => to_unsigned(690, 10), 750 => to_unsigned(388, 10), 751 => to_unsigned(1015, 10), 752 => to_unsigned(708, 10), 753 => to_unsigned(871, 10), 754 => to_unsigned(957, 10), 755 => to_unsigned(557, 10), 756 => to_unsigned(302, 10), 757 => to_unsigned(820, 10), 758 => to_unsigned(184, 10), 759 => to_unsigned(587, 10), 760 => to_unsigned(660, 10), 761 => to_unsigned(392, 10), 762 => to_unsigned(377, 10), 763 => to_unsigned(736, 10), 764 => to_unsigned(418, 10), 765 => to_unsigned(875, 10), 766 => to_unsigned(613, 10), 767 => to_unsigned(532, 10), 768 => to_unsigned(51, 10), 769 => to_unsigned(851, 10), 770 => to_unsigned(63, 10), 771 => to_unsigned(644, 10), 772 => to_unsigned(42, 10), 773 => to_unsigned(301, 10), 774 => to_unsigned(929, 10), 775 => to_unsigned(625, 10), 776 => to_unsigned(975, 10), 777 => to_unsigned(241, 10), 778 => to_unsigned(996, 10), 779 => to_unsigned(823, 10), 780 => to_unsigned(88, 10), 781 => to_unsigned(36, 10), 782 => to_unsigned(215, 10), 783 => to_unsigned(352, 10), 784 => to_unsigned(55, 10), 785 => to_unsigned(1005, 10), 786 => to_unsigned(476, 10), 787 => to_unsigned(130, 10), 788 => to_unsigned(134, 10), 789 => to_unsigned(66, 10), 790 => to_unsigned(555, 10), 791 => to_unsigned(919, 10), 792 => to_unsigned(719, 10), 793 => to_unsigned(686, 10), 794 => to_unsigned(987, 10), 795 => to_unsigned(494, 10), 796 => to_unsigned(307, 10), 797 => to_unsigned(963, 10), 798 => to_unsigned(427, 10), 799 => to_unsigned(989, 10), 800 => to_unsigned(620, 10), 801 => to_unsigned(118, 10), 802 => to_unsigned(745, 10), 803 => to_unsigned(573, 10), 804 => to_unsigned(130, 10), 805 => to_unsigned(854, 10), 806 => to_unsigned(320, 10), 807 => to_unsigned(948, 10), 808 => to_unsigned(447, 10), 809 => to_unsigned(183, 10), 810 => to_unsigned(313, 10), 811 => to_unsigned(172, 10), 812 => to_unsigned(241, 10), 813 => to_unsigned(1010, 10), 814 => to_unsigned(832, 10), 815 => to_unsigned(993, 10), 816 => to_unsigned(463, 10), 817 => to_unsigned(314, 10), 818 => to_unsigned(646, 10), 819 => to_unsigned(498, 10), 820 => to_unsigned(449, 10), 821 => to_unsigned(0, 10), 822 => to_unsigned(85, 10), 823 => to_unsigned(368, 10), 824 => to_unsigned(785, 10), 825 => to_unsigned(1018, 10), 826 => to_unsigned(774, 10), 827 => to_unsigned(62, 10), 828 => to_unsigned(184, 10), 829 => to_unsigned(588, 10), 830 => to_unsigned(9, 10), 831 => to_unsigned(14, 10), 832 => to_unsigned(966, 10), 833 => to_unsigned(506, 10), 834 => to_unsigned(626, 10), 835 => to_unsigned(479, 10), 836 => to_unsigned(705, 10), 837 => to_unsigned(478, 10), 838 => to_unsigned(820, 10), 839 => to_unsigned(352, 10), 840 => to_unsigned(152, 10), 841 => to_unsigned(739, 10), 842 => to_unsigned(971, 10), 843 => to_unsigned(276, 10), 844 => to_unsigned(578, 10), 845 => to_unsigned(242, 10), 846 => to_unsigned(696, 10), 847 => to_unsigned(844, 10), 848 => to_unsigned(240, 10), 849 => to_unsigned(785, 10), 850 => to_unsigned(20, 10), 851 => to_unsigned(111, 10), 852 => to_unsigned(224, 10), 853 => to_unsigned(577, 10), 854 => to_unsigned(65, 10), 855 => to_unsigned(610, 10), 856 => to_unsigned(711, 10), 857 => to_unsigned(306, 10), 858 => to_unsigned(445, 10), 859 => to_unsigned(407, 10), 860 => to_unsigned(359, 10), 861 => to_unsigned(321, 10), 862 => to_unsigned(360, 10), 863 => to_unsigned(689, 10), 864 => to_unsigned(854, 10), 865 => to_unsigned(653, 10), 866 => to_unsigned(40, 10), 867 => to_unsigned(906, 10), 868 => to_unsigned(101, 10), 869 => to_unsigned(194, 10), 870 => to_unsigned(815, 10), 871 => to_unsigned(613, 10), 872 => to_unsigned(834, 10), 873 => to_unsigned(287, 10), 874 => to_unsigned(48, 10), 875 => to_unsigned(675, 10), 876 => to_unsigned(667, 10), 877 => to_unsigned(217, 10), 878 => to_unsigned(266, 10), 879 => to_unsigned(358, 10), 880 => to_unsigned(742, 10), 881 => to_unsigned(554, 10), 882 => to_unsigned(472, 10), 883 => to_unsigned(286, 10), 884 => to_unsigned(121, 10), 885 => to_unsigned(314, 10), 886 => to_unsigned(778, 10), 887 => to_unsigned(45, 10), 888 => to_unsigned(874, 10), 889 => to_unsigned(1018, 10), 890 => to_unsigned(387, 10), 891 => to_unsigned(902, 10), 892 => to_unsigned(313, 10), 893 => to_unsigned(9, 10), 894 => to_unsigned(299, 10), 895 => to_unsigned(385, 10), 896 => to_unsigned(585, 10), 897 => to_unsigned(561, 10), 898 => to_unsigned(857, 10), 899 => to_unsigned(464, 10), 900 => to_unsigned(775, 10), 901 => to_unsigned(232, 10), 902 => to_unsigned(235, 10), 903 => to_unsigned(897, 10), 904 => to_unsigned(59, 10), 905 => to_unsigned(576, 10), 906 => to_unsigned(343, 10), 907 => to_unsigned(115, 10), 908 => to_unsigned(47, 10), 909 => to_unsigned(174, 10), 910 => to_unsigned(26, 10), 911 => to_unsigned(562, 10), 912 => to_unsigned(306, 10), 913 => to_unsigned(212, 10), 914 => to_unsigned(43, 10), 915 => to_unsigned(408, 10), 916 => to_unsigned(682, 10), 917 => to_unsigned(198, 10), 918 => to_unsigned(596, 10), 919 => to_unsigned(47, 10), 920 => to_unsigned(369, 10), 921 => to_unsigned(121, 10), 922 => to_unsigned(875, 10), 923 => to_unsigned(484, 10), 924 => to_unsigned(389, 10), 925 => to_unsigned(238, 10), 926 => to_unsigned(308, 10), 927 => to_unsigned(327, 10), 928 => to_unsigned(28, 10), 929 => to_unsigned(54, 10), 930 => to_unsigned(904, 10), 931 => to_unsigned(623, 10), 932 => to_unsigned(743, 10), 933 => to_unsigned(502, 10), 934 => to_unsigned(800, 10), 935 => to_unsigned(526, 10), 936 => to_unsigned(721, 10), 937 => to_unsigned(412, 10), 938 => to_unsigned(837, 10), 939 => to_unsigned(502, 10), 940 => to_unsigned(861, 10), 941 => to_unsigned(557, 10), 942 => to_unsigned(173, 10), 943 => to_unsigned(616, 10), 944 => to_unsigned(531, 10), 945 => to_unsigned(974, 10), 946 => to_unsigned(45, 10), 947 => to_unsigned(88, 10), 948 => to_unsigned(455, 10), 949 => to_unsigned(890, 10), 950 => to_unsigned(760, 10), 951 => to_unsigned(111, 10), 952 => to_unsigned(78, 10), 953 => to_unsigned(858, 10), 954 => to_unsigned(415, 10), 955 => to_unsigned(397, 10), 956 => to_unsigned(478, 10), 957 => to_unsigned(646, 10), 958 => to_unsigned(316, 10), 959 => to_unsigned(437, 10), 960 => to_unsigned(637, 10), 961 => to_unsigned(994, 10), 962 => to_unsigned(998, 10), 963 => to_unsigned(236, 10), 964 => to_unsigned(642, 10), 965 => to_unsigned(549, 10), 966 => to_unsigned(743, 10), 967 => to_unsigned(385, 10), 968 => to_unsigned(890, 10), 969 => to_unsigned(385, 10), 970 => to_unsigned(790, 10), 971 => to_unsigned(816, 10), 972 => to_unsigned(682, 10), 973 => to_unsigned(891, 10), 974 => to_unsigned(494, 10), 975 => to_unsigned(878, 10), 976 => to_unsigned(755, 10), 977 => to_unsigned(121, 10), 978 => to_unsigned(522, 10), 979 => to_unsigned(462, 10), 980 => to_unsigned(244, 10), 981 => to_unsigned(533, 10), 982 => to_unsigned(949, 10), 983 => to_unsigned(679, 10), 984 => to_unsigned(987, 10), 985 => to_unsigned(855, 10), 986 => to_unsigned(702, 10), 987 => to_unsigned(116, 10), 988 => to_unsigned(574, 10), 989 => to_unsigned(512, 10), 990 => to_unsigned(357, 10), 991 => to_unsigned(263, 10), 992 => to_unsigned(779, 10), 993 => to_unsigned(503, 10), 994 => to_unsigned(879, 10), 995 => to_unsigned(387, 10), 996 => to_unsigned(339, 10), 997 => to_unsigned(416, 10), 998 => to_unsigned(621, 10), 999 => to_unsigned(1000, 10), 1000 => to_unsigned(1008, 10), 1001 => to_unsigned(51, 10), 1002 => to_unsigned(327, 10), 1003 => to_unsigned(871, 10), 1004 => to_unsigned(392, 10), 1005 => to_unsigned(266, 10), 1006 => to_unsigned(853, 10), 1007 => to_unsigned(740, 10), 1008 => to_unsigned(717, 10), 1009 => to_unsigned(990, 10), 1010 => to_unsigned(861, 10), 1011 => to_unsigned(880, 10), 1012 => to_unsigned(794, 10), 1013 => to_unsigned(126, 10), 1014 => to_unsigned(520, 10), 1015 => to_unsigned(979, 10), 1016 => to_unsigned(958, 10), 1017 => to_unsigned(790, 10), 1018 => to_unsigned(559, 10), 1019 => to_unsigned(298, 10), 1020 => to_unsigned(490, 10), 1021 => to_unsigned(10, 10), 1022 => to_unsigned(538, 10), 1023 => to_unsigned(538, 10), 1024 => to_unsigned(25, 10), 1025 => to_unsigned(708, 10), 1026 => to_unsigned(485, 10), 1027 => to_unsigned(422, 10), 1028 => to_unsigned(786, 10), 1029 => to_unsigned(370, 10), 1030 => to_unsigned(991, 10), 1031 => to_unsigned(636, 10), 1032 => to_unsigned(952, 10), 1033 => to_unsigned(79, 10), 1034 => to_unsigned(172, 10), 1035 => to_unsigned(750, 10), 1036 => to_unsigned(986, 10), 1037 => to_unsigned(699, 10), 1038 => to_unsigned(514, 10), 1039 => to_unsigned(25, 10), 1040 => to_unsigned(417, 10), 1041 => to_unsigned(513, 10), 1042 => to_unsigned(437, 10), 1043 => to_unsigned(908, 10), 1044 => to_unsigned(705, 10), 1045 => to_unsigned(125, 10), 1046 => to_unsigned(331, 10), 1047 => to_unsigned(257, 10), 1048 => to_unsigned(323, 10), 1049 => to_unsigned(146, 10), 1050 => to_unsigned(31, 10), 1051 => to_unsigned(631, 10), 1052 => to_unsigned(138, 10), 1053 => to_unsigned(639, 10), 1054 => to_unsigned(193, 10), 1055 => to_unsigned(63, 10), 1056 => to_unsigned(512, 10), 1057 => to_unsigned(140, 10), 1058 => to_unsigned(340, 10), 1059 => to_unsigned(282, 10), 1060 => to_unsigned(346, 10), 1061 => to_unsigned(321, 10), 1062 => to_unsigned(695, 10), 1063 => to_unsigned(184, 10), 1064 => to_unsigned(118, 10), 1065 => to_unsigned(676, 10), 1066 => to_unsigned(764, 10), 1067 => to_unsigned(423, 10), 1068 => to_unsigned(819, 10), 1069 => to_unsigned(310, 10), 1070 => to_unsigned(784, 10), 1071 => to_unsigned(444, 10), 1072 => to_unsigned(693, 10), 1073 => to_unsigned(993, 10), 1074 => to_unsigned(925, 10), 1075 => to_unsigned(574, 10), 1076 => to_unsigned(1009, 10), 1077 => to_unsigned(612, 10), 1078 => to_unsigned(340, 10), 1079 => to_unsigned(510, 10), 1080 => to_unsigned(425, 10), 1081 => to_unsigned(858, 10), 1082 => to_unsigned(327, 10), 1083 => to_unsigned(560, 10), 1084 => to_unsigned(889, 10), 1085 => to_unsigned(797, 10), 1086 => to_unsigned(814, 10), 1087 => to_unsigned(968, 10), 1088 => to_unsigned(925, 10), 1089 => to_unsigned(591, 10), 1090 => to_unsigned(60, 10), 1091 => to_unsigned(208, 10), 1092 => to_unsigned(734, 10), 1093 => to_unsigned(265, 10), 1094 => to_unsigned(93, 10), 1095 => to_unsigned(411, 10), 1096 => to_unsigned(95, 10), 1097 => to_unsigned(5, 10), 1098 => to_unsigned(981, 10), 1099 => to_unsigned(140, 10), 1100 => to_unsigned(592, 10), 1101 => to_unsigned(268, 10), 1102 => to_unsigned(184, 10), 1103 => to_unsigned(889, 10), 1104 => to_unsigned(751, 10), 1105 => to_unsigned(284, 10), 1106 => to_unsigned(329, 10), 1107 => to_unsigned(153, 10), 1108 => to_unsigned(872, 10), 1109 => to_unsigned(548, 10), 1110 => to_unsigned(676, 10), 1111 => to_unsigned(548, 10), 1112 => to_unsigned(814, 10), 1113 => to_unsigned(811, 10), 1114 => to_unsigned(60, 10), 1115 => to_unsigned(1013, 10), 1116 => to_unsigned(721, 10), 1117 => to_unsigned(24, 10), 1118 => to_unsigned(855, 10), 1119 => to_unsigned(756, 10), 1120 => to_unsigned(659, 10), 1121 => to_unsigned(462, 10), 1122 => to_unsigned(923, 10), 1123 => to_unsigned(855, 10), 1124 => to_unsigned(270, 10), 1125 => to_unsigned(169, 10), 1126 => to_unsigned(235, 10), 1127 => to_unsigned(400, 10), 1128 => to_unsigned(349, 10), 1129 => to_unsigned(28, 10), 1130 => to_unsigned(751, 10), 1131 => to_unsigned(332, 10), 1132 => to_unsigned(576, 10), 1133 => to_unsigned(1003, 10), 1134 => to_unsigned(551, 10), 1135 => to_unsigned(859, 10), 1136 => to_unsigned(84, 10), 1137 => to_unsigned(595, 10), 1138 => to_unsigned(392, 10), 1139 => to_unsigned(709, 10), 1140 => to_unsigned(7, 10), 1141 => to_unsigned(478, 10), 1142 => to_unsigned(386, 10), 1143 => to_unsigned(227, 10), 1144 => to_unsigned(584, 10), 1145 => to_unsigned(144, 10), 1146 => to_unsigned(656, 10), 1147 => to_unsigned(103, 10), 1148 => to_unsigned(7, 10), 1149 => to_unsigned(744, 10), 1150 => to_unsigned(619, 10), 1151 => to_unsigned(186, 10), 1152 => to_unsigned(576, 10), 1153 => to_unsigned(726, 10), 1154 => to_unsigned(612, 10), 1155 => to_unsigned(305, 10), 1156 => to_unsigned(628, 10), 1157 => to_unsigned(1009, 10), 1158 => to_unsigned(677, 10), 1159 => to_unsigned(57, 10), 1160 => to_unsigned(57, 10), 1161 => to_unsigned(1017, 10), 1162 => to_unsigned(845, 10), 1163 => to_unsigned(890, 10), 1164 => to_unsigned(554, 10), 1165 => to_unsigned(839, 10), 1166 => to_unsigned(953, 10), 1167 => to_unsigned(645, 10), 1168 => to_unsigned(37, 10), 1169 => to_unsigned(939, 10), 1170 => to_unsigned(13, 10), 1171 => to_unsigned(126, 10), 1172 => to_unsigned(35, 10), 1173 => to_unsigned(407, 10), 1174 => to_unsigned(570, 10), 1175 => to_unsigned(782, 10), 1176 => to_unsigned(297, 10), 1177 => to_unsigned(703, 10), 1178 => to_unsigned(767, 10), 1179 => to_unsigned(965, 10), 1180 => to_unsigned(405, 10), 1181 => to_unsigned(109, 10), 1182 => to_unsigned(922, 10), 1183 => to_unsigned(474, 10), 1184 => to_unsigned(621, 10), 1185 => to_unsigned(10, 10), 1186 => to_unsigned(428, 10), 1187 => to_unsigned(871, 10), 1188 => to_unsigned(409, 10), 1189 => to_unsigned(7, 10), 1190 => to_unsigned(63, 10), 1191 => to_unsigned(954, 10), 1192 => to_unsigned(818, 10), 1193 => to_unsigned(853, 10), 1194 => to_unsigned(938, 10), 1195 => to_unsigned(457, 10), 1196 => to_unsigned(364, 10), 1197 => to_unsigned(604, 10), 1198 => to_unsigned(653, 10), 1199 => to_unsigned(505, 10), 1200 => to_unsigned(831, 10), 1201 => to_unsigned(751, 10), 1202 => to_unsigned(231, 10), 1203 => to_unsigned(880, 10), 1204 => to_unsigned(396, 10), 1205 => to_unsigned(591, 10), 1206 => to_unsigned(59, 10), 1207 => to_unsigned(420, 10), 1208 => to_unsigned(61, 10), 1209 => to_unsigned(73, 10), 1210 => to_unsigned(710, 10), 1211 => to_unsigned(300, 10), 1212 => to_unsigned(436, 10), 1213 => to_unsigned(469, 10), 1214 => to_unsigned(551, 10), 1215 => to_unsigned(790, 10), 1216 => to_unsigned(204, 10), 1217 => to_unsigned(420, 10), 1218 => to_unsigned(730, 10), 1219 => to_unsigned(931, 10), 1220 => to_unsigned(1011, 10), 1221 => to_unsigned(984, 10), 1222 => to_unsigned(136, 10), 1223 => to_unsigned(513, 10), 1224 => to_unsigned(687, 10), 1225 => to_unsigned(407, 10), 1226 => to_unsigned(430, 10), 1227 => to_unsigned(1004, 10), 1228 => to_unsigned(30, 10), 1229 => to_unsigned(902, 10), 1230 => to_unsigned(394, 10), 1231 => to_unsigned(325, 10), 1232 => to_unsigned(981, 10), 1233 => to_unsigned(171, 10), 1234 => to_unsigned(836, 10), 1235 => to_unsigned(321, 10), 1236 => to_unsigned(759, 10), 1237 => to_unsigned(424, 10), 1238 => to_unsigned(430, 10), 1239 => to_unsigned(956, 10), 1240 => to_unsigned(946, 10), 1241 => to_unsigned(76, 10), 1242 => to_unsigned(754, 10), 1243 => to_unsigned(707, 10), 1244 => to_unsigned(630, 10), 1245 => to_unsigned(980, 10), 1246 => to_unsigned(360, 10), 1247 => to_unsigned(695, 10), 1248 => to_unsigned(526, 10), 1249 => to_unsigned(459, 10), 1250 => to_unsigned(840, 10), 1251 => to_unsigned(13, 10), 1252 => to_unsigned(226, 10), 1253 => to_unsigned(675, 10), 1254 => to_unsigned(774, 10), 1255 => to_unsigned(633, 10), 1256 => to_unsigned(328, 10), 1257 => to_unsigned(846, 10), 1258 => to_unsigned(96, 10), 1259 => to_unsigned(881, 10), 1260 => to_unsigned(721, 10), 1261 => to_unsigned(929, 10), 1262 => to_unsigned(371, 10), 1263 => to_unsigned(1018, 10), 1264 => to_unsigned(849, 10), 1265 => to_unsigned(860, 10), 1266 => to_unsigned(210, 10), 1267 => to_unsigned(20, 10), 1268 => to_unsigned(1000, 10), 1269 => to_unsigned(5, 10), 1270 => to_unsigned(601, 10), 1271 => to_unsigned(862, 10), 1272 => to_unsigned(33, 10), 1273 => to_unsigned(994, 10), 1274 => to_unsigned(430, 10), 1275 => to_unsigned(799, 10), 1276 => to_unsigned(269, 10), 1277 => to_unsigned(591, 10), 1278 => to_unsigned(697, 10), 1279 => to_unsigned(324, 10), 1280 => to_unsigned(693, 10), 1281 => to_unsigned(509, 10), 1282 => to_unsigned(890, 10), 1283 => to_unsigned(985, 10), 1284 => to_unsigned(30, 10), 1285 => to_unsigned(591, 10), 1286 => to_unsigned(638, 10), 1287 => to_unsigned(877, 10), 1288 => to_unsigned(922, 10), 1289 => to_unsigned(244, 10), 1290 => to_unsigned(206, 10), 1291 => to_unsigned(1005, 10), 1292 => to_unsigned(957, 10), 1293 => to_unsigned(68, 10), 1294 => to_unsigned(862, 10), 1295 => to_unsigned(407, 10), 1296 => to_unsigned(622, 10), 1297 => to_unsigned(564, 10), 1298 => to_unsigned(622, 10), 1299 => to_unsigned(544, 10), 1300 => to_unsigned(500, 10), 1301 => to_unsigned(698, 10), 1302 => to_unsigned(986, 10), 1303 => to_unsigned(583, 10), 1304 => to_unsigned(716, 10), 1305 => to_unsigned(48, 10), 1306 => to_unsigned(483, 10), 1307 => to_unsigned(359, 10), 1308 => to_unsigned(652, 10), 1309 => to_unsigned(485, 10), 1310 => to_unsigned(225, 10), 1311 => to_unsigned(337, 10), 1312 => to_unsigned(430, 10), 1313 => to_unsigned(520, 10), 1314 => to_unsigned(51, 10), 1315 => to_unsigned(197, 10), 1316 => to_unsigned(764, 10), 1317 => to_unsigned(797, 10), 1318 => to_unsigned(851, 10), 1319 => to_unsigned(336, 10), 1320 => to_unsigned(11, 10), 1321 => to_unsigned(740, 10), 1322 => to_unsigned(149, 10), 1323 => to_unsigned(618, 10), 1324 => to_unsigned(349, 10), 1325 => to_unsigned(648, 10), 1326 => to_unsigned(456, 10), 1327 => to_unsigned(949, 10), 1328 => to_unsigned(583, 10), 1329 => to_unsigned(329, 10), 1330 => to_unsigned(430, 10), 1331 => to_unsigned(113, 10), 1332 => to_unsigned(136, 10), 1333 => to_unsigned(293, 10), 1334 => to_unsigned(492, 10), 1335 => to_unsigned(849, 10), 1336 => to_unsigned(0, 10), 1337 => to_unsigned(477, 10), 1338 => to_unsigned(239, 10), 1339 => to_unsigned(121, 10), 1340 => to_unsigned(241, 10), 1341 => to_unsigned(427, 10), 1342 => to_unsigned(931, 10), 1343 => to_unsigned(1019, 10), 1344 => to_unsigned(857, 10), 1345 => to_unsigned(663, 10), 1346 => to_unsigned(752, 10), 1347 => to_unsigned(698, 10), 1348 => to_unsigned(159, 10), 1349 => to_unsigned(254, 10), 1350 => to_unsigned(838, 10), 1351 => to_unsigned(668, 10), 1352 => to_unsigned(125, 10), 1353 => to_unsigned(580, 10), 1354 => to_unsigned(180, 10), 1355 => to_unsigned(715, 10), 1356 => to_unsigned(209, 10), 1357 => to_unsigned(897, 10), 1358 => to_unsigned(583, 10), 1359 => to_unsigned(438, 10), 1360 => to_unsigned(680, 10), 1361 => to_unsigned(343, 10), 1362 => to_unsigned(790, 10), 1363 => to_unsigned(664, 10), 1364 => to_unsigned(995, 10), 1365 => to_unsigned(310, 10), 1366 => to_unsigned(231, 10), 1367 => to_unsigned(387, 10), 1368 => to_unsigned(498, 10), 1369 => to_unsigned(179, 10), 1370 => to_unsigned(997, 10), 1371 => to_unsigned(186, 10), 1372 => to_unsigned(951, 10), 1373 => to_unsigned(567, 10), 1374 => to_unsigned(224, 10), 1375 => to_unsigned(639, 10), 1376 => to_unsigned(352, 10), 1377 => to_unsigned(322, 10), 1378 => to_unsigned(796, 10), 1379 => to_unsigned(1004, 10), 1380 => to_unsigned(75, 10), 1381 => to_unsigned(509, 10), 1382 => to_unsigned(714, 10), 1383 => to_unsigned(175, 10), 1384 => to_unsigned(558, 10), 1385 => to_unsigned(55, 10), 1386 => to_unsigned(893, 10), 1387 => to_unsigned(851, 10), 1388 => to_unsigned(1016, 10), 1389 => to_unsigned(140, 10), 1390 => to_unsigned(471, 10), 1391 => to_unsigned(305, 10), 1392 => to_unsigned(297, 10), 1393 => to_unsigned(561, 10), 1394 => to_unsigned(323, 10), 1395 => to_unsigned(370, 10), 1396 => to_unsigned(99, 10), 1397 => to_unsigned(823, 10), 1398 => to_unsigned(55, 10), 1399 => to_unsigned(87, 10), 1400 => to_unsigned(505, 10), 1401 => to_unsigned(194, 10), 1402 => to_unsigned(319, 10), 1403 => to_unsigned(370, 10), 1404 => to_unsigned(213, 10), 1405 => to_unsigned(386, 10), 1406 => to_unsigned(539, 10), 1407 => to_unsigned(502, 10), 1408 => to_unsigned(61, 10), 1409 => to_unsigned(515, 10), 1410 => to_unsigned(197, 10), 1411 => to_unsigned(578, 10), 1412 => to_unsigned(846, 10), 1413 => to_unsigned(527, 10), 1414 => to_unsigned(416, 10), 1415 => to_unsigned(780, 10), 1416 => to_unsigned(944, 10), 1417 => to_unsigned(60, 10), 1418 => to_unsigned(954, 10), 1419 => to_unsigned(520, 10), 1420 => to_unsigned(967, 10), 1421 => to_unsigned(683, 10), 1422 => to_unsigned(894, 10), 1423 => to_unsigned(1011, 10), 1424 => to_unsigned(354, 10), 1425 => to_unsigned(205, 10), 1426 => to_unsigned(747, 10), 1427 => to_unsigned(824, 10), 1428 => to_unsigned(499, 10), 1429 => to_unsigned(588, 10), 1430 => to_unsigned(693, 10), 1431 => to_unsigned(805, 10), 1432 => to_unsigned(865, 10), 1433 => to_unsigned(111, 10), 1434 => to_unsigned(888, 10), 1435 => to_unsigned(488, 10), 1436 => to_unsigned(476, 10), 1437 => to_unsigned(588, 10), 1438 => to_unsigned(110, 10), 1439 => to_unsigned(497, 10), 1440 => to_unsigned(695, 10), 1441 => to_unsigned(33, 10), 1442 => to_unsigned(49, 10), 1443 => to_unsigned(995, 10), 1444 => to_unsigned(865, 10), 1445 => to_unsigned(860, 10), 1446 => to_unsigned(2, 10), 1447 => to_unsigned(926, 10), 1448 => to_unsigned(943, 10), 1449 => to_unsigned(132, 10), 1450 => to_unsigned(471, 10), 1451 => to_unsigned(910, 10), 1452 => to_unsigned(164, 10), 1453 => to_unsigned(836, 10), 1454 => to_unsigned(229, 10), 1455 => to_unsigned(760, 10), 1456 => to_unsigned(466, 10), 1457 => to_unsigned(83, 10), 1458 => to_unsigned(382, 10), 1459 => to_unsigned(563, 10), 1460 => to_unsigned(230, 10), 1461 => to_unsigned(593, 10), 1462 => to_unsigned(490, 10), 1463 => to_unsigned(755, 10), 1464 => to_unsigned(408, 10), 1465 => to_unsigned(310, 10), 1466 => to_unsigned(129, 10), 1467 => to_unsigned(102, 10), 1468 => to_unsigned(958, 10), 1469 => to_unsigned(821, 10), 1470 => to_unsigned(160, 10), 1471 => to_unsigned(962, 10), 1472 => to_unsigned(805, 10), 1473 => to_unsigned(329, 10), 1474 => to_unsigned(783, 10), 1475 => to_unsigned(5, 10), 1476 => to_unsigned(390, 10), 1477 => to_unsigned(28, 10), 1478 => to_unsigned(803, 10), 1479 => to_unsigned(292, 10), 1480 => to_unsigned(445, 10), 1481 => to_unsigned(712, 10), 1482 => to_unsigned(183, 10), 1483 => to_unsigned(306, 10), 1484 => to_unsigned(833, 10), 1485 => to_unsigned(326, 10), 1486 => to_unsigned(335, 10), 1487 => to_unsigned(447, 10), 1488 => to_unsigned(775, 10), 1489 => to_unsigned(693, 10), 1490 => to_unsigned(9, 10), 1491 => to_unsigned(752, 10), 1492 => to_unsigned(234, 10), 1493 => to_unsigned(592, 10), 1494 => to_unsigned(363, 10), 1495 => to_unsigned(978, 10), 1496 => to_unsigned(267, 10), 1497 => to_unsigned(597, 10), 1498 => to_unsigned(992, 10), 1499 => to_unsigned(245, 10), 1500 => to_unsigned(273, 10), 1501 => to_unsigned(265, 10), 1502 => to_unsigned(529, 10), 1503 => to_unsigned(763, 10), 1504 => to_unsigned(520, 10), 1505 => to_unsigned(228, 10), 1506 => to_unsigned(939, 10), 1507 => to_unsigned(283, 10), 1508 => to_unsigned(849, 10), 1509 => to_unsigned(553, 10), 1510 => to_unsigned(833, 10), 1511 => to_unsigned(365, 10), 1512 => to_unsigned(348, 10), 1513 => to_unsigned(726, 10), 1514 => to_unsigned(916, 10), 1515 => to_unsigned(355, 10), 1516 => to_unsigned(169, 10), 1517 => to_unsigned(401, 10), 1518 => to_unsigned(1003, 10), 1519 => to_unsigned(265, 10), 1520 => to_unsigned(671, 10), 1521 => to_unsigned(752, 10), 1522 => to_unsigned(32, 10), 1523 => to_unsigned(415, 10), 1524 => to_unsigned(139, 10), 1525 => to_unsigned(543, 10), 1526 => to_unsigned(758, 10), 1527 => to_unsigned(399, 10), 1528 => to_unsigned(952, 10), 1529 => to_unsigned(339, 10), 1530 => to_unsigned(669, 10), 1531 => to_unsigned(659, 10), 1532 => to_unsigned(793, 10), 1533 => to_unsigned(171, 10), 1534 => to_unsigned(597, 10), 1535 => to_unsigned(858, 10), 1536 => to_unsigned(320, 10), 1537 => to_unsigned(337, 10), 1538 => to_unsigned(128, 10), 1539 => to_unsigned(489, 10), 1540 => to_unsigned(121, 10), 1541 => to_unsigned(383, 10), 1542 => to_unsigned(969, 10), 1543 => to_unsigned(118, 10), 1544 => to_unsigned(169, 10), 1545 => to_unsigned(526, 10), 1546 => to_unsigned(171, 10), 1547 => to_unsigned(840, 10), 1548 => to_unsigned(228, 10), 1549 => to_unsigned(235, 10), 1550 => to_unsigned(1014, 10), 1551 => to_unsigned(612, 10), 1552 => to_unsigned(940, 10), 1553 => to_unsigned(971, 10), 1554 => to_unsigned(685, 10), 1555 => to_unsigned(723, 10), 1556 => to_unsigned(789, 10), 1557 => to_unsigned(140, 10), 1558 => to_unsigned(130, 10), 1559 => to_unsigned(1015, 10), 1560 => to_unsigned(258, 10), 1561 => to_unsigned(900, 10), 1562 => to_unsigned(201, 10), 1563 => to_unsigned(108, 10), 1564 => to_unsigned(44, 10), 1565 => to_unsigned(532, 10), 1566 => to_unsigned(212, 10), 1567 => to_unsigned(959, 10), 1568 => to_unsigned(60, 10), 1569 => to_unsigned(686, 10), 1570 => to_unsigned(213, 10), 1571 => to_unsigned(674, 10), 1572 => to_unsigned(695, 10), 1573 => to_unsigned(88, 10), 1574 => to_unsigned(1021, 10), 1575 => to_unsigned(678, 10), 1576 => to_unsigned(48, 10), 1577 => to_unsigned(928, 10), 1578 => to_unsigned(228, 10), 1579 => to_unsigned(422, 10), 1580 => to_unsigned(148, 10), 1581 => to_unsigned(232, 10), 1582 => to_unsigned(275, 10), 1583 => to_unsigned(14, 10), 1584 => to_unsigned(193, 10), 1585 => to_unsigned(1022, 10), 1586 => to_unsigned(410, 10), 1587 => to_unsigned(497, 10), 1588 => to_unsigned(777, 10), 1589 => to_unsigned(748, 10), 1590 => to_unsigned(1000, 10), 1591 => to_unsigned(871, 10), 1592 => to_unsigned(716, 10), 1593 => to_unsigned(372, 10), 1594 => to_unsigned(184, 10), 1595 => to_unsigned(796, 10), 1596 => to_unsigned(940, 10), 1597 => to_unsigned(132, 10), 1598 => to_unsigned(857, 10), 1599 => to_unsigned(800, 10), 1600 => to_unsigned(192, 10), 1601 => to_unsigned(359, 10), 1602 => to_unsigned(386, 10), 1603 => to_unsigned(875, 10), 1604 => to_unsigned(694, 10), 1605 => to_unsigned(49, 10), 1606 => to_unsigned(116, 10), 1607 => to_unsigned(764, 10), 1608 => to_unsigned(973, 10), 1609 => to_unsigned(162, 10), 1610 => to_unsigned(943, 10), 1611 => to_unsigned(358, 10), 1612 => to_unsigned(978, 10), 1613 => to_unsigned(932, 10), 1614 => to_unsigned(400, 10), 1615 => to_unsigned(952, 10), 1616 => to_unsigned(565, 10), 1617 => to_unsigned(931, 10), 1618 => to_unsigned(125, 10), 1619 => to_unsigned(48, 10), 1620 => to_unsigned(104, 10), 1621 => to_unsigned(937, 10), 1622 => to_unsigned(151, 10), 1623 => to_unsigned(481, 10), 1624 => to_unsigned(574, 10), 1625 => to_unsigned(706, 10), 1626 => to_unsigned(982, 10), 1627 => to_unsigned(862, 10), 1628 => to_unsigned(861, 10), 1629 => to_unsigned(776, 10), 1630 => to_unsigned(210, 10), 1631 => to_unsigned(636, 10), 1632 => to_unsigned(610, 10), 1633 => to_unsigned(871, 10), 1634 => to_unsigned(912, 10), 1635 => to_unsigned(824, 10), 1636 => to_unsigned(225, 10), 1637 => to_unsigned(22, 10), 1638 => to_unsigned(543, 10), 1639 => to_unsigned(947, 10), 1640 => to_unsigned(859, 10), 1641 => to_unsigned(250, 10), 1642 => to_unsigned(516, 10), 1643 => to_unsigned(66, 10), 1644 => to_unsigned(857, 10), 1645 => to_unsigned(794, 10), 1646 => to_unsigned(883, 10), 1647 => to_unsigned(511, 10), 1648 => to_unsigned(597, 10), 1649 => to_unsigned(739, 10), 1650 => to_unsigned(493, 10), 1651 => to_unsigned(873, 10), 1652 => to_unsigned(152, 10), 1653 => to_unsigned(581, 10), 1654 => to_unsigned(768, 10), 1655 => to_unsigned(826, 10), 1656 => to_unsigned(867, 10), 1657 => to_unsigned(317, 10), 1658 => to_unsigned(770, 10), 1659 => to_unsigned(660, 10), 1660 => to_unsigned(472, 10), 1661 => to_unsigned(781, 10), 1662 => to_unsigned(424, 10), 1663 => to_unsigned(714, 10), 1664 => to_unsigned(887, 10), 1665 => to_unsigned(229, 10), 1666 => to_unsigned(734, 10), 1667 => to_unsigned(723, 10), 1668 => to_unsigned(842, 10), 1669 => to_unsigned(403, 10), 1670 => to_unsigned(310, 10), 1671 => to_unsigned(699, 10), 1672 => to_unsigned(703, 10), 1673 => to_unsigned(539, 10), 1674 => to_unsigned(34, 10), 1675 => to_unsigned(161, 10), 1676 => to_unsigned(652, 10), 1677 => to_unsigned(218, 10), 1678 => to_unsigned(803, 10), 1679 => to_unsigned(375, 10), 1680 => to_unsigned(247, 10), 1681 => to_unsigned(333, 10), 1682 => to_unsigned(290, 10), 1683 => to_unsigned(748, 10), 1684 => to_unsigned(122, 10), 1685 => to_unsigned(304, 10), 1686 => to_unsigned(609, 10), 1687 => to_unsigned(456, 10), 1688 => to_unsigned(184, 10), 1689 => to_unsigned(666, 10), 1690 => to_unsigned(796, 10), 1691 => to_unsigned(412, 10), 1692 => to_unsigned(947, 10), 1693 => to_unsigned(720, 10), 1694 => to_unsigned(329, 10), 1695 => to_unsigned(680, 10), 1696 => to_unsigned(872, 10), 1697 => to_unsigned(324, 10), 1698 => to_unsigned(261, 10), 1699 => to_unsigned(453, 10), 1700 => to_unsigned(787, 10), 1701 => to_unsigned(356, 10), 1702 => to_unsigned(194, 10), 1703 => to_unsigned(226, 10), 1704 => to_unsigned(243, 10), 1705 => to_unsigned(373, 10), 1706 => to_unsigned(160, 10), 1707 => to_unsigned(467, 10), 1708 => to_unsigned(182, 10), 1709 => to_unsigned(293, 10), 1710 => to_unsigned(432, 10), 1711 => to_unsigned(708, 10), 1712 => to_unsigned(759, 10), 1713 => to_unsigned(4, 10), 1714 => to_unsigned(946, 10), 1715 => to_unsigned(760, 10), 1716 => to_unsigned(969, 10), 1717 => to_unsigned(754, 10), 1718 => to_unsigned(1013, 10), 1719 => to_unsigned(71, 10), 1720 => to_unsigned(128, 10), 1721 => to_unsigned(450, 10), 1722 => to_unsigned(1021, 10), 1723 => to_unsigned(259, 10), 1724 => to_unsigned(584, 10), 1725 => to_unsigned(618, 10), 1726 => to_unsigned(6, 10), 1727 => to_unsigned(739, 10), 1728 => to_unsigned(30, 10), 1729 => to_unsigned(212, 10), 1730 => to_unsigned(759, 10), 1731 => to_unsigned(170, 10), 1732 => to_unsigned(306, 10), 1733 => to_unsigned(602, 10), 1734 => to_unsigned(170, 10), 1735 => to_unsigned(1002, 10), 1736 => to_unsigned(37, 10), 1737 => to_unsigned(294, 10), 1738 => to_unsigned(996, 10), 1739 => to_unsigned(975, 10), 1740 => to_unsigned(242, 10), 1741 => to_unsigned(258, 10), 1742 => to_unsigned(57, 10), 1743 => to_unsigned(661, 10), 1744 => to_unsigned(428, 10), 1745 => to_unsigned(176, 10), 1746 => to_unsigned(908, 10), 1747 => to_unsigned(143, 10), 1748 => to_unsigned(139, 10), 1749 => to_unsigned(405, 10), 1750 => to_unsigned(385, 10), 1751 => to_unsigned(77, 10), 1752 => to_unsigned(529, 10), 1753 => to_unsigned(121, 10), 1754 => to_unsigned(165, 10), 1755 => to_unsigned(933, 10), 1756 => to_unsigned(729, 10), 1757 => to_unsigned(884, 10), 1758 => to_unsigned(377, 10), 1759 => to_unsigned(972, 10), 1760 => to_unsigned(909, 10), 1761 => to_unsigned(951, 10), 1762 => to_unsigned(737, 10), 1763 => to_unsigned(899, 10), 1764 => to_unsigned(304, 10), 1765 => to_unsigned(176, 10), 1766 => to_unsigned(804, 10), 1767 => to_unsigned(1023, 10), 1768 => to_unsigned(421, 10), 1769 => to_unsigned(999, 10), 1770 => to_unsigned(418, 10), 1771 => to_unsigned(421, 10), 1772 => to_unsigned(394, 10), 1773 => to_unsigned(546, 10), 1774 => to_unsigned(861, 10), 1775 => to_unsigned(737, 10), 1776 => to_unsigned(796, 10), 1777 => to_unsigned(46, 10), 1778 => to_unsigned(1013, 10), 1779 => to_unsigned(29, 10), 1780 => to_unsigned(438, 10), 1781 => to_unsigned(1009, 10), 1782 => to_unsigned(734, 10), 1783 => to_unsigned(38, 10), 1784 => to_unsigned(704, 10), 1785 => to_unsigned(349, 10), 1786 => to_unsigned(576, 10), 1787 => to_unsigned(207, 10), 1788 => to_unsigned(448, 10), 1789 => to_unsigned(486, 10), 1790 => to_unsigned(399, 10), 1791 => to_unsigned(6, 10), 1792 => to_unsigned(518, 10), 1793 => to_unsigned(648, 10), 1794 => to_unsigned(672, 10), 1795 => to_unsigned(558, 10), 1796 => to_unsigned(294, 10), 1797 => to_unsigned(366, 10), 1798 => to_unsigned(235, 10), 1799 => to_unsigned(162, 10), 1800 => to_unsigned(501, 10), 1801 => to_unsigned(896, 10), 1802 => to_unsigned(688, 10), 1803 => to_unsigned(867, 10), 1804 => to_unsigned(916, 10), 1805 => to_unsigned(973, 10), 1806 => to_unsigned(435, 10), 1807 => to_unsigned(183, 10), 1808 => to_unsigned(727, 10), 1809 => to_unsigned(485, 10), 1810 => to_unsigned(12, 10), 1811 => to_unsigned(538, 10), 1812 => to_unsigned(670, 10), 1813 => to_unsigned(669, 10), 1814 => to_unsigned(633, 10), 1815 => to_unsigned(559, 10), 1816 => to_unsigned(215, 10), 1817 => to_unsigned(719, 10), 1818 => to_unsigned(301, 10), 1819 => to_unsigned(775, 10), 1820 => to_unsigned(757, 10), 1821 => to_unsigned(568, 10), 1822 => to_unsigned(916, 10), 1823 => to_unsigned(235, 10), 1824 => to_unsigned(248, 10), 1825 => to_unsigned(771, 10), 1826 => to_unsigned(479, 10), 1827 => to_unsigned(375, 10), 1828 => to_unsigned(314, 10), 1829 => to_unsigned(768, 10), 1830 => to_unsigned(420, 10), 1831 => to_unsigned(764, 10), 1832 => to_unsigned(263, 10), 1833 => to_unsigned(637, 10), 1834 => to_unsigned(283, 10), 1835 => to_unsigned(530, 10), 1836 => to_unsigned(219, 10), 1837 => to_unsigned(942, 10), 1838 => to_unsigned(802, 10), 1839 => to_unsigned(338, 10), 1840 => to_unsigned(239, 10), 1841 => to_unsigned(370, 10), 1842 => to_unsigned(512, 10), 1843 => to_unsigned(605, 10), 1844 => to_unsigned(1017, 10), 1845 => to_unsigned(374, 10), 1846 => to_unsigned(477, 10), 1847 => to_unsigned(1015, 10), 1848 => to_unsigned(796, 10), 1849 => to_unsigned(143, 10), 1850 => to_unsigned(1020, 10), 1851 => to_unsigned(939, 10), 1852 => to_unsigned(194, 10), 1853 => to_unsigned(49, 10), 1854 => to_unsigned(839, 10), 1855 => to_unsigned(774, 10), 1856 => to_unsigned(196, 10), 1857 => to_unsigned(624, 10), 1858 => to_unsigned(621, 10), 1859 => to_unsigned(665, 10), 1860 => to_unsigned(942, 10), 1861 => to_unsigned(464, 10), 1862 => to_unsigned(764, 10), 1863 => to_unsigned(75, 10), 1864 => to_unsigned(489, 10), 1865 => to_unsigned(836, 10), 1866 => to_unsigned(286, 10), 1867 => to_unsigned(762, 10), 1868 => to_unsigned(408, 10), 1869 => to_unsigned(372, 10), 1870 => to_unsigned(774, 10), 1871 => to_unsigned(182, 10), 1872 => to_unsigned(311, 10), 1873 => to_unsigned(626, 10), 1874 => to_unsigned(480, 10), 1875 => to_unsigned(983, 10), 1876 => to_unsigned(83, 10), 1877 => to_unsigned(357, 10), 1878 => to_unsigned(166, 10), 1879 => to_unsigned(550, 10), 1880 => to_unsigned(826, 10), 1881 => to_unsigned(836, 10), 1882 => to_unsigned(204, 10), 1883 => to_unsigned(465, 10), 1884 => to_unsigned(702, 10), 1885 => to_unsigned(648, 10), 1886 => to_unsigned(545, 10), 1887 => to_unsigned(201, 10), 1888 => to_unsigned(551, 10), 1889 => to_unsigned(36, 10), 1890 => to_unsigned(978, 10), 1891 => to_unsigned(512, 10), 1892 => to_unsigned(632, 10), 1893 => to_unsigned(528, 10), 1894 => to_unsigned(619, 10), 1895 => to_unsigned(327, 10), 1896 => to_unsigned(818, 10), 1897 => to_unsigned(439, 10), 1898 => to_unsigned(305, 10), 1899 => to_unsigned(434, 10), 1900 => to_unsigned(743, 10), 1901 => to_unsigned(210, 10), 1902 => to_unsigned(388, 10), 1903 => to_unsigned(153, 10), 1904 => to_unsigned(778, 10), 1905 => to_unsigned(96, 10), 1906 => to_unsigned(45, 10), 1907 => to_unsigned(341, 10), 1908 => to_unsigned(354, 10), 1909 => to_unsigned(436, 10), 1910 => to_unsigned(270, 10), 1911 => to_unsigned(286, 10), 1912 => to_unsigned(74, 10), 1913 => to_unsigned(327, 10), 1914 => to_unsigned(80, 10), 1915 => to_unsigned(1004, 10), 1916 => to_unsigned(27, 10), 1917 => to_unsigned(876, 10), 1918 => to_unsigned(52, 10), 1919 => to_unsigned(416, 10), 1920 => to_unsigned(423, 10), 1921 => to_unsigned(631, 10), 1922 => to_unsigned(440, 10), 1923 => to_unsigned(1021, 10), 1924 => to_unsigned(535, 10), 1925 => to_unsigned(242, 10), 1926 => to_unsigned(829, 10), 1927 => to_unsigned(838, 10), 1928 => to_unsigned(140, 10), 1929 => to_unsigned(627, 10), 1930 => to_unsigned(388, 10), 1931 => to_unsigned(914, 10), 1932 => to_unsigned(590, 10), 1933 => to_unsigned(788, 10), 1934 => to_unsigned(869, 10), 1935 => to_unsigned(184, 10), 1936 => to_unsigned(803, 10), 1937 => to_unsigned(326, 10), 1938 => to_unsigned(236, 10), 1939 => to_unsigned(29, 10), 1940 => to_unsigned(123, 10), 1941 => to_unsigned(138, 10), 1942 => to_unsigned(218, 10), 1943 => to_unsigned(386, 10), 1944 => to_unsigned(470, 10), 1945 => to_unsigned(613, 10), 1946 => to_unsigned(401, 10), 1947 => to_unsigned(46, 10), 1948 => to_unsigned(737, 10), 1949 => to_unsigned(284, 10), 1950 => to_unsigned(178, 10), 1951 => to_unsigned(962, 10), 1952 => to_unsigned(41, 10), 1953 => to_unsigned(456, 10), 1954 => to_unsigned(402, 10), 1955 => to_unsigned(396, 10), 1956 => to_unsigned(209, 10), 1957 => to_unsigned(493, 10), 1958 => to_unsigned(693, 10), 1959 => to_unsigned(284, 10), 1960 => to_unsigned(360, 10), 1961 => to_unsigned(249, 10), 1962 => to_unsigned(274, 10), 1963 => to_unsigned(591, 10), 1964 => to_unsigned(828, 10), 1965 => to_unsigned(384, 10), 1966 => to_unsigned(630, 10), 1967 => to_unsigned(940, 10), 1968 => to_unsigned(644, 10), 1969 => to_unsigned(461, 10), 1970 => to_unsigned(430, 10), 1971 => to_unsigned(749, 10), 1972 => to_unsigned(203, 10), 1973 => to_unsigned(667, 10), 1974 => to_unsigned(747, 10), 1975 => to_unsigned(955, 10), 1976 => to_unsigned(903, 10), 1977 => to_unsigned(693, 10), 1978 => to_unsigned(664, 10), 1979 => to_unsigned(11, 10), 1980 => to_unsigned(794, 10), 1981 => to_unsigned(99, 10), 1982 => to_unsigned(959, 10), 1983 => to_unsigned(655, 10), 1984 => to_unsigned(204, 10), 1985 => to_unsigned(718, 10), 1986 => to_unsigned(710, 10), 1987 => to_unsigned(274, 10), 1988 => to_unsigned(371, 10), 1989 => to_unsigned(508, 10), 1990 => to_unsigned(616, 10), 1991 => to_unsigned(15, 10), 1992 => to_unsigned(942, 10), 1993 => to_unsigned(980, 10), 1994 => to_unsigned(849, 10), 1995 => to_unsigned(968, 10), 1996 => to_unsigned(860, 10), 1997 => to_unsigned(910, 10), 1998 => to_unsigned(161, 10), 1999 => to_unsigned(309, 10), 2000 => to_unsigned(95, 10), 2001 => to_unsigned(651, 10), 2002 => to_unsigned(309, 10), 2003 => to_unsigned(9, 10), 2004 => to_unsigned(108, 10), 2005 => to_unsigned(288, 10), 2006 => to_unsigned(751, 10), 2007 => to_unsigned(104, 10), 2008 => to_unsigned(341, 10), 2009 => to_unsigned(615, 10), 2010 => to_unsigned(650, 10), 2011 => to_unsigned(225, 10), 2012 => to_unsigned(393, 10), 2013 => to_unsigned(540, 10), 2014 => to_unsigned(130, 10), 2015 => to_unsigned(890, 10), 2016 => to_unsigned(653, 10), 2017 => to_unsigned(250, 10), 2018 => to_unsigned(234, 10), 2019 => to_unsigned(779, 10), 2020 => to_unsigned(846, 10), 2021 => to_unsigned(109, 10), 2022 => to_unsigned(985, 10), 2023 => to_unsigned(0, 10), 2024 => to_unsigned(984, 10), 2025 => to_unsigned(747, 10), 2026 => to_unsigned(455, 10), 2027 => to_unsigned(18, 10), 2028 => to_unsigned(691, 10), 2029 => to_unsigned(897, 10), 2030 => to_unsigned(703, 10), 2031 => to_unsigned(4, 10), 2032 => to_unsigned(806, 10), 2033 => to_unsigned(677, 10), 2034 => to_unsigned(633, 10), 2035 => to_unsigned(380, 10), 2036 => to_unsigned(338, 10), 2037 => to_unsigned(229, 10), 2038 => to_unsigned(184, 10), 2039 => to_unsigned(265, 10), 2040 => to_unsigned(721, 10), 2041 => to_unsigned(104, 10), 2042 => to_unsigned(102, 10), 2043 => to_unsigned(852, 10), 2044 => to_unsigned(781, 10), 2045 => to_unsigned(559, 10), 2046 => to_unsigned(282, 10), 2047 => to_unsigned(825, 10)),
            5 => (0 => to_unsigned(707, 10), 1 => to_unsigned(273, 10), 2 => to_unsigned(800, 10), 3 => to_unsigned(782, 10), 4 => to_unsigned(971, 10), 5 => to_unsigned(359, 10), 6 => to_unsigned(169, 10), 7 => to_unsigned(410, 10), 8 => to_unsigned(568, 10), 9 => to_unsigned(851, 10), 10 => to_unsigned(3, 10), 11 => to_unsigned(658, 10), 12 => to_unsigned(46, 10), 13 => to_unsigned(32, 10), 14 => to_unsigned(369, 10), 15 => to_unsigned(440, 10), 16 => to_unsigned(786, 10), 17 => to_unsigned(1012, 10), 18 => to_unsigned(450, 10), 19 => to_unsigned(312, 10), 20 => to_unsigned(991, 10), 21 => to_unsigned(1020, 10), 22 => to_unsigned(68, 10), 23 => to_unsigned(324, 10), 24 => to_unsigned(774, 10), 25 => to_unsigned(499, 10), 26 => to_unsigned(454, 10), 27 => to_unsigned(129, 10), 28 => to_unsigned(589, 10), 29 => to_unsigned(514, 10), 30 => to_unsigned(437, 10), 31 => to_unsigned(848, 10), 32 => to_unsigned(591, 10), 33 => to_unsigned(14, 10), 34 => to_unsigned(114, 10), 35 => to_unsigned(263, 10), 36 => to_unsigned(459, 10), 37 => to_unsigned(594, 10), 38 => to_unsigned(419, 10), 39 => to_unsigned(631, 10), 40 => to_unsigned(131, 10), 41 => to_unsigned(896, 10), 42 => to_unsigned(173, 10), 43 => to_unsigned(692, 10), 44 => to_unsigned(147, 10), 45 => to_unsigned(743, 10), 46 => to_unsigned(757, 10), 47 => to_unsigned(722, 10), 48 => to_unsigned(368, 10), 49 => to_unsigned(266, 10), 50 => to_unsigned(237, 10), 51 => to_unsigned(45, 10), 52 => to_unsigned(225, 10), 53 => to_unsigned(599, 10), 54 => to_unsigned(24, 10), 55 => to_unsigned(982, 10), 56 => to_unsigned(589, 10), 57 => to_unsigned(479, 10), 58 => to_unsigned(511, 10), 59 => to_unsigned(523, 10), 60 => to_unsigned(133, 10), 61 => to_unsigned(309, 10), 62 => to_unsigned(882, 10), 63 => to_unsigned(546, 10), 64 => to_unsigned(120, 10), 65 => to_unsigned(843, 10), 66 => to_unsigned(929, 10), 67 => to_unsigned(390, 10), 68 => to_unsigned(408, 10), 69 => to_unsigned(64, 10), 70 => to_unsigned(517, 10), 71 => to_unsigned(431, 10), 72 => to_unsigned(866, 10), 73 => to_unsigned(31, 10), 74 => to_unsigned(347, 10), 75 => to_unsigned(782, 10), 76 => to_unsigned(648, 10), 77 => to_unsigned(254, 10), 78 => to_unsigned(659, 10), 79 => to_unsigned(756, 10), 80 => to_unsigned(343, 10), 81 => to_unsigned(999, 10), 82 => to_unsigned(886, 10), 83 => to_unsigned(772, 10), 84 => to_unsigned(664, 10), 85 => to_unsigned(396, 10), 86 => to_unsigned(841, 10), 87 => to_unsigned(77, 10), 88 => to_unsigned(147, 10), 89 => to_unsigned(1023, 10), 90 => to_unsigned(747, 10), 91 => to_unsigned(37, 10), 92 => to_unsigned(343, 10), 93 => to_unsigned(141, 10), 94 => to_unsigned(146, 10), 95 => to_unsigned(575, 10), 96 => to_unsigned(492, 10), 97 => to_unsigned(205, 10), 98 => to_unsigned(369, 10), 99 => to_unsigned(314, 10), 100 => to_unsigned(910, 10), 101 => to_unsigned(938, 10), 102 => to_unsigned(15, 10), 103 => to_unsigned(385, 10), 104 => to_unsigned(438, 10), 105 => to_unsigned(205, 10), 106 => to_unsigned(47, 10), 107 => to_unsigned(435, 10), 108 => to_unsigned(547, 10), 109 => to_unsigned(696, 10), 110 => to_unsigned(193, 10), 111 => to_unsigned(910, 10), 112 => to_unsigned(135, 10), 113 => to_unsigned(524, 10), 114 => to_unsigned(286, 10), 115 => to_unsigned(500, 10), 116 => to_unsigned(287, 10), 117 => to_unsigned(509, 10), 118 => to_unsigned(16, 10), 119 => to_unsigned(197, 10), 120 => to_unsigned(491, 10), 121 => to_unsigned(425, 10), 122 => to_unsigned(389, 10), 123 => to_unsigned(792, 10), 124 => to_unsigned(800, 10), 125 => to_unsigned(651, 10), 126 => to_unsigned(52, 10), 127 => to_unsigned(892, 10), 128 => to_unsigned(165, 10), 129 => to_unsigned(359, 10), 130 => to_unsigned(497, 10), 131 => to_unsigned(860, 10), 132 => to_unsigned(930, 10), 133 => to_unsigned(157, 10), 134 => to_unsigned(885, 10), 135 => to_unsigned(199, 10), 136 => to_unsigned(60, 10), 137 => to_unsigned(479, 10), 138 => to_unsigned(419, 10), 139 => to_unsigned(428, 10), 140 => to_unsigned(70, 10), 141 => to_unsigned(642, 10), 142 => to_unsigned(524, 10), 143 => to_unsigned(764, 10), 144 => to_unsigned(915, 10), 145 => to_unsigned(884, 10), 146 => to_unsigned(992, 10), 147 => to_unsigned(869, 10), 148 => to_unsigned(104, 10), 149 => to_unsigned(339, 10), 150 => to_unsigned(840, 10), 151 => to_unsigned(951, 10), 152 => to_unsigned(16, 10), 153 => to_unsigned(613, 10), 154 => to_unsigned(98, 10), 155 => to_unsigned(593, 10), 156 => to_unsigned(57, 10), 157 => to_unsigned(125, 10), 158 => to_unsigned(621, 10), 159 => to_unsigned(866, 10), 160 => to_unsigned(233, 10), 161 => to_unsigned(584, 10), 162 => to_unsigned(165, 10), 163 => to_unsigned(735, 10), 164 => to_unsigned(307, 10), 165 => to_unsigned(323, 10), 166 => to_unsigned(817, 10), 167 => to_unsigned(408, 10), 168 => to_unsigned(457, 10), 169 => to_unsigned(733, 10), 170 => to_unsigned(262, 10), 171 => to_unsigned(59, 10), 172 => to_unsigned(1005, 10), 173 => to_unsigned(419, 10), 174 => to_unsigned(781, 10), 175 => to_unsigned(273, 10), 176 => to_unsigned(926, 10), 177 => to_unsigned(210, 10), 178 => to_unsigned(593, 10), 179 => to_unsigned(920, 10), 180 => to_unsigned(683, 10), 181 => to_unsigned(788, 10), 182 => to_unsigned(591, 10), 183 => to_unsigned(612, 10), 184 => to_unsigned(978, 10), 185 => to_unsigned(261, 10), 186 => to_unsigned(85, 10), 187 => to_unsigned(767, 10), 188 => to_unsigned(497, 10), 189 => to_unsigned(437, 10), 190 => to_unsigned(479, 10), 191 => to_unsigned(721, 10), 192 => to_unsigned(642, 10), 193 => to_unsigned(380, 10), 194 => to_unsigned(169, 10), 195 => to_unsigned(950, 10), 196 => to_unsigned(281, 10), 197 => to_unsigned(275, 10), 198 => to_unsigned(205, 10), 199 => to_unsigned(220, 10), 200 => to_unsigned(721, 10), 201 => to_unsigned(1009, 10), 202 => to_unsigned(725, 10), 203 => to_unsigned(837, 10), 204 => to_unsigned(400, 10), 205 => to_unsigned(697, 10), 206 => to_unsigned(967, 10), 207 => to_unsigned(81, 10), 208 => to_unsigned(227, 10), 209 => to_unsigned(303, 10), 210 => to_unsigned(730, 10), 211 => to_unsigned(589, 10), 212 => to_unsigned(405, 10), 213 => to_unsigned(390, 10), 214 => to_unsigned(6, 10), 215 => to_unsigned(314, 10), 216 => to_unsigned(404, 10), 217 => to_unsigned(962, 10), 218 => to_unsigned(195, 10), 219 => to_unsigned(881, 10), 220 => to_unsigned(832, 10), 221 => to_unsigned(1021, 10), 222 => to_unsigned(930, 10), 223 => to_unsigned(868, 10), 224 => to_unsigned(421, 10), 225 => to_unsigned(943, 10), 226 => to_unsigned(393, 10), 227 => to_unsigned(188, 10), 228 => to_unsigned(654, 10), 229 => to_unsigned(957, 10), 230 => to_unsigned(60, 10), 231 => to_unsigned(782, 10), 232 => to_unsigned(120, 10), 233 => to_unsigned(620, 10), 234 => to_unsigned(825, 10), 235 => to_unsigned(736, 10), 236 => to_unsigned(28, 10), 237 => to_unsigned(671, 10), 238 => to_unsigned(605, 10), 239 => to_unsigned(318, 10), 240 => to_unsigned(239, 10), 241 => to_unsigned(480, 10), 242 => to_unsigned(626, 10), 243 => to_unsigned(994, 10), 244 => to_unsigned(849, 10), 245 => to_unsigned(272, 10), 246 => to_unsigned(413, 10), 247 => to_unsigned(95, 10), 248 => to_unsigned(856, 10), 249 => to_unsigned(75, 10), 250 => to_unsigned(884, 10), 251 => to_unsigned(172, 10), 252 => to_unsigned(309, 10), 253 => to_unsigned(790, 10), 254 => to_unsigned(645, 10), 255 => to_unsigned(437, 10), 256 => to_unsigned(9, 10), 257 => to_unsigned(616, 10), 258 => to_unsigned(212, 10), 259 => to_unsigned(889, 10), 260 => to_unsigned(215, 10), 261 => to_unsigned(959, 10), 262 => to_unsigned(53, 10), 263 => to_unsigned(120, 10), 264 => to_unsigned(835, 10), 265 => to_unsigned(423, 10), 266 => to_unsigned(446, 10), 267 => to_unsigned(405, 10), 268 => to_unsigned(755, 10), 269 => to_unsigned(58, 10), 270 => to_unsigned(504, 10), 271 => to_unsigned(267, 10), 272 => to_unsigned(804, 10), 273 => to_unsigned(138, 10), 274 => to_unsigned(440, 10), 275 => to_unsigned(710, 10), 276 => to_unsigned(635, 10), 277 => to_unsigned(500, 10), 278 => to_unsigned(746, 10), 279 => to_unsigned(822, 10), 280 => to_unsigned(697, 10), 281 => to_unsigned(421, 10), 282 => to_unsigned(967, 10), 283 => to_unsigned(648, 10), 284 => to_unsigned(608, 10), 285 => to_unsigned(913, 10), 286 => to_unsigned(44, 10), 287 => to_unsigned(936, 10), 288 => to_unsigned(121, 10), 289 => to_unsigned(60, 10), 290 => to_unsigned(346, 10), 291 => to_unsigned(992, 10), 292 => to_unsigned(308, 10), 293 => to_unsigned(134, 10), 294 => to_unsigned(405, 10), 295 => to_unsigned(889, 10), 296 => to_unsigned(496, 10), 297 => to_unsigned(713, 10), 298 => to_unsigned(99, 10), 299 => to_unsigned(138, 10), 300 => to_unsigned(743, 10), 301 => to_unsigned(935, 10), 302 => to_unsigned(489, 10), 303 => to_unsigned(563, 10), 304 => to_unsigned(178, 10), 305 => to_unsigned(478, 10), 306 => to_unsigned(598, 10), 307 => to_unsigned(212, 10), 308 => to_unsigned(909, 10), 309 => to_unsigned(648, 10), 310 => to_unsigned(426, 10), 311 => to_unsigned(972, 10), 312 => to_unsigned(218, 10), 313 => to_unsigned(25, 10), 314 => to_unsigned(857, 10), 315 => to_unsigned(756, 10), 316 => to_unsigned(54, 10), 317 => to_unsigned(472, 10), 318 => to_unsigned(51, 10), 319 => to_unsigned(218, 10), 320 => to_unsigned(909, 10), 321 => to_unsigned(295, 10), 322 => to_unsigned(370, 10), 323 => to_unsigned(570, 10), 324 => to_unsigned(975, 10), 325 => to_unsigned(801, 10), 326 => to_unsigned(773, 10), 327 => to_unsigned(882, 10), 328 => to_unsigned(921, 10), 329 => to_unsigned(806, 10), 330 => to_unsigned(1014, 10), 331 => to_unsigned(729, 10), 332 => to_unsigned(695, 10), 333 => to_unsigned(321, 10), 334 => to_unsigned(337, 10), 335 => to_unsigned(908, 10), 336 => to_unsigned(555, 10), 337 => to_unsigned(733, 10), 338 => to_unsigned(288, 10), 339 => to_unsigned(851, 10), 340 => to_unsigned(405, 10), 341 => to_unsigned(268, 10), 342 => to_unsigned(749, 10), 343 => to_unsigned(320, 10), 344 => to_unsigned(401, 10), 345 => to_unsigned(517, 10), 346 => to_unsigned(649, 10), 347 => to_unsigned(126, 10), 348 => to_unsigned(100, 10), 349 => to_unsigned(394, 10), 350 => to_unsigned(578, 10), 351 => to_unsigned(72, 10), 352 => to_unsigned(95, 10), 353 => to_unsigned(23, 10), 354 => to_unsigned(194, 10), 355 => to_unsigned(253, 10), 356 => to_unsigned(642, 10), 357 => to_unsigned(490, 10), 358 => to_unsigned(217, 10), 359 => to_unsigned(813, 10), 360 => to_unsigned(413, 10), 361 => to_unsigned(935, 10), 362 => to_unsigned(573, 10), 363 => to_unsigned(318, 10), 364 => to_unsigned(80, 10), 365 => to_unsigned(852, 10), 366 => to_unsigned(151, 10), 367 => to_unsigned(489, 10), 368 => to_unsigned(293, 10), 369 => to_unsigned(993, 10), 370 => to_unsigned(996, 10), 371 => to_unsigned(477, 10), 372 => to_unsigned(82, 10), 373 => to_unsigned(219, 10), 374 => to_unsigned(608, 10), 375 => to_unsigned(371, 10), 376 => to_unsigned(82, 10), 377 => to_unsigned(656, 10), 378 => to_unsigned(0, 10), 379 => to_unsigned(907, 10), 380 => to_unsigned(287, 10), 381 => to_unsigned(192, 10), 382 => to_unsigned(682, 10), 383 => to_unsigned(263, 10), 384 => to_unsigned(468, 10), 385 => to_unsigned(242, 10), 386 => to_unsigned(514, 10), 387 => to_unsigned(637, 10), 388 => to_unsigned(237, 10), 389 => to_unsigned(51, 10), 390 => to_unsigned(695, 10), 391 => to_unsigned(154, 10), 392 => to_unsigned(807, 10), 393 => to_unsigned(238, 10), 394 => to_unsigned(360, 10), 395 => to_unsigned(1022, 10), 396 => to_unsigned(925, 10), 397 => to_unsigned(466, 10), 398 => to_unsigned(169, 10), 399 => to_unsigned(537, 10), 400 => to_unsigned(940, 10), 401 => to_unsigned(770, 10), 402 => to_unsigned(334, 10), 403 => to_unsigned(426, 10), 404 => to_unsigned(898, 10), 405 => to_unsigned(98, 10), 406 => to_unsigned(915, 10), 407 => to_unsigned(502, 10), 408 => to_unsigned(811, 10), 409 => to_unsigned(777, 10), 410 => to_unsigned(844, 10), 411 => to_unsigned(106, 10), 412 => to_unsigned(129, 10), 413 => to_unsigned(410, 10), 414 => to_unsigned(192, 10), 415 => to_unsigned(153, 10), 416 => to_unsigned(381, 10), 417 => to_unsigned(708, 10), 418 => to_unsigned(849, 10), 419 => to_unsigned(40, 10), 420 => to_unsigned(518, 10), 421 => to_unsigned(263, 10), 422 => to_unsigned(441, 10), 423 => to_unsigned(556, 10), 424 => to_unsigned(433, 10), 425 => to_unsigned(586, 10), 426 => to_unsigned(651, 10), 427 => to_unsigned(743, 10), 428 => to_unsigned(337, 10), 429 => to_unsigned(919, 10), 430 => to_unsigned(30, 10), 431 => to_unsigned(41, 10), 432 => to_unsigned(829, 10), 433 => to_unsigned(136, 10), 434 => to_unsigned(338, 10), 435 => to_unsigned(217, 10), 436 => to_unsigned(925, 10), 437 => to_unsigned(121, 10), 438 => to_unsigned(801, 10), 439 => to_unsigned(195, 10), 440 => to_unsigned(792, 10), 441 => to_unsigned(640, 10), 442 => to_unsigned(941, 10), 443 => to_unsigned(329, 10), 444 => to_unsigned(712, 10), 445 => to_unsigned(29, 10), 446 => to_unsigned(270, 10), 447 => to_unsigned(547, 10), 448 => to_unsigned(598, 10), 449 => to_unsigned(130, 10), 450 => to_unsigned(275, 10), 451 => to_unsigned(539, 10), 452 => to_unsigned(666, 10), 453 => to_unsigned(405, 10), 454 => to_unsigned(447, 10), 455 => to_unsigned(306, 10), 456 => to_unsigned(8, 10), 457 => to_unsigned(190, 10), 458 => to_unsigned(349, 10), 459 => to_unsigned(743, 10), 460 => to_unsigned(849, 10), 461 => to_unsigned(74, 10), 462 => to_unsigned(552, 10), 463 => to_unsigned(909, 10), 464 => to_unsigned(145, 10), 465 => to_unsigned(633, 10), 466 => to_unsigned(79, 10), 467 => to_unsigned(567, 10), 468 => to_unsigned(212, 10), 469 => to_unsigned(226, 10), 470 => to_unsigned(732, 10), 471 => to_unsigned(419, 10), 472 => to_unsigned(266, 10), 473 => to_unsigned(894, 10), 474 => to_unsigned(199, 10), 475 => to_unsigned(47, 10), 476 => to_unsigned(589, 10), 477 => to_unsigned(633, 10), 478 => to_unsigned(568, 10), 479 => to_unsigned(117, 10), 480 => to_unsigned(770, 10), 481 => to_unsigned(199, 10), 482 => to_unsigned(761, 10), 483 => to_unsigned(983, 10), 484 => to_unsigned(695, 10), 485 => to_unsigned(665, 10), 486 => to_unsigned(285, 10), 487 => to_unsigned(222, 10), 488 => to_unsigned(607, 10), 489 => to_unsigned(219, 10), 490 => to_unsigned(225, 10), 491 => to_unsigned(405, 10), 492 => to_unsigned(321, 10), 493 => to_unsigned(257, 10), 494 => to_unsigned(377, 10), 495 => to_unsigned(139, 10), 496 => to_unsigned(495, 10), 497 => to_unsigned(587, 10), 498 => to_unsigned(874, 10), 499 => to_unsigned(152, 10), 500 => to_unsigned(321, 10), 501 => to_unsigned(237, 10), 502 => to_unsigned(957, 10), 503 => to_unsigned(144, 10), 504 => to_unsigned(782, 10), 505 => to_unsigned(453, 10), 506 => to_unsigned(979, 10), 507 => to_unsigned(525, 10), 508 => to_unsigned(785, 10), 509 => to_unsigned(421, 10), 510 => to_unsigned(619, 10), 511 => to_unsigned(795, 10), 512 => to_unsigned(813, 10), 513 => to_unsigned(73, 10), 514 => to_unsigned(305, 10), 515 => to_unsigned(165, 10), 516 => to_unsigned(61, 10), 517 => to_unsigned(784, 10), 518 => to_unsigned(433, 10), 519 => to_unsigned(458, 10), 520 => to_unsigned(921, 10), 521 => to_unsigned(636, 10), 522 => to_unsigned(664, 10), 523 => to_unsigned(101, 10), 524 => to_unsigned(389, 10), 525 => to_unsigned(58, 10), 526 => to_unsigned(128, 10), 527 => to_unsigned(842, 10), 528 => to_unsigned(429, 10), 529 => to_unsigned(551, 10), 530 => to_unsigned(946, 10), 531 => to_unsigned(908, 10), 532 => to_unsigned(470, 10), 533 => to_unsigned(278, 10), 534 => to_unsigned(313, 10), 535 => to_unsigned(448, 10), 536 => to_unsigned(482, 10), 537 => to_unsigned(645, 10), 538 => to_unsigned(897, 10), 539 => to_unsigned(963, 10), 540 => to_unsigned(334, 10), 541 => to_unsigned(382, 10), 542 => to_unsigned(856, 10), 543 => to_unsigned(306, 10), 544 => to_unsigned(301, 10), 545 => to_unsigned(867, 10), 546 => to_unsigned(714, 10), 547 => to_unsigned(860, 10), 548 => to_unsigned(596, 10), 549 => to_unsigned(623, 10), 550 => to_unsigned(829, 10), 551 => to_unsigned(947, 10), 552 => to_unsigned(272, 10), 553 => to_unsigned(538, 10), 554 => to_unsigned(261, 10), 555 => to_unsigned(413, 10), 556 => to_unsigned(596, 10), 557 => to_unsigned(935, 10), 558 => to_unsigned(630, 10), 559 => to_unsigned(891, 10), 560 => to_unsigned(231, 10), 561 => to_unsigned(336, 10), 562 => to_unsigned(436, 10), 563 => to_unsigned(20, 10), 564 => to_unsigned(313, 10), 565 => to_unsigned(251, 10), 566 => to_unsigned(970, 10), 567 => to_unsigned(183, 10), 568 => to_unsigned(276, 10), 569 => to_unsigned(459, 10), 570 => to_unsigned(140, 10), 571 => to_unsigned(625, 10), 572 => to_unsigned(725, 10), 573 => to_unsigned(145, 10), 574 => to_unsigned(61, 10), 575 => to_unsigned(833, 10), 576 => to_unsigned(79, 10), 577 => to_unsigned(976, 10), 578 => to_unsigned(997, 10), 579 => to_unsigned(412, 10), 580 => to_unsigned(624, 10), 581 => to_unsigned(610, 10), 582 => to_unsigned(91, 10), 583 => to_unsigned(682, 10), 584 => to_unsigned(216, 10), 585 => to_unsigned(879, 10), 586 => to_unsigned(723, 10), 587 => to_unsigned(718, 10), 588 => to_unsigned(631, 10), 589 => to_unsigned(580, 10), 590 => to_unsigned(241, 10), 591 => to_unsigned(950, 10), 592 => to_unsigned(302, 10), 593 => to_unsigned(451, 10), 594 => to_unsigned(854, 10), 595 => to_unsigned(336, 10), 596 => to_unsigned(78, 10), 597 => to_unsigned(369, 10), 598 => to_unsigned(579, 10), 599 => to_unsigned(687, 10), 600 => to_unsigned(337, 10), 601 => to_unsigned(726, 10), 602 => to_unsigned(805, 10), 603 => to_unsigned(590, 10), 604 => to_unsigned(169, 10), 605 => to_unsigned(87, 10), 606 => to_unsigned(632, 10), 607 => to_unsigned(624, 10), 608 => to_unsigned(353, 10), 609 => to_unsigned(499, 10), 610 => to_unsigned(644, 10), 611 => to_unsigned(771, 10), 612 => to_unsigned(938, 10), 613 => to_unsigned(418, 10), 614 => to_unsigned(376, 10), 615 => to_unsigned(356, 10), 616 => to_unsigned(860, 10), 617 => to_unsigned(695, 10), 618 => to_unsigned(396, 10), 619 => to_unsigned(487, 10), 620 => to_unsigned(204, 10), 621 => to_unsigned(454, 10), 622 => to_unsigned(221, 10), 623 => to_unsigned(456, 10), 624 => to_unsigned(25, 10), 625 => to_unsigned(537, 10), 626 => to_unsigned(278, 10), 627 => to_unsigned(5, 10), 628 => to_unsigned(371, 10), 629 => to_unsigned(819, 10), 630 => to_unsigned(136, 10), 631 => to_unsigned(381, 10), 632 => to_unsigned(726, 10), 633 => to_unsigned(828, 10), 634 => to_unsigned(372, 10), 635 => to_unsigned(650, 10), 636 => to_unsigned(23, 10), 637 => to_unsigned(597, 10), 638 => to_unsigned(507, 10), 639 => to_unsigned(311, 10), 640 => to_unsigned(881, 10), 641 => to_unsigned(427, 10), 642 => to_unsigned(278, 10), 643 => to_unsigned(812, 10), 644 => to_unsigned(492, 10), 645 => to_unsigned(264, 10), 646 => to_unsigned(81, 10), 647 => to_unsigned(367, 10), 648 => to_unsigned(923, 10), 649 => to_unsigned(851, 10), 650 => to_unsigned(601, 10), 651 => to_unsigned(177, 10), 652 => to_unsigned(1001, 10), 653 => to_unsigned(622, 10), 654 => to_unsigned(382, 10), 655 => to_unsigned(443, 10), 656 => to_unsigned(596, 10), 657 => to_unsigned(779, 10), 658 => to_unsigned(352, 10), 659 => to_unsigned(513, 10), 660 => to_unsigned(462, 10), 661 => to_unsigned(641, 10), 662 => to_unsigned(101, 10), 663 => to_unsigned(101, 10), 664 => to_unsigned(617, 10), 665 => to_unsigned(179, 10), 666 => to_unsigned(378, 10), 667 => to_unsigned(553, 10), 668 => to_unsigned(624, 10), 669 => to_unsigned(562, 10), 670 => to_unsigned(921, 10), 671 => to_unsigned(874, 10), 672 => to_unsigned(125, 10), 673 => to_unsigned(608, 10), 674 => to_unsigned(635, 10), 675 => to_unsigned(214, 10), 676 => to_unsigned(887, 10), 677 => to_unsigned(80, 10), 678 => to_unsigned(403, 10), 679 => to_unsigned(321, 10), 680 => to_unsigned(524, 10), 681 => to_unsigned(259, 10), 682 => to_unsigned(181, 10), 683 => to_unsigned(794, 10), 684 => to_unsigned(496, 10), 685 => to_unsigned(650, 10), 686 => to_unsigned(176, 10), 687 => to_unsigned(229, 10), 688 => to_unsigned(179, 10), 689 => to_unsigned(713, 10), 690 => to_unsigned(974, 10), 691 => to_unsigned(758, 10), 692 => to_unsigned(480, 10), 693 => to_unsigned(255, 10), 694 => to_unsigned(720, 10), 695 => to_unsigned(240, 10), 696 => to_unsigned(519, 10), 697 => to_unsigned(684, 10), 698 => to_unsigned(433, 10), 699 => to_unsigned(170, 10), 700 => to_unsigned(155, 10), 701 => to_unsigned(161, 10), 702 => to_unsigned(349, 10), 703 => to_unsigned(915, 10), 704 => to_unsigned(544, 10), 705 => to_unsigned(13, 10), 706 => to_unsigned(30, 10), 707 => to_unsigned(712, 10), 708 => to_unsigned(314, 10), 709 => to_unsigned(519, 10), 710 => to_unsigned(578, 10), 711 => to_unsigned(431, 10), 712 => to_unsigned(731, 10), 713 => to_unsigned(663, 10), 714 => to_unsigned(728, 10), 715 => to_unsigned(499, 10), 716 => to_unsigned(1015, 10), 717 => to_unsigned(311, 10), 718 => to_unsigned(158, 10), 719 => to_unsigned(284, 10), 720 => to_unsigned(324, 10), 721 => to_unsigned(676, 10), 722 => to_unsigned(423, 10), 723 => to_unsigned(604, 10), 724 => to_unsigned(168, 10), 725 => to_unsigned(511, 10), 726 => to_unsigned(892, 10), 727 => to_unsigned(50, 10), 728 => to_unsigned(826, 10), 729 => to_unsigned(731, 10), 730 => to_unsigned(810, 10), 731 => to_unsigned(946, 10), 732 => to_unsigned(55, 10), 733 => to_unsigned(153, 10), 734 => to_unsigned(66, 10), 735 => to_unsigned(729, 10), 736 => to_unsigned(275, 10), 737 => to_unsigned(201, 10), 738 => to_unsigned(81, 10), 739 => to_unsigned(939, 10), 740 => to_unsigned(272, 10), 741 => to_unsigned(1013, 10), 742 => to_unsigned(985, 10), 743 => to_unsigned(786, 10), 744 => to_unsigned(822, 10), 745 => to_unsigned(518, 10), 746 => to_unsigned(187, 10), 747 => to_unsigned(333, 10), 748 => to_unsigned(768, 10), 749 => to_unsigned(800, 10), 750 => to_unsigned(255, 10), 751 => to_unsigned(190, 10), 752 => to_unsigned(363, 10), 753 => to_unsigned(312, 10), 754 => to_unsigned(251, 10), 755 => to_unsigned(629, 10), 756 => to_unsigned(766, 10), 757 => to_unsigned(437, 10), 758 => to_unsigned(241, 10), 759 => to_unsigned(549, 10), 760 => to_unsigned(982, 10), 761 => to_unsigned(507, 10), 762 => to_unsigned(104, 10), 763 => to_unsigned(295, 10), 764 => to_unsigned(772, 10), 765 => to_unsigned(450, 10), 766 => to_unsigned(503, 10), 767 => to_unsigned(393, 10), 768 => to_unsigned(588, 10), 769 => to_unsigned(92, 10), 770 => to_unsigned(37, 10), 771 => to_unsigned(451, 10), 772 => to_unsigned(82, 10), 773 => to_unsigned(147, 10), 774 => to_unsigned(733, 10), 775 => to_unsigned(193, 10), 776 => to_unsigned(885, 10), 777 => to_unsigned(944, 10), 778 => to_unsigned(137, 10), 779 => to_unsigned(463, 10), 780 => to_unsigned(972, 10), 781 => to_unsigned(449, 10), 782 => to_unsigned(554, 10), 783 => to_unsigned(359, 10), 784 => to_unsigned(51, 10), 785 => to_unsigned(276, 10), 786 => to_unsigned(16, 10), 787 => to_unsigned(102, 10), 788 => to_unsigned(902, 10), 789 => to_unsigned(976, 10), 790 => to_unsigned(976, 10), 791 => to_unsigned(554, 10), 792 => to_unsigned(97, 10), 793 => to_unsigned(6, 10), 794 => to_unsigned(666, 10), 795 => to_unsigned(472, 10), 796 => to_unsigned(186, 10), 797 => to_unsigned(346, 10), 798 => to_unsigned(473, 10), 799 => to_unsigned(913, 10), 800 => to_unsigned(707, 10), 801 => to_unsigned(442, 10), 802 => to_unsigned(817, 10), 803 => to_unsigned(158, 10), 804 => to_unsigned(139, 10), 805 => to_unsigned(20, 10), 806 => to_unsigned(933, 10), 807 => to_unsigned(999, 10), 808 => to_unsigned(826, 10), 809 => to_unsigned(657, 10), 810 => to_unsigned(251, 10), 811 => to_unsigned(998, 10), 812 => to_unsigned(87, 10), 813 => to_unsigned(730, 10), 814 => to_unsigned(369, 10), 815 => to_unsigned(895, 10), 816 => to_unsigned(519, 10), 817 => to_unsigned(960, 10), 818 => to_unsigned(766, 10), 819 => to_unsigned(909, 10), 820 => to_unsigned(972, 10), 821 => to_unsigned(556, 10), 822 => to_unsigned(533, 10), 823 => to_unsigned(868, 10), 824 => to_unsigned(664, 10), 825 => to_unsigned(380, 10), 826 => to_unsigned(301, 10), 827 => to_unsigned(253, 10), 828 => to_unsigned(324, 10), 829 => to_unsigned(956, 10), 830 => to_unsigned(420, 10), 831 => to_unsigned(425, 10), 832 => to_unsigned(1008, 10), 833 => to_unsigned(826, 10), 834 => to_unsigned(794, 10), 835 => to_unsigned(929, 10), 836 => to_unsigned(368, 10), 837 => to_unsigned(459, 10), 838 => to_unsigned(54, 10), 839 => to_unsigned(912, 10), 840 => to_unsigned(231, 10), 841 => to_unsigned(75, 10), 842 => to_unsigned(874, 10), 843 => to_unsigned(877, 10), 844 => to_unsigned(263, 10), 845 => to_unsigned(861, 10), 846 => to_unsigned(907, 10), 847 => to_unsigned(160, 10), 848 => to_unsigned(312, 10), 849 => to_unsigned(60, 10), 850 => to_unsigned(640, 10), 851 => to_unsigned(408, 10), 852 => to_unsigned(484, 10), 853 => to_unsigned(815, 10), 854 => to_unsigned(350, 10), 855 => to_unsigned(378, 10), 856 => to_unsigned(460, 10), 857 => to_unsigned(348, 10), 858 => to_unsigned(614, 10), 859 => to_unsigned(186, 10), 860 => to_unsigned(626, 10), 861 => to_unsigned(863, 10), 862 => to_unsigned(387, 10), 863 => to_unsigned(842, 10), 864 => to_unsigned(968, 10), 865 => to_unsigned(412, 10), 866 => to_unsigned(985, 10), 867 => to_unsigned(110, 10), 868 => to_unsigned(75, 10), 869 => to_unsigned(954, 10), 870 => to_unsigned(378, 10), 871 => to_unsigned(68, 10), 872 => to_unsigned(221, 10), 873 => to_unsigned(795, 10), 874 => to_unsigned(912, 10), 875 => to_unsigned(38, 10), 876 => to_unsigned(7, 10), 877 => to_unsigned(282, 10), 878 => to_unsigned(177, 10), 879 => to_unsigned(603, 10), 880 => to_unsigned(954, 10), 881 => to_unsigned(49, 10), 882 => to_unsigned(604, 10), 883 => to_unsigned(975, 10), 884 => to_unsigned(466, 10), 885 => to_unsigned(158, 10), 886 => to_unsigned(51, 10), 887 => to_unsigned(83, 10), 888 => to_unsigned(480, 10), 889 => to_unsigned(569, 10), 890 => to_unsigned(411, 10), 891 => to_unsigned(375, 10), 892 => to_unsigned(509, 10), 893 => to_unsigned(382, 10), 894 => to_unsigned(72, 10), 895 => to_unsigned(388, 10), 896 => to_unsigned(411, 10), 897 => to_unsigned(551, 10), 898 => to_unsigned(705, 10), 899 => to_unsigned(913, 10), 900 => to_unsigned(841, 10), 901 => to_unsigned(437, 10), 902 => to_unsigned(226, 10), 903 => to_unsigned(726, 10), 904 => to_unsigned(628, 10), 905 => to_unsigned(64, 10), 906 => to_unsigned(732, 10), 907 => to_unsigned(992, 10), 908 => to_unsigned(547, 10), 909 => to_unsigned(34, 10), 910 => to_unsigned(867, 10), 911 => to_unsigned(847, 10), 912 => to_unsigned(49, 10), 913 => to_unsigned(472, 10), 914 => to_unsigned(860, 10), 915 => to_unsigned(886, 10), 916 => to_unsigned(646, 10), 917 => to_unsigned(144, 10), 918 => to_unsigned(456, 10), 919 => to_unsigned(721, 10), 920 => to_unsigned(441, 10), 921 => to_unsigned(162, 10), 922 => to_unsigned(66, 10), 923 => to_unsigned(776, 10), 924 => to_unsigned(587, 10), 925 => to_unsigned(104, 10), 926 => to_unsigned(560, 10), 927 => to_unsigned(568, 10), 928 => to_unsigned(199, 10), 929 => to_unsigned(217, 10), 930 => to_unsigned(311, 10), 931 => to_unsigned(724, 10), 932 => to_unsigned(619, 10), 933 => to_unsigned(166, 10), 934 => to_unsigned(176, 10), 935 => to_unsigned(753, 10), 936 => to_unsigned(249, 10), 937 => to_unsigned(727, 10), 938 => to_unsigned(98, 10), 939 => to_unsigned(636, 10), 940 => to_unsigned(996, 10), 941 => to_unsigned(641, 10), 942 => to_unsigned(112, 10), 943 => to_unsigned(1013, 10), 944 => to_unsigned(855, 10), 945 => to_unsigned(1009, 10), 946 => to_unsigned(110, 10), 947 => to_unsigned(698, 10), 948 => to_unsigned(900, 10), 949 => to_unsigned(425, 10), 950 => to_unsigned(492, 10), 951 => to_unsigned(525, 10), 952 => to_unsigned(172, 10), 953 => to_unsigned(910, 10), 954 => to_unsigned(738, 10), 955 => to_unsigned(32, 10), 956 => to_unsigned(243, 10), 957 => to_unsigned(688, 10), 958 => to_unsigned(312, 10), 959 => to_unsigned(481, 10), 960 => to_unsigned(784, 10), 961 => to_unsigned(130, 10), 962 => to_unsigned(710, 10), 963 => to_unsigned(404, 10), 964 => to_unsigned(935, 10), 965 => to_unsigned(1023, 10), 966 => to_unsigned(550, 10), 967 => to_unsigned(642, 10), 968 => to_unsigned(434, 10), 969 => to_unsigned(393, 10), 970 => to_unsigned(90, 10), 971 => to_unsigned(112, 10), 972 => to_unsigned(574, 10), 973 => to_unsigned(233, 10), 974 => to_unsigned(121, 10), 975 => to_unsigned(611, 10), 976 => to_unsigned(167, 10), 977 => to_unsigned(659, 10), 978 => to_unsigned(115, 10), 979 => to_unsigned(227, 10), 980 => to_unsigned(972, 10), 981 => to_unsigned(513, 10), 982 => to_unsigned(152, 10), 983 => to_unsigned(987, 10), 984 => to_unsigned(320, 10), 985 => to_unsigned(10, 10), 986 => to_unsigned(547, 10), 987 => to_unsigned(707, 10), 988 => to_unsigned(281, 10), 989 => to_unsigned(155, 10), 990 => to_unsigned(182, 10), 991 => to_unsigned(89, 10), 992 => to_unsigned(761, 10), 993 => to_unsigned(267, 10), 994 => to_unsigned(208, 10), 995 => to_unsigned(342, 10), 996 => to_unsigned(703, 10), 997 => to_unsigned(520, 10), 998 => to_unsigned(994, 10), 999 => to_unsigned(20, 10), 1000 => to_unsigned(312, 10), 1001 => to_unsigned(832, 10), 1002 => to_unsigned(477, 10), 1003 => to_unsigned(443, 10), 1004 => to_unsigned(735, 10), 1005 => to_unsigned(613, 10), 1006 => to_unsigned(539, 10), 1007 => to_unsigned(166, 10), 1008 => to_unsigned(971, 10), 1009 => to_unsigned(302, 10), 1010 => to_unsigned(904, 10), 1011 => to_unsigned(296, 10), 1012 => to_unsigned(418, 10), 1013 => to_unsigned(1017, 10), 1014 => to_unsigned(648, 10), 1015 => to_unsigned(888, 10), 1016 => to_unsigned(51, 10), 1017 => to_unsigned(797, 10), 1018 => to_unsigned(99, 10), 1019 => to_unsigned(701, 10), 1020 => to_unsigned(215, 10), 1021 => to_unsigned(92, 10), 1022 => to_unsigned(292, 10), 1023 => to_unsigned(175, 10), 1024 => to_unsigned(853, 10), 1025 => to_unsigned(407, 10), 1026 => to_unsigned(363, 10), 1027 => to_unsigned(926, 10), 1028 => to_unsigned(549, 10), 1029 => to_unsigned(25, 10), 1030 => to_unsigned(812, 10), 1031 => to_unsigned(260, 10), 1032 => to_unsigned(404, 10), 1033 => to_unsigned(252, 10), 1034 => to_unsigned(379, 10), 1035 => to_unsigned(92, 10), 1036 => to_unsigned(793, 10), 1037 => to_unsigned(836, 10), 1038 => to_unsigned(207, 10), 1039 => to_unsigned(898, 10), 1040 => to_unsigned(839, 10), 1041 => to_unsigned(304, 10), 1042 => to_unsigned(450, 10), 1043 => to_unsigned(223, 10), 1044 => to_unsigned(666, 10), 1045 => to_unsigned(959, 10), 1046 => to_unsigned(895, 10), 1047 => to_unsigned(774, 10), 1048 => to_unsigned(2, 10), 1049 => to_unsigned(875, 10), 1050 => to_unsigned(365, 10), 1051 => to_unsigned(985, 10), 1052 => to_unsigned(59, 10), 1053 => to_unsigned(614, 10), 1054 => to_unsigned(399, 10), 1055 => to_unsigned(379, 10), 1056 => to_unsigned(923, 10), 1057 => to_unsigned(667, 10), 1058 => to_unsigned(220, 10), 1059 => to_unsigned(729, 10), 1060 => to_unsigned(192, 10), 1061 => to_unsigned(294, 10), 1062 => to_unsigned(187, 10), 1063 => to_unsigned(395, 10), 1064 => to_unsigned(277, 10), 1065 => to_unsigned(774, 10), 1066 => to_unsigned(47, 10), 1067 => to_unsigned(153, 10), 1068 => to_unsigned(1015, 10), 1069 => to_unsigned(915, 10), 1070 => to_unsigned(306, 10), 1071 => to_unsigned(259, 10), 1072 => to_unsigned(608, 10), 1073 => to_unsigned(402, 10), 1074 => to_unsigned(669, 10), 1075 => to_unsigned(890, 10), 1076 => to_unsigned(64, 10), 1077 => to_unsigned(140, 10), 1078 => to_unsigned(44, 10), 1079 => to_unsigned(227, 10), 1080 => to_unsigned(744, 10), 1081 => to_unsigned(312, 10), 1082 => to_unsigned(75, 10), 1083 => to_unsigned(771, 10), 1084 => to_unsigned(685, 10), 1085 => to_unsigned(569, 10), 1086 => to_unsigned(157, 10), 1087 => to_unsigned(410, 10), 1088 => to_unsigned(648, 10), 1089 => to_unsigned(449, 10), 1090 => to_unsigned(961, 10), 1091 => to_unsigned(1012, 10), 1092 => to_unsigned(582, 10), 1093 => to_unsigned(511, 10), 1094 => to_unsigned(472, 10), 1095 => to_unsigned(952, 10), 1096 => to_unsigned(847, 10), 1097 => to_unsigned(74, 10), 1098 => to_unsigned(786, 10), 1099 => to_unsigned(628, 10), 1100 => to_unsigned(214, 10), 1101 => to_unsigned(681, 10), 1102 => to_unsigned(841, 10), 1103 => to_unsigned(71, 10), 1104 => to_unsigned(321, 10), 1105 => to_unsigned(965, 10), 1106 => to_unsigned(393, 10), 1107 => to_unsigned(133, 10), 1108 => to_unsigned(623, 10), 1109 => to_unsigned(687, 10), 1110 => to_unsigned(756, 10), 1111 => to_unsigned(52, 10), 1112 => to_unsigned(191, 10), 1113 => to_unsigned(942, 10), 1114 => to_unsigned(979, 10), 1115 => to_unsigned(939, 10), 1116 => to_unsigned(92, 10), 1117 => to_unsigned(936, 10), 1118 => to_unsigned(621, 10), 1119 => to_unsigned(210, 10), 1120 => to_unsigned(587, 10), 1121 => to_unsigned(198, 10), 1122 => to_unsigned(178, 10), 1123 => to_unsigned(531, 10), 1124 => to_unsigned(246, 10), 1125 => to_unsigned(329, 10), 1126 => to_unsigned(947, 10), 1127 => to_unsigned(827, 10), 1128 => to_unsigned(353, 10), 1129 => to_unsigned(276, 10), 1130 => to_unsigned(482, 10), 1131 => to_unsigned(1016, 10), 1132 => to_unsigned(332, 10), 1133 => to_unsigned(573, 10), 1134 => to_unsigned(457, 10), 1135 => to_unsigned(860, 10), 1136 => to_unsigned(835, 10), 1137 => to_unsigned(976, 10), 1138 => to_unsigned(302, 10), 1139 => to_unsigned(781, 10), 1140 => to_unsigned(560, 10), 1141 => to_unsigned(372, 10), 1142 => to_unsigned(309, 10), 1143 => to_unsigned(319, 10), 1144 => to_unsigned(174, 10), 1145 => to_unsigned(181, 10), 1146 => to_unsigned(723, 10), 1147 => to_unsigned(243, 10), 1148 => to_unsigned(929, 10), 1149 => to_unsigned(656, 10), 1150 => to_unsigned(296, 10), 1151 => to_unsigned(514, 10), 1152 => to_unsigned(573, 10), 1153 => to_unsigned(399, 10), 1154 => to_unsigned(848, 10), 1155 => to_unsigned(756, 10), 1156 => to_unsigned(880, 10), 1157 => to_unsigned(181, 10), 1158 => to_unsigned(907, 10), 1159 => to_unsigned(133, 10), 1160 => to_unsigned(191, 10), 1161 => to_unsigned(468, 10), 1162 => to_unsigned(463, 10), 1163 => to_unsigned(61, 10), 1164 => to_unsigned(653, 10), 1165 => to_unsigned(27, 10), 1166 => to_unsigned(150, 10), 1167 => to_unsigned(126, 10), 1168 => to_unsigned(762, 10), 1169 => to_unsigned(342, 10), 1170 => to_unsigned(711, 10), 1171 => to_unsigned(42, 10), 1172 => to_unsigned(663, 10), 1173 => to_unsigned(472, 10), 1174 => to_unsigned(865, 10), 1175 => to_unsigned(854, 10), 1176 => to_unsigned(230, 10), 1177 => to_unsigned(900, 10), 1178 => to_unsigned(867, 10), 1179 => to_unsigned(37, 10), 1180 => to_unsigned(612, 10), 1181 => to_unsigned(673, 10), 1182 => to_unsigned(630, 10), 1183 => to_unsigned(116, 10), 1184 => to_unsigned(941, 10), 1185 => to_unsigned(552, 10), 1186 => to_unsigned(36, 10), 1187 => to_unsigned(533, 10), 1188 => to_unsigned(860, 10), 1189 => to_unsigned(40, 10), 1190 => to_unsigned(60, 10), 1191 => to_unsigned(986, 10), 1192 => to_unsigned(133, 10), 1193 => to_unsigned(465, 10), 1194 => to_unsigned(203, 10), 1195 => to_unsigned(773, 10), 1196 => to_unsigned(983, 10), 1197 => to_unsigned(943, 10), 1198 => to_unsigned(355, 10), 1199 => to_unsigned(629, 10), 1200 => to_unsigned(797, 10), 1201 => to_unsigned(513, 10), 1202 => to_unsigned(180, 10), 1203 => to_unsigned(665, 10), 1204 => to_unsigned(55, 10), 1205 => to_unsigned(164, 10), 1206 => to_unsigned(727, 10), 1207 => to_unsigned(346, 10), 1208 => to_unsigned(770, 10), 1209 => to_unsigned(25, 10), 1210 => to_unsigned(76, 10), 1211 => to_unsigned(954, 10), 1212 => to_unsigned(948, 10), 1213 => to_unsigned(634, 10), 1214 => to_unsigned(52, 10), 1215 => to_unsigned(534, 10), 1216 => to_unsigned(331, 10), 1217 => to_unsigned(375, 10), 1218 => to_unsigned(865, 10), 1219 => to_unsigned(567, 10), 1220 => to_unsigned(21, 10), 1221 => to_unsigned(442, 10), 1222 => to_unsigned(417, 10), 1223 => to_unsigned(102, 10), 1224 => to_unsigned(951, 10), 1225 => to_unsigned(698, 10), 1226 => to_unsigned(856, 10), 1227 => to_unsigned(418, 10), 1228 => to_unsigned(264, 10), 1229 => to_unsigned(62, 10), 1230 => to_unsigned(904, 10), 1231 => to_unsigned(934, 10), 1232 => to_unsigned(96, 10), 1233 => to_unsigned(717, 10), 1234 => to_unsigned(291, 10), 1235 => to_unsigned(158, 10), 1236 => to_unsigned(127, 10), 1237 => to_unsigned(359, 10), 1238 => to_unsigned(638, 10), 1239 => to_unsigned(1008, 10), 1240 => to_unsigned(969, 10), 1241 => to_unsigned(381, 10), 1242 => to_unsigned(365, 10), 1243 => to_unsigned(404, 10), 1244 => to_unsigned(720, 10), 1245 => to_unsigned(271, 10), 1246 => to_unsigned(869, 10), 1247 => to_unsigned(88, 10), 1248 => to_unsigned(179, 10), 1249 => to_unsigned(477, 10), 1250 => to_unsigned(491, 10), 1251 => to_unsigned(464, 10), 1252 => to_unsigned(266, 10), 1253 => to_unsigned(68, 10), 1254 => to_unsigned(148, 10), 1255 => to_unsigned(472, 10), 1256 => to_unsigned(727, 10), 1257 => to_unsigned(557, 10), 1258 => to_unsigned(612, 10), 1259 => to_unsigned(117, 10), 1260 => to_unsigned(510, 10), 1261 => to_unsigned(413, 10), 1262 => to_unsigned(811, 10), 1263 => to_unsigned(179, 10), 1264 => to_unsigned(405, 10), 1265 => to_unsigned(842, 10), 1266 => to_unsigned(106, 10), 1267 => to_unsigned(889, 10), 1268 => to_unsigned(642, 10), 1269 => to_unsigned(325, 10), 1270 => to_unsigned(493, 10), 1271 => to_unsigned(712, 10), 1272 => to_unsigned(150, 10), 1273 => to_unsigned(226, 10), 1274 => to_unsigned(228, 10), 1275 => to_unsigned(557, 10), 1276 => to_unsigned(224, 10), 1277 => to_unsigned(43, 10), 1278 => to_unsigned(122, 10), 1279 => to_unsigned(707, 10), 1280 => to_unsigned(30, 10), 1281 => to_unsigned(42, 10), 1282 => to_unsigned(940, 10), 1283 => to_unsigned(630, 10), 1284 => to_unsigned(417, 10), 1285 => to_unsigned(303, 10), 1286 => to_unsigned(739, 10), 1287 => to_unsigned(49, 10), 1288 => to_unsigned(289, 10), 1289 => to_unsigned(356, 10), 1290 => to_unsigned(552, 10), 1291 => to_unsigned(905, 10), 1292 => to_unsigned(1, 10), 1293 => to_unsigned(381, 10), 1294 => to_unsigned(47, 10), 1295 => to_unsigned(532, 10), 1296 => to_unsigned(902, 10), 1297 => to_unsigned(715, 10), 1298 => to_unsigned(763, 10), 1299 => to_unsigned(419, 10), 1300 => to_unsigned(292, 10), 1301 => to_unsigned(385, 10), 1302 => to_unsigned(939, 10), 1303 => to_unsigned(69, 10), 1304 => to_unsigned(759, 10), 1305 => to_unsigned(190, 10), 1306 => to_unsigned(83, 10), 1307 => to_unsigned(741, 10), 1308 => to_unsigned(859, 10), 1309 => to_unsigned(870, 10), 1310 => to_unsigned(507, 10), 1311 => to_unsigned(770, 10), 1312 => to_unsigned(153, 10), 1313 => to_unsigned(705, 10), 1314 => to_unsigned(961, 10), 1315 => to_unsigned(888, 10), 1316 => to_unsigned(525, 10), 1317 => to_unsigned(588, 10), 1318 => to_unsigned(311, 10), 1319 => to_unsigned(633, 10), 1320 => to_unsigned(139, 10), 1321 => to_unsigned(147, 10), 1322 => to_unsigned(723, 10), 1323 => to_unsigned(768, 10), 1324 => to_unsigned(254, 10), 1325 => to_unsigned(817, 10), 1326 => to_unsigned(171, 10), 1327 => to_unsigned(656, 10), 1328 => to_unsigned(161, 10), 1329 => to_unsigned(745, 10), 1330 => to_unsigned(467, 10), 1331 => to_unsigned(281, 10), 1332 => to_unsigned(451, 10), 1333 => to_unsigned(962, 10), 1334 => to_unsigned(902, 10), 1335 => to_unsigned(435, 10), 1336 => to_unsigned(585, 10), 1337 => to_unsigned(640, 10), 1338 => to_unsigned(975, 10), 1339 => to_unsigned(1007, 10), 1340 => to_unsigned(103, 10), 1341 => to_unsigned(198, 10), 1342 => to_unsigned(542, 10), 1343 => to_unsigned(787, 10), 1344 => to_unsigned(274, 10), 1345 => to_unsigned(486, 10), 1346 => to_unsigned(321, 10), 1347 => to_unsigned(725, 10), 1348 => to_unsigned(158, 10), 1349 => to_unsigned(616, 10), 1350 => to_unsigned(674, 10), 1351 => to_unsigned(785, 10), 1352 => to_unsigned(104, 10), 1353 => to_unsigned(640, 10), 1354 => to_unsigned(981, 10), 1355 => to_unsigned(413, 10), 1356 => to_unsigned(178, 10), 1357 => to_unsigned(512, 10), 1358 => to_unsigned(157, 10), 1359 => to_unsigned(867, 10), 1360 => to_unsigned(128, 10), 1361 => to_unsigned(957, 10), 1362 => to_unsigned(637, 10), 1363 => to_unsigned(102, 10), 1364 => to_unsigned(462, 10), 1365 => to_unsigned(248, 10), 1366 => to_unsigned(483, 10), 1367 => to_unsigned(948, 10), 1368 => to_unsigned(86, 10), 1369 => to_unsigned(788, 10), 1370 => to_unsigned(432, 10), 1371 => to_unsigned(797, 10), 1372 => to_unsigned(892, 10), 1373 => to_unsigned(398, 10), 1374 => to_unsigned(818, 10), 1375 => to_unsigned(231, 10), 1376 => to_unsigned(724, 10), 1377 => to_unsigned(279, 10), 1378 => to_unsigned(419, 10), 1379 => to_unsigned(204, 10), 1380 => to_unsigned(171, 10), 1381 => to_unsigned(617, 10), 1382 => to_unsigned(693, 10), 1383 => to_unsigned(157, 10), 1384 => to_unsigned(258, 10), 1385 => to_unsigned(689, 10), 1386 => to_unsigned(326, 10), 1387 => to_unsigned(56, 10), 1388 => to_unsigned(49, 10), 1389 => to_unsigned(1023, 10), 1390 => to_unsigned(486, 10), 1391 => to_unsigned(445, 10), 1392 => to_unsigned(301, 10), 1393 => to_unsigned(819, 10), 1394 => to_unsigned(116, 10), 1395 => to_unsigned(30, 10), 1396 => to_unsigned(307, 10), 1397 => to_unsigned(377, 10), 1398 => to_unsigned(166, 10), 1399 => to_unsigned(260, 10), 1400 => to_unsigned(801, 10), 1401 => to_unsigned(636, 10), 1402 => to_unsigned(383, 10), 1403 => to_unsigned(623, 10), 1404 => to_unsigned(28, 10), 1405 => to_unsigned(958, 10), 1406 => to_unsigned(984, 10), 1407 => to_unsigned(41, 10), 1408 => to_unsigned(567, 10), 1409 => to_unsigned(1008, 10), 1410 => to_unsigned(451, 10), 1411 => to_unsigned(657, 10), 1412 => to_unsigned(685, 10), 1413 => to_unsigned(773, 10), 1414 => to_unsigned(993, 10), 1415 => to_unsigned(458, 10), 1416 => to_unsigned(0, 10), 1417 => to_unsigned(545, 10), 1418 => to_unsigned(338, 10), 1419 => to_unsigned(834, 10), 1420 => to_unsigned(109, 10), 1421 => to_unsigned(3, 10), 1422 => to_unsigned(511, 10), 1423 => to_unsigned(147, 10), 1424 => to_unsigned(91, 10), 1425 => to_unsigned(882, 10), 1426 => to_unsigned(362, 10), 1427 => to_unsigned(530, 10), 1428 => to_unsigned(680, 10), 1429 => to_unsigned(219, 10), 1430 => to_unsigned(954, 10), 1431 => to_unsigned(761, 10), 1432 => to_unsigned(388, 10), 1433 => to_unsigned(268, 10), 1434 => to_unsigned(657, 10), 1435 => to_unsigned(21, 10), 1436 => to_unsigned(435, 10), 1437 => to_unsigned(478, 10), 1438 => to_unsigned(118, 10), 1439 => to_unsigned(614, 10), 1440 => to_unsigned(1001, 10), 1441 => to_unsigned(10, 10), 1442 => to_unsigned(99, 10), 1443 => to_unsigned(569, 10), 1444 => to_unsigned(425, 10), 1445 => to_unsigned(188, 10), 1446 => to_unsigned(916, 10), 1447 => to_unsigned(597, 10), 1448 => to_unsigned(840, 10), 1449 => to_unsigned(946, 10), 1450 => to_unsigned(249, 10), 1451 => to_unsigned(401, 10), 1452 => to_unsigned(261, 10), 1453 => to_unsigned(526, 10), 1454 => to_unsigned(164, 10), 1455 => to_unsigned(209, 10), 1456 => to_unsigned(485, 10), 1457 => to_unsigned(535, 10), 1458 => to_unsigned(439, 10), 1459 => to_unsigned(662, 10), 1460 => to_unsigned(349, 10), 1461 => to_unsigned(273, 10), 1462 => to_unsigned(467, 10), 1463 => to_unsigned(775, 10), 1464 => to_unsigned(641, 10), 1465 => to_unsigned(559, 10), 1466 => to_unsigned(598, 10), 1467 => to_unsigned(649, 10), 1468 => to_unsigned(776, 10), 1469 => to_unsigned(339, 10), 1470 => to_unsigned(319, 10), 1471 => to_unsigned(748, 10), 1472 => to_unsigned(921, 10), 1473 => to_unsigned(819, 10), 1474 => to_unsigned(469, 10), 1475 => to_unsigned(282, 10), 1476 => to_unsigned(383, 10), 1477 => to_unsigned(651, 10), 1478 => to_unsigned(489, 10), 1479 => to_unsigned(14, 10), 1480 => to_unsigned(29, 10), 1481 => to_unsigned(562, 10), 1482 => to_unsigned(633, 10), 1483 => to_unsigned(246, 10), 1484 => to_unsigned(44, 10), 1485 => to_unsigned(122, 10), 1486 => to_unsigned(82, 10), 1487 => to_unsigned(478, 10), 1488 => to_unsigned(231, 10), 1489 => to_unsigned(481, 10), 1490 => to_unsigned(20, 10), 1491 => to_unsigned(34, 10), 1492 => to_unsigned(802, 10), 1493 => to_unsigned(374, 10), 1494 => to_unsigned(158, 10), 1495 => to_unsigned(559, 10), 1496 => to_unsigned(445, 10), 1497 => to_unsigned(115, 10), 1498 => to_unsigned(762, 10), 1499 => to_unsigned(469, 10), 1500 => to_unsigned(996, 10), 1501 => to_unsigned(901, 10), 1502 => to_unsigned(583, 10), 1503 => to_unsigned(960, 10), 1504 => to_unsigned(225, 10), 1505 => to_unsigned(44, 10), 1506 => to_unsigned(264, 10), 1507 => to_unsigned(836, 10), 1508 => to_unsigned(425, 10), 1509 => to_unsigned(533, 10), 1510 => to_unsigned(18, 10), 1511 => to_unsigned(765, 10), 1512 => to_unsigned(747, 10), 1513 => to_unsigned(609, 10), 1514 => to_unsigned(931, 10), 1515 => to_unsigned(919, 10), 1516 => to_unsigned(735, 10), 1517 => to_unsigned(853, 10), 1518 => to_unsigned(554, 10), 1519 => to_unsigned(1018, 10), 1520 => to_unsigned(301, 10), 1521 => to_unsigned(208, 10), 1522 => to_unsigned(572, 10), 1523 => to_unsigned(728, 10), 1524 => to_unsigned(222, 10), 1525 => to_unsigned(183, 10), 1526 => to_unsigned(972, 10), 1527 => to_unsigned(562, 10), 1528 => to_unsigned(580, 10), 1529 => to_unsigned(628, 10), 1530 => to_unsigned(409, 10), 1531 => to_unsigned(535, 10), 1532 => to_unsigned(525, 10), 1533 => to_unsigned(260, 10), 1534 => to_unsigned(987, 10), 1535 => to_unsigned(816, 10), 1536 => to_unsigned(694, 10), 1537 => to_unsigned(431, 10), 1538 => to_unsigned(426, 10), 1539 => to_unsigned(819, 10), 1540 => to_unsigned(434, 10), 1541 => to_unsigned(884, 10), 1542 => to_unsigned(831, 10), 1543 => to_unsigned(565, 10), 1544 => to_unsigned(841, 10), 1545 => to_unsigned(408, 10), 1546 => to_unsigned(684, 10), 1547 => to_unsigned(167, 10), 1548 => to_unsigned(71, 10), 1549 => to_unsigned(121, 10), 1550 => to_unsigned(1014, 10), 1551 => to_unsigned(167, 10), 1552 => to_unsigned(130, 10), 1553 => to_unsigned(22, 10), 1554 => to_unsigned(915, 10), 1555 => to_unsigned(85, 10), 1556 => to_unsigned(84, 10), 1557 => to_unsigned(208, 10), 1558 => to_unsigned(655, 10), 1559 => to_unsigned(866, 10), 1560 => to_unsigned(194, 10), 1561 => to_unsigned(101, 10), 1562 => to_unsigned(204, 10), 1563 => to_unsigned(58, 10), 1564 => to_unsigned(663, 10), 1565 => to_unsigned(524, 10), 1566 => to_unsigned(419, 10), 1567 => to_unsigned(999, 10), 1568 => to_unsigned(493, 10), 1569 => to_unsigned(62, 10), 1570 => to_unsigned(460, 10), 1571 => to_unsigned(419, 10), 1572 => to_unsigned(554, 10), 1573 => to_unsigned(827, 10), 1574 => to_unsigned(757, 10), 1575 => to_unsigned(475, 10), 1576 => to_unsigned(675, 10), 1577 => to_unsigned(825, 10), 1578 => to_unsigned(980, 10), 1579 => to_unsigned(562, 10), 1580 => to_unsigned(810, 10), 1581 => to_unsigned(175, 10), 1582 => to_unsigned(348, 10), 1583 => to_unsigned(364, 10), 1584 => to_unsigned(585, 10), 1585 => to_unsigned(172, 10), 1586 => to_unsigned(924, 10), 1587 => to_unsigned(299, 10), 1588 => to_unsigned(314, 10), 1589 => to_unsigned(477, 10), 1590 => to_unsigned(172, 10), 1591 => to_unsigned(86, 10), 1592 => to_unsigned(604, 10), 1593 => to_unsigned(684, 10), 1594 => to_unsigned(999, 10), 1595 => to_unsigned(563, 10), 1596 => to_unsigned(924, 10), 1597 => to_unsigned(675, 10), 1598 => to_unsigned(262, 10), 1599 => to_unsigned(106, 10), 1600 => to_unsigned(614, 10), 1601 => to_unsigned(297, 10), 1602 => to_unsigned(934, 10), 1603 => to_unsigned(491, 10), 1604 => to_unsigned(44, 10), 1605 => to_unsigned(242, 10), 1606 => to_unsigned(691, 10), 1607 => to_unsigned(36, 10), 1608 => to_unsigned(384, 10), 1609 => to_unsigned(64, 10), 1610 => to_unsigned(111, 10), 1611 => to_unsigned(697, 10), 1612 => to_unsigned(783, 10), 1613 => to_unsigned(900, 10), 1614 => to_unsigned(303, 10), 1615 => to_unsigned(58, 10), 1616 => to_unsigned(734, 10), 1617 => to_unsigned(109, 10), 1618 => to_unsigned(799, 10), 1619 => to_unsigned(403, 10), 1620 => to_unsigned(434, 10), 1621 => to_unsigned(225, 10), 1622 => to_unsigned(211, 10), 1623 => to_unsigned(917, 10), 1624 => to_unsigned(121, 10), 1625 => to_unsigned(990, 10), 1626 => to_unsigned(349, 10), 1627 => to_unsigned(1022, 10), 1628 => to_unsigned(218, 10), 1629 => to_unsigned(480, 10), 1630 => to_unsigned(848, 10), 1631 => to_unsigned(143, 10), 1632 => to_unsigned(356, 10), 1633 => to_unsigned(271, 10), 1634 => to_unsigned(518, 10), 1635 => to_unsigned(798, 10), 1636 => to_unsigned(187, 10), 1637 => to_unsigned(505, 10), 1638 => to_unsigned(175, 10), 1639 => to_unsigned(20, 10), 1640 => to_unsigned(221, 10), 1641 => to_unsigned(360, 10), 1642 => to_unsigned(533, 10), 1643 => to_unsigned(316, 10), 1644 => to_unsigned(671, 10), 1645 => to_unsigned(323, 10), 1646 => to_unsigned(387, 10), 1647 => to_unsigned(1021, 10), 1648 => to_unsigned(772, 10), 1649 => to_unsigned(237, 10), 1650 => to_unsigned(660, 10), 1651 => to_unsigned(829, 10), 1652 => to_unsigned(450, 10), 1653 => to_unsigned(395, 10), 1654 => to_unsigned(524, 10), 1655 => to_unsigned(933, 10), 1656 => to_unsigned(776, 10), 1657 => to_unsigned(982, 10), 1658 => to_unsigned(939, 10), 1659 => to_unsigned(168, 10), 1660 => to_unsigned(311, 10), 1661 => to_unsigned(652, 10), 1662 => to_unsigned(639, 10), 1663 => to_unsigned(986, 10), 1664 => to_unsigned(346, 10), 1665 => to_unsigned(116, 10), 1666 => to_unsigned(977, 10), 1667 => to_unsigned(935, 10), 1668 => to_unsigned(695, 10), 1669 => to_unsigned(126, 10), 1670 => to_unsigned(771, 10), 1671 => to_unsigned(133, 10), 1672 => to_unsigned(791, 10), 1673 => to_unsigned(304, 10), 1674 => to_unsigned(173, 10), 1675 => to_unsigned(999, 10), 1676 => to_unsigned(937, 10), 1677 => to_unsigned(938, 10), 1678 => to_unsigned(691, 10), 1679 => to_unsigned(814, 10), 1680 => to_unsigned(693, 10), 1681 => to_unsigned(612, 10), 1682 => to_unsigned(74, 10), 1683 => to_unsigned(372, 10), 1684 => to_unsigned(708, 10), 1685 => to_unsigned(215, 10), 1686 => to_unsigned(848, 10), 1687 => to_unsigned(758, 10), 1688 => to_unsigned(189, 10), 1689 => to_unsigned(653, 10), 1690 => to_unsigned(684, 10), 1691 => to_unsigned(303, 10), 1692 => to_unsigned(3, 10), 1693 => to_unsigned(474, 10), 1694 => to_unsigned(674, 10), 1695 => to_unsigned(368, 10), 1696 => to_unsigned(371, 10), 1697 => to_unsigned(618, 10), 1698 => to_unsigned(684, 10), 1699 => to_unsigned(770, 10), 1700 => to_unsigned(77, 10), 1701 => to_unsigned(214, 10), 1702 => to_unsigned(780, 10), 1703 => to_unsigned(521, 10), 1704 => to_unsigned(592, 10), 1705 => to_unsigned(643, 10), 1706 => to_unsigned(192, 10), 1707 => to_unsigned(313, 10), 1708 => to_unsigned(524, 10), 1709 => to_unsigned(930, 10), 1710 => to_unsigned(316, 10), 1711 => to_unsigned(640, 10), 1712 => to_unsigned(21, 10), 1713 => to_unsigned(924, 10), 1714 => to_unsigned(503, 10), 1715 => to_unsigned(193, 10), 1716 => to_unsigned(410, 10), 1717 => to_unsigned(448, 10), 1718 => to_unsigned(725, 10), 1719 => to_unsigned(534, 10), 1720 => to_unsigned(115, 10), 1721 => to_unsigned(418, 10), 1722 => to_unsigned(1002, 10), 1723 => to_unsigned(481, 10), 1724 => to_unsigned(345, 10), 1725 => to_unsigned(839, 10), 1726 => to_unsigned(267, 10), 1727 => to_unsigned(237, 10), 1728 => to_unsigned(725, 10), 1729 => to_unsigned(1014, 10), 1730 => to_unsigned(598, 10), 1731 => to_unsigned(903, 10), 1732 => to_unsigned(417, 10), 1733 => to_unsigned(155, 10), 1734 => to_unsigned(953, 10), 1735 => to_unsigned(455, 10), 1736 => to_unsigned(486, 10), 1737 => to_unsigned(454, 10), 1738 => to_unsigned(488, 10), 1739 => to_unsigned(921, 10), 1740 => to_unsigned(259, 10), 1741 => to_unsigned(904, 10), 1742 => to_unsigned(429, 10), 1743 => to_unsigned(590, 10), 1744 => to_unsigned(978, 10), 1745 => to_unsigned(571, 10), 1746 => to_unsigned(839, 10), 1747 => to_unsigned(575, 10), 1748 => to_unsigned(658, 10), 1749 => to_unsigned(275, 10), 1750 => to_unsigned(422, 10), 1751 => to_unsigned(637, 10), 1752 => to_unsigned(414, 10), 1753 => to_unsigned(142, 10), 1754 => to_unsigned(247, 10), 1755 => to_unsigned(399, 10), 1756 => to_unsigned(324, 10), 1757 => to_unsigned(734, 10), 1758 => to_unsigned(738, 10), 1759 => to_unsigned(368, 10), 1760 => to_unsigned(139, 10), 1761 => to_unsigned(81, 10), 1762 => to_unsigned(367, 10), 1763 => to_unsigned(245, 10), 1764 => to_unsigned(585, 10), 1765 => to_unsigned(229, 10), 1766 => to_unsigned(417, 10), 1767 => to_unsigned(205, 10), 1768 => to_unsigned(421, 10), 1769 => to_unsigned(977, 10), 1770 => to_unsigned(164, 10), 1771 => to_unsigned(285, 10), 1772 => to_unsigned(50, 10), 1773 => to_unsigned(171, 10), 1774 => to_unsigned(510, 10), 1775 => to_unsigned(408, 10), 1776 => to_unsigned(886, 10), 1777 => to_unsigned(698, 10), 1778 => to_unsigned(487, 10), 1779 => to_unsigned(641, 10), 1780 => to_unsigned(499, 10), 1781 => to_unsigned(611, 10), 1782 => to_unsigned(358, 10), 1783 => to_unsigned(183, 10), 1784 => to_unsigned(700, 10), 1785 => to_unsigned(881, 10), 1786 => to_unsigned(511, 10), 1787 => to_unsigned(432, 10), 1788 => to_unsigned(427, 10), 1789 => to_unsigned(618, 10), 1790 => to_unsigned(818, 10), 1791 => to_unsigned(97, 10), 1792 => to_unsigned(802, 10), 1793 => to_unsigned(486, 10), 1794 => to_unsigned(863, 10), 1795 => to_unsigned(507, 10), 1796 => to_unsigned(710, 10), 1797 => to_unsigned(92, 10), 1798 => to_unsigned(172, 10), 1799 => to_unsigned(243, 10), 1800 => to_unsigned(333, 10), 1801 => to_unsigned(1012, 10), 1802 => to_unsigned(173, 10), 1803 => to_unsigned(104, 10), 1804 => to_unsigned(597, 10), 1805 => to_unsigned(953, 10), 1806 => to_unsigned(724, 10), 1807 => to_unsigned(594, 10), 1808 => to_unsigned(191, 10), 1809 => to_unsigned(343, 10), 1810 => to_unsigned(4, 10), 1811 => to_unsigned(603, 10), 1812 => to_unsigned(280, 10), 1813 => to_unsigned(780, 10), 1814 => to_unsigned(925, 10), 1815 => to_unsigned(988, 10), 1816 => to_unsigned(662, 10), 1817 => to_unsigned(969, 10), 1818 => to_unsigned(101, 10), 1819 => to_unsigned(402, 10), 1820 => to_unsigned(34, 10), 1821 => to_unsigned(527, 10), 1822 => to_unsigned(858, 10), 1823 => to_unsigned(11, 10), 1824 => to_unsigned(17, 10), 1825 => to_unsigned(668, 10), 1826 => to_unsigned(45, 10), 1827 => to_unsigned(403, 10), 1828 => to_unsigned(336, 10), 1829 => to_unsigned(658, 10), 1830 => to_unsigned(884, 10), 1831 => to_unsigned(499, 10), 1832 => to_unsigned(504, 10), 1833 => to_unsigned(472, 10), 1834 => to_unsigned(5, 10), 1835 => to_unsigned(186, 10), 1836 => to_unsigned(81, 10), 1837 => to_unsigned(58, 10), 1838 => to_unsigned(814, 10), 1839 => to_unsigned(125, 10), 1840 => to_unsigned(411, 10), 1841 => to_unsigned(592, 10), 1842 => to_unsigned(725, 10), 1843 => to_unsigned(94, 10), 1844 => to_unsigned(887, 10), 1845 => to_unsigned(828, 10), 1846 => to_unsigned(876, 10), 1847 => to_unsigned(897, 10), 1848 => to_unsigned(643, 10), 1849 => to_unsigned(232, 10), 1850 => to_unsigned(944, 10), 1851 => to_unsigned(191, 10), 1852 => to_unsigned(968, 10), 1853 => to_unsigned(348, 10), 1854 => to_unsigned(526, 10), 1855 => to_unsigned(750, 10), 1856 => to_unsigned(357, 10), 1857 => to_unsigned(336, 10), 1858 => to_unsigned(649, 10), 1859 => to_unsigned(182, 10), 1860 => to_unsigned(257, 10), 1861 => to_unsigned(469, 10), 1862 => to_unsigned(7, 10), 1863 => to_unsigned(776, 10), 1864 => to_unsigned(950, 10), 1865 => to_unsigned(537, 10), 1866 => to_unsigned(729, 10), 1867 => to_unsigned(930, 10), 1868 => to_unsigned(841, 10), 1869 => to_unsigned(315, 10), 1870 => to_unsigned(739, 10), 1871 => to_unsigned(280, 10), 1872 => to_unsigned(1006, 10), 1873 => to_unsigned(665, 10), 1874 => to_unsigned(61, 10), 1875 => to_unsigned(321, 10), 1876 => to_unsigned(902, 10), 1877 => to_unsigned(465, 10), 1878 => to_unsigned(740, 10), 1879 => to_unsigned(474, 10), 1880 => to_unsigned(998, 10), 1881 => to_unsigned(636, 10), 1882 => to_unsigned(816, 10), 1883 => to_unsigned(203, 10), 1884 => to_unsigned(454, 10), 1885 => to_unsigned(386, 10), 1886 => to_unsigned(523, 10), 1887 => to_unsigned(867, 10), 1888 => to_unsigned(533, 10), 1889 => to_unsigned(365, 10), 1890 => to_unsigned(588, 10), 1891 => to_unsigned(1009, 10), 1892 => to_unsigned(722, 10), 1893 => to_unsigned(940, 10), 1894 => to_unsigned(830, 10), 1895 => to_unsigned(215, 10), 1896 => to_unsigned(680, 10), 1897 => to_unsigned(709, 10), 1898 => to_unsigned(727, 10), 1899 => to_unsigned(970, 10), 1900 => to_unsigned(962, 10), 1901 => to_unsigned(813, 10), 1902 => to_unsigned(392, 10), 1903 => to_unsigned(826, 10), 1904 => to_unsigned(478, 10), 1905 => to_unsigned(207, 10), 1906 => to_unsigned(830, 10), 1907 => to_unsigned(363, 10), 1908 => to_unsigned(359, 10), 1909 => to_unsigned(182, 10), 1910 => to_unsigned(956, 10), 1911 => to_unsigned(728, 10), 1912 => to_unsigned(960, 10), 1913 => to_unsigned(307, 10), 1914 => to_unsigned(97, 10), 1915 => to_unsigned(213, 10), 1916 => to_unsigned(430, 10), 1917 => to_unsigned(48, 10), 1918 => to_unsigned(688, 10), 1919 => to_unsigned(1002, 10), 1920 => to_unsigned(245, 10), 1921 => to_unsigned(618, 10), 1922 => to_unsigned(679, 10), 1923 => to_unsigned(291, 10), 1924 => to_unsigned(349, 10), 1925 => to_unsigned(358, 10), 1926 => to_unsigned(492, 10), 1927 => to_unsigned(469, 10), 1928 => to_unsigned(665, 10), 1929 => to_unsigned(293, 10), 1930 => to_unsigned(780, 10), 1931 => to_unsigned(313, 10), 1932 => to_unsigned(277, 10), 1933 => to_unsigned(24, 10), 1934 => to_unsigned(791, 10), 1935 => to_unsigned(34, 10), 1936 => to_unsigned(757, 10), 1937 => to_unsigned(557, 10), 1938 => to_unsigned(863, 10), 1939 => to_unsigned(1004, 10), 1940 => to_unsigned(510, 10), 1941 => to_unsigned(1013, 10), 1942 => to_unsigned(324, 10), 1943 => to_unsigned(319, 10), 1944 => to_unsigned(1021, 10), 1945 => to_unsigned(737, 10), 1946 => to_unsigned(966, 10), 1947 => to_unsigned(750, 10), 1948 => to_unsigned(159, 10), 1949 => to_unsigned(666, 10), 1950 => to_unsigned(568, 10), 1951 => to_unsigned(764, 10), 1952 => to_unsigned(980, 10), 1953 => to_unsigned(992, 10), 1954 => to_unsigned(70, 10), 1955 => to_unsigned(899, 10), 1956 => to_unsigned(336, 10), 1957 => to_unsigned(946, 10), 1958 => to_unsigned(750, 10), 1959 => to_unsigned(632, 10), 1960 => to_unsigned(254, 10), 1961 => to_unsigned(382, 10), 1962 => to_unsigned(63, 10), 1963 => to_unsigned(248, 10), 1964 => to_unsigned(88, 10), 1965 => to_unsigned(646, 10), 1966 => to_unsigned(30, 10), 1967 => to_unsigned(897, 10), 1968 => to_unsigned(737, 10), 1969 => to_unsigned(1003, 10), 1970 => to_unsigned(383, 10), 1971 => to_unsigned(696, 10), 1972 => to_unsigned(6, 10), 1973 => to_unsigned(536, 10), 1974 => to_unsigned(160, 10), 1975 => to_unsigned(583, 10), 1976 => to_unsigned(106, 10), 1977 => to_unsigned(898, 10), 1978 => to_unsigned(970, 10), 1979 => to_unsigned(305, 10), 1980 => to_unsigned(833, 10), 1981 => to_unsigned(98, 10), 1982 => to_unsigned(66, 10), 1983 => to_unsigned(991, 10), 1984 => to_unsigned(670, 10), 1985 => to_unsigned(571, 10), 1986 => to_unsigned(290, 10), 1987 => to_unsigned(942, 10), 1988 => to_unsigned(861, 10), 1989 => to_unsigned(458, 10), 1990 => to_unsigned(61, 10), 1991 => to_unsigned(76, 10), 1992 => to_unsigned(921, 10), 1993 => to_unsigned(84, 10), 1994 => to_unsigned(950, 10), 1995 => to_unsigned(648, 10), 1996 => to_unsigned(712, 10), 1997 => to_unsigned(670, 10), 1998 => to_unsigned(507, 10), 1999 => to_unsigned(742, 10), 2000 => to_unsigned(585, 10), 2001 => to_unsigned(357, 10), 2002 => to_unsigned(504, 10), 2003 => to_unsigned(979, 10), 2004 => to_unsigned(15, 10), 2005 => to_unsigned(84, 10), 2006 => to_unsigned(847, 10), 2007 => to_unsigned(377, 10), 2008 => to_unsigned(782, 10), 2009 => to_unsigned(767, 10), 2010 => to_unsigned(242, 10), 2011 => to_unsigned(915, 10), 2012 => to_unsigned(1005, 10), 2013 => to_unsigned(626, 10), 2014 => to_unsigned(178, 10), 2015 => to_unsigned(24, 10), 2016 => to_unsigned(0, 10), 2017 => to_unsigned(1017, 10), 2018 => to_unsigned(87, 10), 2019 => to_unsigned(936, 10), 2020 => to_unsigned(761, 10), 2021 => to_unsigned(52, 10), 2022 => to_unsigned(154, 10), 2023 => to_unsigned(731, 10), 2024 => to_unsigned(682, 10), 2025 => to_unsigned(360, 10), 2026 => to_unsigned(867, 10), 2027 => to_unsigned(804, 10), 2028 => to_unsigned(455, 10), 2029 => to_unsigned(447, 10), 2030 => to_unsigned(203, 10), 2031 => to_unsigned(571, 10), 2032 => to_unsigned(996, 10), 2033 => to_unsigned(29, 10), 2034 => to_unsigned(442, 10), 2035 => to_unsigned(341, 10), 2036 => to_unsigned(912, 10), 2037 => to_unsigned(107, 10), 2038 => to_unsigned(70, 10), 2039 => to_unsigned(660, 10), 2040 => to_unsigned(754, 10), 2041 => to_unsigned(920, 10), 2042 => to_unsigned(291, 10), 2043 => to_unsigned(497, 10), 2044 => to_unsigned(80, 10), 2045 => to_unsigned(426, 10), 2046 => to_unsigned(664, 10), 2047 => to_unsigned(815, 10)),
            6 => (0 => to_unsigned(27, 10), 1 => to_unsigned(5, 10), 2 => to_unsigned(479, 10), 3 => to_unsigned(409, 10), 4 => to_unsigned(199, 10), 5 => to_unsigned(992, 10), 6 => to_unsigned(639, 10), 7 => to_unsigned(236, 10), 8 => to_unsigned(537, 10), 9 => to_unsigned(406, 10), 10 => to_unsigned(911, 10), 11 => to_unsigned(740, 10), 12 => to_unsigned(943, 10), 13 => to_unsigned(15, 10), 14 => to_unsigned(501, 10), 15 => to_unsigned(431, 10), 16 => to_unsigned(938, 10), 17 => to_unsigned(946, 10), 18 => to_unsigned(875, 10), 19 => to_unsigned(984, 10), 20 => to_unsigned(494, 10), 21 => to_unsigned(653, 10), 22 => to_unsigned(535, 10), 23 => to_unsigned(1001, 10), 24 => to_unsigned(953, 10), 25 => to_unsigned(49, 10), 26 => to_unsigned(1004, 10), 27 => to_unsigned(52, 10), 28 => to_unsigned(618, 10), 29 => to_unsigned(722, 10), 30 => to_unsigned(401, 10), 31 => to_unsigned(490, 10), 32 => to_unsigned(136, 10), 33 => to_unsigned(533, 10), 34 => to_unsigned(740, 10), 35 => to_unsigned(269, 10), 36 => to_unsigned(1008, 10), 37 => to_unsigned(615, 10), 38 => to_unsigned(739, 10), 39 => to_unsigned(80, 10), 40 => to_unsigned(549, 10), 41 => to_unsigned(696, 10), 42 => to_unsigned(461, 10), 43 => to_unsigned(161, 10), 44 => to_unsigned(843, 10), 45 => to_unsigned(832, 10), 46 => to_unsigned(910, 10), 47 => to_unsigned(43, 10), 48 => to_unsigned(920, 10), 49 => to_unsigned(91, 10), 50 => to_unsigned(788, 10), 51 => to_unsigned(798, 10), 52 => to_unsigned(782, 10), 53 => to_unsigned(684, 10), 54 => to_unsigned(94, 10), 55 => to_unsigned(1023, 10), 56 => to_unsigned(144, 10), 57 => to_unsigned(639, 10), 58 => to_unsigned(638, 10), 59 => to_unsigned(384, 10), 60 => to_unsigned(635, 10), 61 => to_unsigned(755, 10), 62 => to_unsigned(688, 10), 63 => to_unsigned(427, 10), 64 => to_unsigned(895, 10), 65 => to_unsigned(132, 10), 66 => to_unsigned(196, 10), 67 => to_unsigned(658, 10), 68 => to_unsigned(547, 10), 69 => to_unsigned(914, 10), 70 => to_unsigned(385, 10), 71 => to_unsigned(955, 10), 72 => to_unsigned(289, 10), 73 => to_unsigned(428, 10), 74 => to_unsigned(852, 10), 75 => to_unsigned(987, 10), 76 => to_unsigned(756, 10), 77 => to_unsigned(169, 10), 78 => to_unsigned(843, 10), 79 => to_unsigned(416, 10), 80 => to_unsigned(807, 10), 81 => to_unsigned(7, 10), 82 => to_unsigned(755, 10), 83 => to_unsigned(53, 10), 84 => to_unsigned(809, 10), 85 => to_unsigned(281, 10), 86 => to_unsigned(190, 10), 87 => to_unsigned(981, 10), 88 => to_unsigned(822, 10), 89 => to_unsigned(297, 10), 90 => to_unsigned(288, 10), 91 => to_unsigned(878, 10), 92 => to_unsigned(521, 10), 93 => to_unsigned(639, 10), 94 => to_unsigned(237, 10), 95 => to_unsigned(425, 10), 96 => to_unsigned(1002, 10), 97 => to_unsigned(583, 10), 98 => to_unsigned(313, 10), 99 => to_unsigned(305, 10), 100 => to_unsigned(108, 10), 101 => to_unsigned(719, 10), 102 => to_unsigned(800, 10), 103 => to_unsigned(823, 10), 104 => to_unsigned(88, 10), 105 => to_unsigned(782, 10), 106 => to_unsigned(980, 10), 107 => to_unsigned(792, 10), 108 => to_unsigned(598, 10), 109 => to_unsigned(738, 10), 110 => to_unsigned(566, 10), 111 => to_unsigned(607, 10), 112 => to_unsigned(770, 10), 113 => to_unsigned(498, 10), 114 => to_unsigned(562, 10), 115 => to_unsigned(568, 10), 116 => to_unsigned(651, 10), 117 => to_unsigned(563, 10), 118 => to_unsigned(663, 10), 119 => to_unsigned(811, 10), 120 => to_unsigned(827, 10), 121 => to_unsigned(184, 10), 122 => to_unsigned(387, 10), 123 => to_unsigned(967, 10), 124 => to_unsigned(521, 10), 125 => to_unsigned(138, 10), 126 => to_unsigned(990, 10), 127 => to_unsigned(257, 10), 128 => to_unsigned(404, 10), 129 => to_unsigned(210, 10), 130 => to_unsigned(638, 10), 131 => to_unsigned(301, 10), 132 => to_unsigned(293, 10), 133 => to_unsigned(23, 10), 134 => to_unsigned(446, 10), 135 => to_unsigned(248, 10), 136 => to_unsigned(940, 10), 137 => to_unsigned(616, 10), 138 => to_unsigned(441, 10), 139 => to_unsigned(346, 10), 140 => to_unsigned(556, 10), 141 => to_unsigned(381, 10), 142 => to_unsigned(837, 10), 143 => to_unsigned(429, 10), 144 => to_unsigned(660, 10), 145 => to_unsigned(49, 10), 146 => to_unsigned(326, 10), 147 => to_unsigned(307, 10), 148 => to_unsigned(197, 10), 149 => to_unsigned(141, 10), 150 => to_unsigned(387, 10), 151 => to_unsigned(96, 10), 152 => to_unsigned(53, 10), 153 => to_unsigned(284, 10), 154 => to_unsigned(817, 10), 155 => to_unsigned(511, 10), 156 => to_unsigned(152, 10), 157 => to_unsigned(823, 10), 158 => to_unsigned(444, 10), 159 => to_unsigned(318, 10), 160 => to_unsigned(315, 10), 161 => to_unsigned(557, 10), 162 => to_unsigned(795, 10), 163 => to_unsigned(485, 10), 164 => to_unsigned(826, 10), 165 => to_unsigned(642, 10), 166 => to_unsigned(557, 10), 167 => to_unsigned(225, 10), 168 => to_unsigned(361, 10), 169 => to_unsigned(892, 10), 170 => to_unsigned(531, 10), 171 => to_unsigned(976, 10), 172 => to_unsigned(717, 10), 173 => to_unsigned(976, 10), 174 => to_unsigned(33, 10), 175 => to_unsigned(55, 10), 176 => to_unsigned(563, 10), 177 => to_unsigned(301, 10), 178 => to_unsigned(630, 10), 179 => to_unsigned(759, 10), 180 => to_unsigned(134, 10), 181 => to_unsigned(860, 10), 182 => to_unsigned(576, 10), 183 => to_unsigned(926, 10), 184 => to_unsigned(693, 10), 185 => to_unsigned(685, 10), 186 => to_unsigned(235, 10), 187 => to_unsigned(200, 10), 188 => to_unsigned(708, 10), 189 => to_unsigned(634, 10), 190 => to_unsigned(201, 10), 191 => to_unsigned(915, 10), 192 => to_unsigned(199, 10), 193 => to_unsigned(549, 10), 194 => to_unsigned(725, 10), 195 => to_unsigned(309, 10), 196 => to_unsigned(999, 10), 197 => to_unsigned(402, 10), 198 => to_unsigned(35, 10), 199 => to_unsigned(858, 10), 200 => to_unsigned(169, 10), 201 => to_unsigned(64, 10), 202 => to_unsigned(642, 10), 203 => to_unsigned(863, 10), 204 => to_unsigned(868, 10), 205 => to_unsigned(161, 10), 206 => to_unsigned(454, 10), 207 => to_unsigned(361, 10), 208 => to_unsigned(589, 10), 209 => to_unsigned(673, 10), 210 => to_unsigned(319, 10), 211 => to_unsigned(280, 10), 212 => to_unsigned(742, 10), 213 => to_unsigned(226, 10), 214 => to_unsigned(212, 10), 215 => to_unsigned(144, 10), 216 => to_unsigned(398, 10), 217 => to_unsigned(910, 10), 218 => to_unsigned(724, 10), 219 => to_unsigned(524, 10), 220 => to_unsigned(660, 10), 221 => to_unsigned(272, 10), 222 => to_unsigned(500, 10), 223 => to_unsigned(109, 10), 224 => to_unsigned(348, 10), 225 => to_unsigned(766, 10), 226 => to_unsigned(398, 10), 227 => to_unsigned(677, 10), 228 => to_unsigned(917, 10), 229 => to_unsigned(777, 10), 230 => to_unsigned(60, 10), 231 => to_unsigned(108, 10), 232 => to_unsigned(484, 10), 233 => to_unsigned(22, 10), 234 => to_unsigned(726, 10), 235 => to_unsigned(134, 10), 236 => to_unsigned(495, 10), 237 => to_unsigned(857, 10), 238 => to_unsigned(582, 10), 239 => to_unsigned(144, 10), 240 => to_unsigned(969, 10), 241 => to_unsigned(312, 10), 242 => to_unsigned(629, 10), 243 => to_unsigned(612, 10), 244 => to_unsigned(581, 10), 245 => to_unsigned(292, 10), 246 => to_unsigned(545, 10), 247 => to_unsigned(1007, 10), 248 => to_unsigned(21, 10), 249 => to_unsigned(495, 10), 250 => to_unsigned(826, 10), 251 => to_unsigned(253, 10), 252 => to_unsigned(474, 10), 253 => to_unsigned(570, 10), 254 => to_unsigned(835, 10), 255 => to_unsigned(201, 10), 256 => to_unsigned(831, 10), 257 => to_unsigned(712, 10), 258 => to_unsigned(324, 10), 259 => to_unsigned(133, 10), 260 => to_unsigned(847, 10), 261 => to_unsigned(423, 10), 262 => to_unsigned(643, 10), 263 => to_unsigned(300, 10), 264 => to_unsigned(656, 10), 265 => to_unsigned(1011, 10), 266 => to_unsigned(123, 10), 267 => to_unsigned(674, 10), 268 => to_unsigned(543, 10), 269 => to_unsigned(246, 10), 270 => to_unsigned(329, 10), 271 => to_unsigned(431, 10), 272 => to_unsigned(420, 10), 273 => to_unsigned(414, 10), 274 => to_unsigned(649, 10), 275 => to_unsigned(422, 10), 276 => to_unsigned(672, 10), 277 => to_unsigned(514, 10), 278 => to_unsigned(953, 10), 279 => to_unsigned(523, 10), 280 => to_unsigned(750, 10), 281 => to_unsigned(822, 10), 282 => to_unsigned(243, 10), 283 => to_unsigned(344, 10), 284 => to_unsigned(216, 10), 285 => to_unsigned(955, 10), 286 => to_unsigned(183, 10), 287 => to_unsigned(937, 10), 288 => to_unsigned(753, 10), 289 => to_unsigned(667, 10), 290 => to_unsigned(77, 10), 291 => to_unsigned(171, 10), 292 => to_unsigned(383, 10), 293 => to_unsigned(107, 10), 294 => to_unsigned(175, 10), 295 => to_unsigned(452, 10), 296 => to_unsigned(274, 10), 297 => to_unsigned(453, 10), 298 => to_unsigned(262, 10), 299 => to_unsigned(76, 10), 300 => to_unsigned(356, 10), 301 => to_unsigned(43, 10), 302 => to_unsigned(714, 10), 303 => to_unsigned(559, 10), 304 => to_unsigned(747, 10), 305 => to_unsigned(1019, 10), 306 => to_unsigned(952, 10), 307 => to_unsigned(226, 10), 308 => to_unsigned(289, 10), 309 => to_unsigned(211, 10), 310 => to_unsigned(402, 10), 311 => to_unsigned(141, 10), 312 => to_unsigned(488, 10), 313 => to_unsigned(53, 10), 314 => to_unsigned(401, 10), 315 => to_unsigned(446, 10), 316 => to_unsigned(181, 10), 317 => to_unsigned(1017, 10), 318 => to_unsigned(486, 10), 319 => to_unsigned(129, 10), 320 => to_unsigned(202, 10), 321 => to_unsigned(651, 10), 322 => to_unsigned(887, 10), 323 => to_unsigned(784, 10), 324 => to_unsigned(687, 10), 325 => to_unsigned(789, 10), 326 => to_unsigned(403, 10), 327 => to_unsigned(830, 10), 328 => to_unsigned(607, 10), 329 => to_unsigned(818, 10), 330 => to_unsigned(874, 10), 331 => to_unsigned(585, 10), 332 => to_unsigned(677, 10), 333 => to_unsigned(429, 10), 334 => to_unsigned(854, 10), 335 => to_unsigned(851, 10), 336 => to_unsigned(640, 10), 337 => to_unsigned(262, 10), 338 => to_unsigned(258, 10), 339 => to_unsigned(627, 10), 340 => to_unsigned(426, 10), 341 => to_unsigned(119, 10), 342 => to_unsigned(48, 10), 343 => to_unsigned(321, 10), 344 => to_unsigned(841, 10), 345 => to_unsigned(177, 10), 346 => to_unsigned(599, 10), 347 => to_unsigned(599, 10), 348 => to_unsigned(101, 10), 349 => to_unsigned(539, 10), 350 => to_unsigned(92, 10), 351 => to_unsigned(190, 10), 352 => to_unsigned(251, 10), 353 => to_unsigned(357, 10), 354 => to_unsigned(933, 10), 355 => to_unsigned(999, 10), 356 => to_unsigned(809, 10), 357 => to_unsigned(751, 10), 358 => to_unsigned(706, 10), 359 => to_unsigned(855, 10), 360 => to_unsigned(947, 10), 361 => to_unsigned(994, 10), 362 => to_unsigned(576, 10), 363 => to_unsigned(868, 10), 364 => to_unsigned(963, 10), 365 => to_unsigned(1004, 10), 366 => to_unsigned(192, 10), 367 => to_unsigned(1015, 10), 368 => to_unsigned(537, 10), 369 => to_unsigned(27, 10), 370 => to_unsigned(100, 10), 371 => to_unsigned(176, 10), 372 => to_unsigned(321, 10), 373 => to_unsigned(760, 10), 374 => to_unsigned(519, 10), 375 => to_unsigned(865, 10), 376 => to_unsigned(668, 10), 377 => to_unsigned(676, 10), 378 => to_unsigned(749, 10), 379 => to_unsigned(422, 10), 380 => to_unsigned(616, 10), 381 => to_unsigned(573, 10), 382 => to_unsigned(37, 10), 383 => to_unsigned(99, 10), 384 => to_unsigned(465, 10), 385 => to_unsigned(187, 10), 386 => to_unsigned(90, 10), 387 => to_unsigned(565, 10), 388 => to_unsigned(562, 10), 389 => to_unsigned(319, 10), 390 => to_unsigned(1023, 10), 391 => to_unsigned(269, 10), 392 => to_unsigned(542, 10), 393 => to_unsigned(83, 10), 394 => to_unsigned(276, 10), 395 => to_unsigned(302, 10), 396 => to_unsigned(12, 10), 397 => to_unsigned(945, 10), 398 => to_unsigned(300, 10), 399 => to_unsigned(617, 10), 400 => to_unsigned(509, 10), 401 => to_unsigned(1011, 10), 402 => to_unsigned(188, 10), 403 => to_unsigned(970, 10), 404 => to_unsigned(813, 10), 405 => to_unsigned(246, 10), 406 => to_unsigned(301, 10), 407 => to_unsigned(532, 10), 408 => to_unsigned(318, 10), 409 => to_unsigned(603, 10), 410 => to_unsigned(407, 10), 411 => to_unsigned(162, 10), 412 => to_unsigned(162, 10), 413 => to_unsigned(977, 10), 414 => to_unsigned(574, 10), 415 => to_unsigned(486, 10), 416 => to_unsigned(348, 10), 417 => to_unsigned(64, 10), 418 => to_unsigned(444, 10), 419 => to_unsigned(826, 10), 420 => to_unsigned(1017, 10), 421 => to_unsigned(236, 10), 422 => to_unsigned(435, 10), 423 => to_unsigned(423, 10), 424 => to_unsigned(847, 10), 425 => to_unsigned(355, 10), 426 => to_unsigned(267, 10), 427 => to_unsigned(534, 10), 428 => to_unsigned(444, 10), 429 => to_unsigned(312, 10), 430 => to_unsigned(269, 10), 431 => to_unsigned(254, 10), 432 => to_unsigned(380, 10), 433 => to_unsigned(41, 10), 434 => to_unsigned(485, 10), 435 => to_unsigned(247, 10), 436 => to_unsigned(392, 10), 437 => to_unsigned(961, 10), 438 => to_unsigned(231, 10), 439 => to_unsigned(486, 10), 440 => to_unsigned(537, 10), 441 => to_unsigned(928, 10), 442 => to_unsigned(529, 10), 443 => to_unsigned(725, 10), 444 => to_unsigned(364, 10), 445 => to_unsigned(706, 10), 446 => to_unsigned(12, 10), 447 => to_unsigned(484, 10), 448 => to_unsigned(780, 10), 449 => to_unsigned(0, 10), 450 => to_unsigned(195, 10), 451 => to_unsigned(100, 10), 452 => to_unsigned(958, 10), 453 => to_unsigned(117, 10), 454 => to_unsigned(506, 10), 455 => to_unsigned(761, 10), 456 => to_unsigned(193, 10), 457 => to_unsigned(936, 10), 458 => to_unsigned(327, 10), 459 => to_unsigned(968, 10), 460 => to_unsigned(988, 10), 461 => to_unsigned(292, 10), 462 => to_unsigned(1023, 10), 463 => to_unsigned(481, 10), 464 => to_unsigned(645, 10), 465 => to_unsigned(605, 10), 466 => to_unsigned(966, 10), 467 => to_unsigned(669, 10), 468 => to_unsigned(981, 10), 469 => to_unsigned(637, 10), 470 => to_unsigned(488, 10), 471 => to_unsigned(142, 10), 472 => to_unsigned(182, 10), 473 => to_unsigned(34, 10), 474 => to_unsigned(940, 10), 475 => to_unsigned(687, 10), 476 => to_unsigned(672, 10), 477 => to_unsigned(731, 10), 478 => to_unsigned(140, 10), 479 => to_unsigned(223, 10), 480 => to_unsigned(575, 10), 481 => to_unsigned(463, 10), 482 => to_unsigned(75, 10), 483 => to_unsigned(507, 10), 484 => to_unsigned(236, 10), 485 => to_unsigned(177, 10), 486 => to_unsigned(369, 10), 487 => to_unsigned(416, 10), 488 => to_unsigned(833, 10), 489 => to_unsigned(334, 10), 490 => to_unsigned(809, 10), 491 => to_unsigned(481, 10), 492 => to_unsigned(219, 10), 493 => to_unsigned(827, 10), 494 => to_unsigned(597, 10), 495 => to_unsigned(251, 10), 496 => to_unsigned(353, 10), 497 => to_unsigned(234, 10), 498 => to_unsigned(938, 10), 499 => to_unsigned(997, 10), 500 => to_unsigned(513, 10), 501 => to_unsigned(19, 10), 502 => to_unsigned(395, 10), 503 => to_unsigned(644, 10), 504 => to_unsigned(777, 10), 505 => to_unsigned(795, 10), 506 => to_unsigned(847, 10), 507 => to_unsigned(705, 10), 508 => to_unsigned(867, 10), 509 => to_unsigned(0, 10), 510 => to_unsigned(336, 10), 511 => to_unsigned(584, 10), 512 => to_unsigned(273, 10), 513 => to_unsigned(742, 10), 514 => to_unsigned(724, 10), 515 => to_unsigned(763, 10), 516 => to_unsigned(50, 10), 517 => to_unsigned(256, 10), 518 => to_unsigned(279, 10), 519 => to_unsigned(557, 10), 520 => to_unsigned(337, 10), 521 => to_unsigned(625, 10), 522 => to_unsigned(200, 10), 523 => to_unsigned(9, 10), 524 => to_unsigned(347, 10), 525 => to_unsigned(841, 10), 526 => to_unsigned(370, 10), 527 => to_unsigned(178, 10), 528 => to_unsigned(934, 10), 529 => to_unsigned(287, 10), 530 => to_unsigned(391, 10), 531 => to_unsigned(1021, 10), 532 => to_unsigned(458, 10), 533 => to_unsigned(237, 10), 534 => to_unsigned(198, 10), 535 => to_unsigned(127, 10), 536 => to_unsigned(198, 10), 537 => to_unsigned(891, 10), 538 => to_unsigned(613, 10), 539 => to_unsigned(958, 10), 540 => to_unsigned(563, 10), 541 => to_unsigned(466, 10), 542 => to_unsigned(427, 10), 543 => to_unsigned(941, 10), 544 => to_unsigned(817, 10), 545 => to_unsigned(351, 10), 546 => to_unsigned(985, 10), 547 => to_unsigned(560, 10), 548 => to_unsigned(485, 10), 549 => to_unsigned(718, 10), 550 => to_unsigned(805, 10), 551 => to_unsigned(432, 10), 552 => to_unsigned(216, 10), 553 => to_unsigned(451, 10), 554 => to_unsigned(894, 10), 555 => to_unsigned(490, 10), 556 => to_unsigned(555, 10), 557 => to_unsigned(698, 10), 558 => to_unsigned(542, 10), 559 => to_unsigned(456, 10), 560 => to_unsigned(592, 10), 561 => to_unsigned(661, 10), 562 => to_unsigned(646, 10), 563 => to_unsigned(253, 10), 564 => to_unsigned(580, 10), 565 => to_unsigned(670, 10), 566 => to_unsigned(508, 10), 567 => to_unsigned(343, 10), 568 => to_unsigned(369, 10), 569 => to_unsigned(694, 10), 570 => to_unsigned(377, 10), 571 => to_unsigned(700, 10), 572 => to_unsigned(193, 10), 573 => to_unsigned(370, 10), 574 => to_unsigned(808, 10), 575 => to_unsigned(391, 10), 576 => to_unsigned(329, 10), 577 => to_unsigned(894, 10), 578 => to_unsigned(807, 10), 579 => to_unsigned(1010, 10), 580 => to_unsigned(237, 10), 581 => to_unsigned(904, 10), 582 => to_unsigned(284, 10), 583 => to_unsigned(528, 10), 584 => to_unsigned(532, 10), 585 => to_unsigned(260, 10), 586 => to_unsigned(419, 10), 587 => to_unsigned(827, 10), 588 => to_unsigned(506, 10), 589 => to_unsigned(488, 10), 590 => to_unsigned(233, 10), 591 => to_unsigned(463, 10), 592 => to_unsigned(622, 10), 593 => to_unsigned(355, 10), 594 => to_unsigned(929, 10), 595 => to_unsigned(332, 10), 596 => to_unsigned(206, 10), 597 => to_unsigned(178, 10), 598 => to_unsigned(866, 10), 599 => to_unsigned(707, 10), 600 => to_unsigned(389, 10), 601 => to_unsigned(927, 10), 602 => to_unsigned(983, 10), 603 => to_unsigned(50, 10), 604 => to_unsigned(1000, 10), 605 => to_unsigned(76, 10), 606 => to_unsigned(704, 10), 607 => to_unsigned(26, 10), 608 => to_unsigned(87, 10), 609 => to_unsigned(14, 10), 610 => to_unsigned(793, 10), 611 => to_unsigned(591, 10), 612 => to_unsigned(584, 10), 613 => to_unsigned(667, 10), 614 => to_unsigned(163, 10), 615 => to_unsigned(893, 10), 616 => to_unsigned(279, 10), 617 => to_unsigned(715, 10), 618 => to_unsigned(107, 10), 619 => to_unsigned(901, 10), 620 => to_unsigned(770, 10), 621 => to_unsigned(180, 10), 622 => to_unsigned(273, 10), 623 => to_unsigned(228, 10), 624 => to_unsigned(167, 10), 625 => to_unsigned(967, 10), 626 => to_unsigned(97, 10), 627 => to_unsigned(671, 10), 628 => to_unsigned(540, 10), 629 => to_unsigned(907, 10), 630 => to_unsigned(635, 10), 631 => to_unsigned(887, 10), 632 => to_unsigned(188, 10), 633 => to_unsigned(747, 10), 634 => to_unsigned(884, 10), 635 => to_unsigned(829, 10), 636 => to_unsigned(284, 10), 637 => to_unsigned(667, 10), 638 => to_unsigned(87, 10), 639 => to_unsigned(992, 10), 640 => to_unsigned(495, 10), 641 => to_unsigned(212, 10), 642 => to_unsigned(446, 10), 643 => to_unsigned(508, 10), 644 => to_unsigned(611, 10), 645 => to_unsigned(250, 10), 646 => to_unsigned(736, 10), 647 => to_unsigned(380, 10), 648 => to_unsigned(259, 10), 649 => to_unsigned(716, 10), 650 => to_unsigned(119, 10), 651 => to_unsigned(161, 10), 652 => to_unsigned(486, 10), 653 => to_unsigned(999, 10), 654 => to_unsigned(315, 10), 655 => to_unsigned(62, 10), 656 => to_unsigned(540, 10), 657 => to_unsigned(115, 10), 658 => to_unsigned(849, 10), 659 => to_unsigned(729, 10), 660 => to_unsigned(186, 10), 661 => to_unsigned(538, 10), 662 => to_unsigned(475, 10), 663 => to_unsigned(66, 10), 664 => to_unsigned(314, 10), 665 => to_unsigned(892, 10), 666 => to_unsigned(659, 10), 667 => to_unsigned(352, 10), 668 => to_unsigned(729, 10), 669 => to_unsigned(987, 10), 670 => to_unsigned(524, 10), 671 => to_unsigned(495, 10), 672 => to_unsigned(893, 10), 673 => to_unsigned(939, 10), 674 => to_unsigned(324, 10), 675 => to_unsigned(5, 10), 676 => to_unsigned(566, 10), 677 => to_unsigned(562, 10), 678 => to_unsigned(404, 10), 679 => to_unsigned(829, 10), 680 => to_unsigned(667, 10), 681 => to_unsigned(387, 10), 682 => to_unsigned(192, 10), 683 => to_unsigned(98, 10), 684 => to_unsigned(814, 10), 685 => to_unsigned(369, 10), 686 => to_unsigned(457, 10), 687 => to_unsigned(958, 10), 688 => to_unsigned(803, 10), 689 => to_unsigned(677, 10), 690 => to_unsigned(1, 10), 691 => to_unsigned(429, 10), 692 => to_unsigned(865, 10), 693 => to_unsigned(474, 10), 694 => to_unsigned(972, 10), 695 => to_unsigned(536, 10), 696 => to_unsigned(151, 10), 697 => to_unsigned(865, 10), 698 => to_unsigned(926, 10), 699 => to_unsigned(136, 10), 700 => to_unsigned(700, 10), 701 => to_unsigned(487, 10), 702 => to_unsigned(159, 10), 703 => to_unsigned(452, 10), 704 => to_unsigned(811, 10), 705 => to_unsigned(974, 10), 706 => to_unsigned(955, 10), 707 => to_unsigned(907, 10), 708 => to_unsigned(733, 10), 709 => to_unsigned(541, 10), 710 => to_unsigned(913, 10), 711 => to_unsigned(105, 10), 712 => to_unsigned(452, 10), 713 => to_unsigned(514, 10), 714 => to_unsigned(396, 10), 715 => to_unsigned(646, 10), 716 => to_unsigned(909, 10), 717 => to_unsigned(371, 10), 718 => to_unsigned(430, 10), 719 => to_unsigned(974, 10), 720 => to_unsigned(263, 10), 721 => to_unsigned(493, 10), 722 => to_unsigned(563, 10), 723 => to_unsigned(598, 10), 724 => to_unsigned(104, 10), 725 => to_unsigned(107, 10), 726 => to_unsigned(774, 10), 727 => to_unsigned(582, 10), 728 => to_unsigned(66, 10), 729 => to_unsigned(695, 10), 730 => to_unsigned(784, 10), 731 => to_unsigned(920, 10), 732 => to_unsigned(770, 10), 733 => to_unsigned(535, 10), 734 => to_unsigned(607, 10), 735 => to_unsigned(938, 10), 736 => to_unsigned(394, 10), 737 => to_unsigned(245, 10), 738 => to_unsigned(773, 10), 739 => to_unsigned(94, 10), 740 => to_unsigned(9, 10), 741 => to_unsigned(767, 10), 742 => to_unsigned(818, 10), 743 => to_unsigned(118, 10), 744 => to_unsigned(237, 10), 745 => to_unsigned(842, 10), 746 => to_unsigned(940, 10), 747 => to_unsigned(944, 10), 748 => to_unsigned(986, 10), 749 => to_unsigned(705, 10), 750 => to_unsigned(252, 10), 751 => to_unsigned(418, 10), 752 => to_unsigned(892, 10), 753 => to_unsigned(936, 10), 754 => to_unsigned(194, 10), 755 => to_unsigned(307, 10), 756 => to_unsigned(704, 10), 757 => to_unsigned(979, 10), 758 => to_unsigned(427, 10), 759 => to_unsigned(104, 10), 760 => to_unsigned(769, 10), 761 => to_unsigned(1006, 10), 762 => to_unsigned(73, 10), 763 => to_unsigned(659, 10), 764 => to_unsigned(108, 10), 765 => to_unsigned(198, 10), 766 => to_unsigned(884, 10), 767 => to_unsigned(714, 10), 768 => to_unsigned(481, 10), 769 => to_unsigned(598, 10), 770 => to_unsigned(672, 10), 771 => to_unsigned(332, 10), 772 => to_unsigned(898, 10), 773 => to_unsigned(583, 10), 774 => to_unsigned(327, 10), 775 => to_unsigned(328, 10), 776 => to_unsigned(1011, 10), 777 => to_unsigned(771, 10), 778 => to_unsigned(689, 10), 779 => to_unsigned(512, 10), 780 => to_unsigned(850, 10), 781 => to_unsigned(208, 10), 782 => to_unsigned(786, 10), 783 => to_unsigned(256, 10), 784 => to_unsigned(283, 10), 785 => to_unsigned(212, 10), 786 => to_unsigned(1018, 10), 787 => to_unsigned(970, 10), 788 => to_unsigned(877, 10), 789 => to_unsigned(52, 10), 790 => to_unsigned(963, 10), 791 => to_unsigned(485, 10), 792 => to_unsigned(531, 10), 793 => to_unsigned(339, 10), 794 => to_unsigned(338, 10), 795 => to_unsigned(496, 10), 796 => to_unsigned(837, 10), 797 => to_unsigned(498, 10), 798 => to_unsigned(642, 10), 799 => to_unsigned(533, 10), 800 => to_unsigned(103, 10), 801 => to_unsigned(802, 10), 802 => to_unsigned(810, 10), 803 => to_unsigned(537, 10), 804 => to_unsigned(866, 10), 805 => to_unsigned(219, 10), 806 => to_unsigned(488, 10), 807 => to_unsigned(254, 10), 808 => to_unsigned(575, 10), 809 => to_unsigned(550, 10), 810 => to_unsigned(665, 10), 811 => to_unsigned(875, 10), 812 => to_unsigned(205, 10), 813 => to_unsigned(302, 10), 814 => to_unsigned(95, 10), 815 => to_unsigned(561, 10), 816 => to_unsigned(843, 10), 817 => to_unsigned(755, 10), 818 => to_unsigned(333, 10), 819 => to_unsigned(318, 10), 820 => to_unsigned(551, 10), 821 => to_unsigned(642, 10), 822 => to_unsigned(643, 10), 823 => to_unsigned(28, 10), 824 => to_unsigned(473, 10), 825 => to_unsigned(774, 10), 826 => to_unsigned(453, 10), 827 => to_unsigned(269, 10), 828 => to_unsigned(562, 10), 829 => to_unsigned(864, 10), 830 => to_unsigned(563, 10), 831 => to_unsigned(427, 10), 832 => to_unsigned(725, 10), 833 => to_unsigned(850, 10), 834 => to_unsigned(92, 10), 835 => to_unsigned(41, 10), 836 => to_unsigned(406, 10), 837 => to_unsigned(891, 10), 838 => to_unsigned(205, 10), 839 => to_unsigned(44, 10), 840 => to_unsigned(549, 10), 841 => to_unsigned(534, 10), 842 => to_unsigned(576, 10), 843 => to_unsigned(546, 10), 844 => to_unsigned(581, 10), 845 => to_unsigned(511, 10), 846 => to_unsigned(104, 10), 847 => to_unsigned(495, 10), 848 => to_unsigned(28, 10), 849 => to_unsigned(531, 10), 850 => to_unsigned(661, 10), 851 => to_unsigned(624, 10), 852 => to_unsigned(811, 10), 853 => to_unsigned(517, 10), 854 => to_unsigned(958, 10), 855 => to_unsigned(16, 10), 856 => to_unsigned(795, 10), 857 => to_unsigned(808, 10), 858 => to_unsigned(979, 10), 859 => to_unsigned(474, 10), 860 => to_unsigned(203, 10), 861 => to_unsigned(792, 10), 862 => to_unsigned(173, 10), 863 => to_unsigned(383, 10), 864 => to_unsigned(876, 10), 865 => to_unsigned(174, 10), 866 => to_unsigned(47, 10), 867 => to_unsigned(751, 10), 868 => to_unsigned(633, 10), 869 => to_unsigned(628, 10), 870 => to_unsigned(870, 10), 871 => to_unsigned(265, 10), 872 => to_unsigned(363, 10), 873 => to_unsigned(613, 10), 874 => to_unsigned(80, 10), 875 => to_unsigned(776, 10), 876 => to_unsigned(408, 10), 877 => to_unsigned(616, 10), 878 => to_unsigned(250, 10), 879 => to_unsigned(59, 10), 880 => to_unsigned(385, 10), 881 => to_unsigned(716, 10), 882 => to_unsigned(153, 10), 883 => to_unsigned(323, 10), 884 => to_unsigned(541, 10), 885 => to_unsigned(686, 10), 886 => to_unsigned(204, 10), 887 => to_unsigned(713, 10), 888 => to_unsigned(307, 10), 889 => to_unsigned(466, 10), 890 => to_unsigned(923, 10), 891 => to_unsigned(817, 10), 892 => to_unsigned(569, 10), 893 => to_unsigned(952, 10), 894 => to_unsigned(728, 10), 895 => to_unsigned(605, 10), 896 => to_unsigned(310, 10), 897 => to_unsigned(309, 10), 898 => to_unsigned(399, 10), 899 => to_unsigned(606, 10), 900 => to_unsigned(734, 10), 901 => to_unsigned(530, 10), 902 => to_unsigned(436, 10), 903 => to_unsigned(717, 10), 904 => to_unsigned(619, 10), 905 => to_unsigned(14, 10), 906 => to_unsigned(136, 10), 907 => to_unsigned(466, 10), 908 => to_unsigned(516, 10), 909 => to_unsigned(333, 10), 910 => to_unsigned(502, 10), 911 => to_unsigned(730, 10), 912 => to_unsigned(569, 10), 913 => to_unsigned(94, 10), 914 => to_unsigned(912, 10), 915 => to_unsigned(782, 10), 916 => to_unsigned(377, 10), 917 => to_unsigned(938, 10), 918 => to_unsigned(225, 10), 919 => to_unsigned(424, 10), 920 => to_unsigned(278, 10), 921 => to_unsigned(97, 10), 922 => to_unsigned(314, 10), 923 => to_unsigned(766, 10), 924 => to_unsigned(109, 10), 925 => to_unsigned(807, 10), 926 => to_unsigned(28, 10), 927 => to_unsigned(863, 10), 928 => to_unsigned(749, 10), 929 => to_unsigned(53, 10), 930 => to_unsigned(508, 10), 931 => to_unsigned(393, 10), 932 => to_unsigned(867, 10), 933 => to_unsigned(484, 10), 934 => to_unsigned(182, 10), 935 => to_unsigned(832, 10), 936 => to_unsigned(169, 10), 937 => to_unsigned(920, 10), 938 => to_unsigned(611, 10), 939 => to_unsigned(808, 10), 940 => to_unsigned(262, 10), 941 => to_unsigned(657, 10), 942 => to_unsigned(225, 10), 943 => to_unsigned(876, 10), 944 => to_unsigned(376, 10), 945 => to_unsigned(61, 10), 946 => to_unsigned(459, 10), 947 => to_unsigned(571, 10), 948 => to_unsigned(231, 10), 949 => to_unsigned(568, 10), 950 => to_unsigned(708, 10), 951 => to_unsigned(825, 10), 952 => to_unsigned(117, 10), 953 => to_unsigned(373, 10), 954 => to_unsigned(169, 10), 955 => to_unsigned(476, 10), 956 => to_unsigned(825, 10), 957 => to_unsigned(864, 10), 958 => to_unsigned(785, 10), 959 => to_unsigned(9, 10), 960 => to_unsigned(561, 10), 961 => to_unsigned(412, 10), 962 => to_unsigned(936, 10), 963 => to_unsigned(723, 10), 964 => to_unsigned(621, 10), 965 => to_unsigned(329, 10), 966 => to_unsigned(651, 10), 967 => to_unsigned(282, 10), 968 => to_unsigned(492, 10), 969 => to_unsigned(150, 10), 970 => to_unsigned(1007, 10), 971 => to_unsigned(200, 10), 972 => to_unsigned(104, 10), 973 => to_unsigned(53, 10), 974 => to_unsigned(706, 10), 975 => to_unsigned(143, 10), 976 => to_unsigned(410, 10), 977 => to_unsigned(174, 10), 978 => to_unsigned(541, 10), 979 => to_unsigned(907, 10), 980 => to_unsigned(442, 10), 981 => to_unsigned(187, 10), 982 => to_unsigned(273, 10), 983 => to_unsigned(753, 10), 984 => to_unsigned(302, 10), 985 => to_unsigned(992, 10), 986 => to_unsigned(167, 10), 987 => to_unsigned(188, 10), 988 => to_unsigned(135, 10), 989 => to_unsigned(709, 10), 990 => to_unsigned(250, 10), 991 => to_unsigned(529, 10), 992 => to_unsigned(264, 10), 993 => to_unsigned(414, 10), 994 => to_unsigned(940, 10), 995 => to_unsigned(240, 10), 996 => to_unsigned(893, 10), 997 => to_unsigned(650, 10), 998 => to_unsigned(354, 10), 999 => to_unsigned(748, 10), 1000 => to_unsigned(914, 10), 1001 => to_unsigned(495, 10), 1002 => to_unsigned(61, 10), 1003 => to_unsigned(133, 10), 1004 => to_unsigned(29, 10), 1005 => to_unsigned(567, 10), 1006 => to_unsigned(641, 10), 1007 => to_unsigned(103, 10), 1008 => to_unsigned(932, 10), 1009 => to_unsigned(158, 10), 1010 => to_unsigned(78, 10), 1011 => to_unsigned(776, 10), 1012 => to_unsigned(232, 10), 1013 => to_unsigned(93, 10), 1014 => to_unsigned(130, 10), 1015 => to_unsigned(763, 10), 1016 => to_unsigned(152, 10), 1017 => to_unsigned(487, 10), 1018 => to_unsigned(298, 10), 1019 => to_unsigned(450, 10), 1020 => to_unsigned(194, 10), 1021 => to_unsigned(727, 10), 1022 => to_unsigned(614, 10), 1023 => to_unsigned(840, 10), 1024 => to_unsigned(124, 10), 1025 => to_unsigned(610, 10), 1026 => to_unsigned(329, 10), 1027 => to_unsigned(542, 10), 1028 => to_unsigned(514, 10), 1029 => to_unsigned(432, 10), 1030 => to_unsigned(913, 10), 1031 => to_unsigned(412, 10), 1032 => to_unsigned(403, 10), 1033 => to_unsigned(497, 10), 1034 => to_unsigned(525, 10), 1035 => to_unsigned(880, 10), 1036 => to_unsigned(68, 10), 1037 => to_unsigned(172, 10), 1038 => to_unsigned(650, 10), 1039 => to_unsigned(835, 10), 1040 => to_unsigned(973, 10), 1041 => to_unsigned(712, 10), 1042 => to_unsigned(9, 10), 1043 => to_unsigned(245, 10), 1044 => to_unsigned(138, 10), 1045 => to_unsigned(962, 10), 1046 => to_unsigned(375, 10), 1047 => to_unsigned(690, 10), 1048 => to_unsigned(564, 10), 1049 => to_unsigned(966, 10), 1050 => to_unsigned(948, 10), 1051 => to_unsigned(677, 10), 1052 => to_unsigned(576, 10), 1053 => to_unsigned(537, 10), 1054 => to_unsigned(925, 10), 1055 => to_unsigned(648, 10), 1056 => to_unsigned(230, 10), 1057 => to_unsigned(774, 10), 1058 => to_unsigned(334, 10), 1059 => to_unsigned(762, 10), 1060 => to_unsigned(305, 10), 1061 => to_unsigned(717, 10), 1062 => to_unsigned(937, 10), 1063 => to_unsigned(994, 10), 1064 => to_unsigned(208, 10), 1065 => to_unsigned(1006, 10), 1066 => to_unsigned(349, 10), 1067 => to_unsigned(193, 10), 1068 => to_unsigned(56, 10), 1069 => to_unsigned(774, 10), 1070 => to_unsigned(626, 10), 1071 => to_unsigned(760, 10), 1072 => to_unsigned(813, 10), 1073 => to_unsigned(679, 10), 1074 => to_unsigned(390, 10), 1075 => to_unsigned(729, 10), 1076 => to_unsigned(716, 10), 1077 => to_unsigned(444, 10), 1078 => to_unsigned(637, 10), 1079 => to_unsigned(193, 10), 1080 => to_unsigned(805, 10), 1081 => to_unsigned(830, 10), 1082 => to_unsigned(952, 10), 1083 => to_unsigned(861, 10), 1084 => to_unsigned(474, 10), 1085 => to_unsigned(187, 10), 1086 => to_unsigned(94, 10), 1087 => to_unsigned(205, 10), 1088 => to_unsigned(239, 10), 1089 => to_unsigned(527, 10), 1090 => to_unsigned(562, 10), 1091 => to_unsigned(829, 10), 1092 => to_unsigned(152, 10), 1093 => to_unsigned(288, 10), 1094 => to_unsigned(892, 10), 1095 => to_unsigned(685, 10), 1096 => to_unsigned(370, 10), 1097 => to_unsigned(838, 10), 1098 => to_unsigned(150, 10), 1099 => to_unsigned(274, 10), 1100 => to_unsigned(494, 10), 1101 => to_unsigned(336, 10), 1102 => to_unsigned(827, 10), 1103 => to_unsigned(316, 10), 1104 => to_unsigned(440, 10), 1105 => to_unsigned(10, 10), 1106 => to_unsigned(848, 10), 1107 => to_unsigned(44, 10), 1108 => to_unsigned(943, 10), 1109 => to_unsigned(703, 10), 1110 => to_unsigned(99, 10), 1111 => to_unsigned(890, 10), 1112 => to_unsigned(214, 10), 1113 => to_unsigned(841, 10), 1114 => to_unsigned(841, 10), 1115 => to_unsigned(447, 10), 1116 => to_unsigned(767, 10), 1117 => to_unsigned(823, 10), 1118 => to_unsigned(360, 10), 1119 => to_unsigned(1022, 10), 1120 => to_unsigned(819, 10), 1121 => to_unsigned(21, 10), 1122 => to_unsigned(889, 10), 1123 => to_unsigned(110, 10), 1124 => to_unsigned(926, 10), 1125 => to_unsigned(610, 10), 1126 => to_unsigned(728, 10), 1127 => to_unsigned(453, 10), 1128 => to_unsigned(550, 10), 1129 => to_unsigned(221, 10), 1130 => to_unsigned(299, 10), 1131 => to_unsigned(862, 10), 1132 => to_unsigned(329, 10), 1133 => to_unsigned(967, 10), 1134 => to_unsigned(139, 10), 1135 => to_unsigned(26, 10), 1136 => to_unsigned(612, 10), 1137 => to_unsigned(364, 10), 1138 => to_unsigned(119, 10), 1139 => to_unsigned(294, 10), 1140 => to_unsigned(758, 10), 1141 => to_unsigned(848, 10), 1142 => to_unsigned(769, 10), 1143 => to_unsigned(1010, 10), 1144 => to_unsigned(293, 10), 1145 => to_unsigned(579, 10), 1146 => to_unsigned(49, 10), 1147 => to_unsigned(618, 10), 1148 => to_unsigned(343, 10), 1149 => to_unsigned(931, 10), 1150 => to_unsigned(821, 10), 1151 => to_unsigned(617, 10), 1152 => to_unsigned(537, 10), 1153 => to_unsigned(780, 10), 1154 => to_unsigned(114, 10), 1155 => to_unsigned(349, 10), 1156 => to_unsigned(850, 10), 1157 => to_unsigned(967, 10), 1158 => to_unsigned(204, 10), 1159 => to_unsigned(736, 10), 1160 => to_unsigned(72, 10), 1161 => to_unsigned(219, 10), 1162 => to_unsigned(688, 10), 1163 => to_unsigned(506, 10), 1164 => to_unsigned(541, 10), 1165 => to_unsigned(528, 10), 1166 => to_unsigned(87, 10), 1167 => to_unsigned(498, 10), 1168 => to_unsigned(478, 10), 1169 => to_unsigned(631, 10), 1170 => to_unsigned(973, 10), 1171 => to_unsigned(49, 10), 1172 => to_unsigned(712, 10), 1173 => to_unsigned(869, 10), 1174 => to_unsigned(272, 10), 1175 => to_unsigned(370, 10), 1176 => to_unsigned(552, 10), 1177 => to_unsigned(990, 10), 1178 => to_unsigned(609, 10), 1179 => to_unsigned(419, 10), 1180 => to_unsigned(894, 10), 1181 => to_unsigned(491, 10), 1182 => to_unsigned(464, 10), 1183 => to_unsigned(619, 10), 1184 => to_unsigned(43, 10), 1185 => to_unsigned(91, 10), 1186 => to_unsigned(674, 10), 1187 => to_unsigned(140, 10), 1188 => to_unsigned(73, 10), 1189 => to_unsigned(357, 10), 1190 => to_unsigned(124, 10), 1191 => to_unsigned(459, 10), 1192 => to_unsigned(608, 10), 1193 => to_unsigned(386, 10), 1194 => to_unsigned(93, 10), 1195 => to_unsigned(934, 10), 1196 => to_unsigned(252, 10), 1197 => to_unsigned(410, 10), 1198 => to_unsigned(80, 10), 1199 => to_unsigned(455, 10), 1200 => to_unsigned(489, 10), 1201 => to_unsigned(602, 10), 1202 => to_unsigned(585, 10), 1203 => to_unsigned(587, 10), 1204 => to_unsigned(963, 10), 1205 => to_unsigned(583, 10), 1206 => to_unsigned(117, 10), 1207 => to_unsigned(35, 10), 1208 => to_unsigned(379, 10), 1209 => to_unsigned(385, 10), 1210 => to_unsigned(815, 10), 1211 => to_unsigned(220, 10), 1212 => to_unsigned(795, 10), 1213 => to_unsigned(595, 10), 1214 => to_unsigned(948, 10), 1215 => to_unsigned(1012, 10), 1216 => to_unsigned(411, 10), 1217 => to_unsigned(758, 10), 1218 => to_unsigned(520, 10), 1219 => to_unsigned(684, 10), 1220 => to_unsigned(781, 10), 1221 => to_unsigned(898, 10), 1222 => to_unsigned(313, 10), 1223 => to_unsigned(571, 10), 1224 => to_unsigned(821, 10), 1225 => to_unsigned(734, 10), 1226 => to_unsigned(555, 10), 1227 => to_unsigned(666, 10), 1228 => to_unsigned(504, 10), 1229 => to_unsigned(773, 10), 1230 => to_unsigned(871, 10), 1231 => to_unsigned(1008, 10), 1232 => to_unsigned(412, 10), 1233 => to_unsigned(281, 10), 1234 => to_unsigned(595, 10), 1235 => to_unsigned(451, 10), 1236 => to_unsigned(994, 10), 1237 => to_unsigned(229, 10), 1238 => to_unsigned(531, 10), 1239 => to_unsigned(205, 10), 1240 => to_unsigned(690, 10), 1241 => to_unsigned(446, 10), 1242 => to_unsigned(621, 10), 1243 => to_unsigned(404, 10), 1244 => to_unsigned(733, 10), 1245 => to_unsigned(341, 10), 1246 => to_unsigned(96, 10), 1247 => to_unsigned(1010, 10), 1248 => to_unsigned(896, 10), 1249 => to_unsigned(195, 10), 1250 => to_unsigned(409, 10), 1251 => to_unsigned(507, 10), 1252 => to_unsigned(376, 10), 1253 => to_unsigned(703, 10), 1254 => to_unsigned(592, 10), 1255 => to_unsigned(867, 10), 1256 => to_unsigned(305, 10), 1257 => to_unsigned(579, 10), 1258 => to_unsigned(707, 10), 1259 => to_unsigned(712, 10), 1260 => to_unsigned(373, 10), 1261 => to_unsigned(672, 10), 1262 => to_unsigned(618, 10), 1263 => to_unsigned(376, 10), 1264 => to_unsigned(975, 10), 1265 => to_unsigned(977, 10), 1266 => to_unsigned(983, 10), 1267 => to_unsigned(867, 10), 1268 => to_unsigned(184, 10), 1269 => to_unsigned(825, 10), 1270 => to_unsigned(145, 10), 1271 => to_unsigned(283, 10), 1272 => to_unsigned(831, 10), 1273 => to_unsigned(60, 10), 1274 => to_unsigned(378, 10), 1275 => to_unsigned(276, 10), 1276 => to_unsigned(572, 10), 1277 => to_unsigned(922, 10), 1278 => to_unsigned(821, 10), 1279 => to_unsigned(14, 10), 1280 => to_unsigned(414, 10), 1281 => to_unsigned(945, 10), 1282 => to_unsigned(235, 10), 1283 => to_unsigned(150, 10), 1284 => to_unsigned(1, 10), 1285 => to_unsigned(953, 10), 1286 => to_unsigned(29, 10), 1287 => to_unsigned(941, 10), 1288 => to_unsigned(118, 10), 1289 => to_unsigned(923, 10), 1290 => to_unsigned(485, 10), 1291 => to_unsigned(904, 10), 1292 => to_unsigned(157, 10), 1293 => to_unsigned(419, 10), 1294 => to_unsigned(893, 10), 1295 => to_unsigned(426, 10), 1296 => to_unsigned(986, 10), 1297 => to_unsigned(42, 10), 1298 => to_unsigned(41, 10), 1299 => to_unsigned(592, 10), 1300 => to_unsigned(343, 10), 1301 => to_unsigned(911, 10), 1302 => to_unsigned(825, 10), 1303 => to_unsigned(79, 10), 1304 => to_unsigned(935, 10), 1305 => to_unsigned(916, 10), 1306 => to_unsigned(875, 10), 1307 => to_unsigned(367, 10), 1308 => to_unsigned(425, 10), 1309 => to_unsigned(428, 10), 1310 => to_unsigned(74, 10), 1311 => to_unsigned(886, 10), 1312 => to_unsigned(331, 10), 1313 => to_unsigned(636, 10), 1314 => to_unsigned(491, 10), 1315 => to_unsigned(654, 10), 1316 => to_unsigned(217, 10), 1317 => to_unsigned(971, 10), 1318 => to_unsigned(77, 10), 1319 => to_unsigned(953, 10), 1320 => to_unsigned(691, 10), 1321 => to_unsigned(516, 10), 1322 => to_unsigned(610, 10), 1323 => to_unsigned(831, 10), 1324 => to_unsigned(322, 10), 1325 => to_unsigned(533, 10), 1326 => to_unsigned(300, 10), 1327 => to_unsigned(52, 10), 1328 => to_unsigned(110, 10), 1329 => to_unsigned(850, 10), 1330 => to_unsigned(243, 10), 1331 => to_unsigned(923, 10), 1332 => to_unsigned(521, 10), 1333 => to_unsigned(305, 10), 1334 => to_unsigned(981, 10), 1335 => to_unsigned(1020, 10), 1336 => to_unsigned(697, 10), 1337 => to_unsigned(863, 10), 1338 => to_unsigned(19, 10), 1339 => to_unsigned(605, 10), 1340 => to_unsigned(445, 10), 1341 => to_unsigned(377, 10), 1342 => to_unsigned(213, 10), 1343 => to_unsigned(855, 10), 1344 => to_unsigned(166, 10), 1345 => to_unsigned(978, 10), 1346 => to_unsigned(141, 10), 1347 => to_unsigned(712, 10), 1348 => to_unsigned(706, 10), 1349 => to_unsigned(32, 10), 1350 => to_unsigned(900, 10), 1351 => to_unsigned(517, 10), 1352 => to_unsigned(295, 10), 1353 => to_unsigned(810, 10), 1354 => to_unsigned(847, 10), 1355 => to_unsigned(50, 10), 1356 => to_unsigned(623, 10), 1357 => to_unsigned(354, 10), 1358 => to_unsigned(586, 10), 1359 => to_unsigned(106, 10), 1360 => to_unsigned(130, 10), 1361 => to_unsigned(112, 10), 1362 => to_unsigned(153, 10), 1363 => to_unsigned(418, 10), 1364 => to_unsigned(578, 10), 1365 => to_unsigned(139, 10), 1366 => to_unsigned(675, 10), 1367 => to_unsigned(747, 10), 1368 => to_unsigned(576, 10), 1369 => to_unsigned(187, 10), 1370 => to_unsigned(488, 10), 1371 => to_unsigned(871, 10), 1372 => to_unsigned(816, 10), 1373 => to_unsigned(68, 10), 1374 => to_unsigned(673, 10), 1375 => to_unsigned(73, 10), 1376 => to_unsigned(518, 10), 1377 => to_unsigned(249, 10), 1378 => to_unsigned(922, 10), 1379 => to_unsigned(131, 10), 1380 => to_unsigned(767, 10), 1381 => to_unsigned(162, 10), 1382 => to_unsigned(844, 10), 1383 => to_unsigned(160, 10), 1384 => to_unsigned(931, 10), 1385 => to_unsigned(547, 10), 1386 => to_unsigned(253, 10), 1387 => to_unsigned(536, 10), 1388 => to_unsigned(435, 10), 1389 => to_unsigned(121, 10), 1390 => to_unsigned(914, 10), 1391 => to_unsigned(99, 10), 1392 => to_unsigned(425, 10), 1393 => to_unsigned(615, 10), 1394 => to_unsigned(166, 10), 1395 => to_unsigned(663, 10), 1396 => to_unsigned(348, 10), 1397 => to_unsigned(696, 10), 1398 => to_unsigned(1019, 10), 1399 => to_unsigned(1018, 10), 1400 => to_unsigned(266, 10), 1401 => to_unsigned(166, 10), 1402 => to_unsigned(756, 10), 1403 => to_unsigned(326, 10), 1404 => to_unsigned(629, 10), 1405 => to_unsigned(49, 10), 1406 => to_unsigned(835, 10), 1407 => to_unsigned(344, 10), 1408 => to_unsigned(779, 10), 1409 => to_unsigned(796, 10), 1410 => to_unsigned(180, 10), 1411 => to_unsigned(349, 10), 1412 => to_unsigned(94, 10), 1413 => to_unsigned(445, 10), 1414 => to_unsigned(780, 10), 1415 => to_unsigned(307, 10), 1416 => to_unsigned(62, 10), 1417 => to_unsigned(919, 10), 1418 => to_unsigned(294, 10), 1419 => to_unsigned(509, 10), 1420 => to_unsigned(799, 10), 1421 => to_unsigned(769, 10), 1422 => to_unsigned(488, 10), 1423 => to_unsigned(504, 10), 1424 => to_unsigned(315, 10), 1425 => to_unsigned(444, 10), 1426 => to_unsigned(375, 10), 1427 => to_unsigned(693, 10), 1428 => to_unsigned(115, 10), 1429 => to_unsigned(93, 10), 1430 => to_unsigned(944, 10), 1431 => to_unsigned(679, 10), 1432 => to_unsigned(362, 10), 1433 => to_unsigned(377, 10), 1434 => to_unsigned(739, 10), 1435 => to_unsigned(489, 10), 1436 => to_unsigned(805, 10), 1437 => to_unsigned(93, 10), 1438 => to_unsigned(25, 10), 1439 => to_unsigned(933, 10), 1440 => to_unsigned(117, 10), 1441 => to_unsigned(430, 10), 1442 => to_unsigned(308, 10), 1443 => to_unsigned(860, 10), 1444 => to_unsigned(602, 10), 1445 => to_unsigned(931, 10), 1446 => to_unsigned(294, 10), 1447 => to_unsigned(115, 10), 1448 => to_unsigned(256, 10), 1449 => to_unsigned(922, 10), 1450 => to_unsigned(366, 10), 1451 => to_unsigned(623, 10), 1452 => to_unsigned(110, 10), 1453 => to_unsigned(437, 10), 1454 => to_unsigned(324, 10), 1455 => to_unsigned(703, 10), 1456 => to_unsigned(798, 10), 1457 => to_unsigned(908, 10), 1458 => to_unsigned(202, 10), 1459 => to_unsigned(832, 10), 1460 => to_unsigned(446, 10), 1461 => to_unsigned(941, 10), 1462 => to_unsigned(275, 10), 1463 => to_unsigned(433, 10), 1464 => to_unsigned(952, 10), 1465 => to_unsigned(640, 10), 1466 => to_unsigned(703, 10), 1467 => to_unsigned(373, 10), 1468 => to_unsigned(480, 10), 1469 => to_unsigned(403, 10), 1470 => to_unsigned(806, 10), 1471 => to_unsigned(309, 10), 1472 => to_unsigned(615, 10), 1473 => to_unsigned(919, 10), 1474 => to_unsigned(430, 10), 1475 => to_unsigned(634, 10), 1476 => to_unsigned(848, 10), 1477 => to_unsigned(756, 10), 1478 => to_unsigned(754, 10), 1479 => to_unsigned(112, 10), 1480 => to_unsigned(602, 10), 1481 => to_unsigned(445, 10), 1482 => to_unsigned(72, 10), 1483 => to_unsigned(924, 10), 1484 => to_unsigned(534, 10), 1485 => to_unsigned(935, 10), 1486 => to_unsigned(226, 10), 1487 => to_unsigned(310, 10), 1488 => to_unsigned(335, 10), 1489 => to_unsigned(71, 10), 1490 => to_unsigned(577, 10), 1491 => to_unsigned(796, 10), 1492 => to_unsigned(826, 10), 1493 => to_unsigned(322, 10), 1494 => to_unsigned(392, 10), 1495 => to_unsigned(889, 10), 1496 => to_unsigned(303, 10), 1497 => to_unsigned(667, 10), 1498 => to_unsigned(403, 10), 1499 => to_unsigned(228, 10), 1500 => to_unsigned(466, 10), 1501 => to_unsigned(934, 10), 1502 => to_unsigned(419, 10), 1503 => to_unsigned(495, 10), 1504 => to_unsigned(496, 10), 1505 => to_unsigned(938, 10), 1506 => to_unsigned(248, 10), 1507 => to_unsigned(127, 10), 1508 => to_unsigned(7, 10), 1509 => to_unsigned(1014, 10), 1510 => to_unsigned(624, 10), 1511 => to_unsigned(621, 10), 1512 => to_unsigned(880, 10), 1513 => to_unsigned(740, 10), 1514 => to_unsigned(822, 10), 1515 => to_unsigned(765, 10), 1516 => to_unsigned(95, 10), 1517 => to_unsigned(516, 10), 1518 => to_unsigned(453, 10), 1519 => to_unsigned(391, 10), 1520 => to_unsigned(279, 10), 1521 => to_unsigned(948, 10), 1522 => to_unsigned(220, 10), 1523 => to_unsigned(313, 10), 1524 => to_unsigned(578, 10), 1525 => to_unsigned(772, 10), 1526 => to_unsigned(324, 10), 1527 => to_unsigned(474, 10), 1528 => to_unsigned(525, 10), 1529 => to_unsigned(538, 10), 1530 => to_unsigned(236, 10), 1531 => to_unsigned(641, 10), 1532 => to_unsigned(534, 10), 1533 => to_unsigned(54, 10), 1534 => to_unsigned(762, 10), 1535 => to_unsigned(46, 10), 1536 => to_unsigned(584, 10), 1537 => to_unsigned(5, 10), 1538 => to_unsigned(196, 10), 1539 => to_unsigned(765, 10), 1540 => to_unsigned(652, 10), 1541 => to_unsigned(402, 10), 1542 => to_unsigned(494, 10), 1543 => to_unsigned(737, 10), 1544 => to_unsigned(130, 10), 1545 => to_unsigned(349, 10), 1546 => to_unsigned(447, 10), 1547 => to_unsigned(303, 10), 1548 => to_unsigned(345, 10), 1549 => to_unsigned(674, 10), 1550 => to_unsigned(442, 10), 1551 => to_unsigned(149, 10), 1552 => to_unsigned(892, 10), 1553 => to_unsigned(968, 10), 1554 => to_unsigned(529, 10), 1555 => to_unsigned(922, 10), 1556 => to_unsigned(760, 10), 1557 => to_unsigned(228, 10), 1558 => to_unsigned(107, 10), 1559 => to_unsigned(157, 10), 1560 => to_unsigned(380, 10), 1561 => to_unsigned(459, 10), 1562 => to_unsigned(224, 10), 1563 => to_unsigned(87, 10), 1564 => to_unsigned(83, 10), 1565 => to_unsigned(768, 10), 1566 => to_unsigned(789, 10), 1567 => to_unsigned(668, 10), 1568 => to_unsigned(289, 10), 1569 => to_unsigned(182, 10), 1570 => to_unsigned(1003, 10), 1571 => to_unsigned(765, 10), 1572 => to_unsigned(146, 10), 1573 => to_unsigned(256, 10), 1574 => to_unsigned(38, 10), 1575 => to_unsigned(850, 10), 1576 => to_unsigned(946, 10), 1577 => to_unsigned(986, 10), 1578 => to_unsigned(845, 10), 1579 => to_unsigned(691, 10), 1580 => to_unsigned(707, 10), 1581 => to_unsigned(769, 10), 1582 => to_unsigned(167, 10), 1583 => to_unsigned(919, 10), 1584 => to_unsigned(172, 10), 1585 => to_unsigned(415, 10), 1586 => to_unsigned(7, 10), 1587 => to_unsigned(158, 10), 1588 => to_unsigned(374, 10), 1589 => to_unsigned(540, 10), 1590 => to_unsigned(182, 10), 1591 => to_unsigned(304, 10), 1592 => to_unsigned(776, 10), 1593 => to_unsigned(218, 10), 1594 => to_unsigned(133, 10), 1595 => to_unsigned(773, 10), 1596 => to_unsigned(245, 10), 1597 => to_unsigned(35, 10), 1598 => to_unsigned(410, 10), 1599 => to_unsigned(115, 10), 1600 => to_unsigned(52, 10), 1601 => to_unsigned(869, 10), 1602 => to_unsigned(80, 10), 1603 => to_unsigned(441, 10), 1604 => to_unsigned(885, 10), 1605 => to_unsigned(995, 10), 1606 => to_unsigned(744, 10), 1607 => to_unsigned(524, 10), 1608 => to_unsigned(924, 10), 1609 => to_unsigned(773, 10), 1610 => to_unsigned(770, 10), 1611 => to_unsigned(50, 10), 1612 => to_unsigned(852, 10), 1613 => to_unsigned(184, 10), 1614 => to_unsigned(254, 10), 1615 => to_unsigned(782, 10), 1616 => to_unsigned(81, 10), 1617 => to_unsigned(90, 10), 1618 => to_unsigned(628, 10), 1619 => to_unsigned(260, 10), 1620 => to_unsigned(174, 10), 1621 => to_unsigned(520, 10), 1622 => to_unsigned(200, 10), 1623 => to_unsigned(531, 10), 1624 => to_unsigned(15, 10), 1625 => to_unsigned(147, 10), 1626 => to_unsigned(370, 10), 1627 => to_unsigned(630, 10), 1628 => to_unsigned(530, 10), 1629 => to_unsigned(857, 10), 1630 => to_unsigned(485, 10), 1631 => to_unsigned(462, 10), 1632 => to_unsigned(664, 10), 1633 => to_unsigned(446, 10), 1634 => to_unsigned(252, 10), 1635 => to_unsigned(453, 10), 1636 => to_unsigned(562, 10), 1637 => to_unsigned(9, 10), 1638 => to_unsigned(27, 10), 1639 => to_unsigned(90, 10), 1640 => to_unsigned(719, 10), 1641 => to_unsigned(803, 10), 1642 => to_unsigned(717, 10), 1643 => to_unsigned(778, 10), 1644 => to_unsigned(523, 10), 1645 => to_unsigned(99, 10), 1646 => to_unsigned(14, 10), 1647 => to_unsigned(242, 10), 1648 => to_unsigned(448, 10), 1649 => to_unsigned(457, 10), 1650 => to_unsigned(434, 10), 1651 => to_unsigned(959, 10), 1652 => to_unsigned(365, 10), 1653 => to_unsigned(577, 10), 1654 => to_unsigned(196, 10), 1655 => to_unsigned(985, 10), 1656 => to_unsigned(667, 10), 1657 => to_unsigned(309, 10), 1658 => to_unsigned(309, 10), 1659 => to_unsigned(1020, 10), 1660 => to_unsigned(100, 10), 1661 => to_unsigned(211, 10), 1662 => to_unsigned(781, 10), 1663 => to_unsigned(472, 10), 1664 => to_unsigned(1009, 10), 1665 => to_unsigned(175, 10), 1666 => to_unsigned(660, 10), 1667 => to_unsigned(384, 10), 1668 => to_unsigned(864, 10), 1669 => to_unsigned(40, 10), 1670 => to_unsigned(478, 10), 1671 => to_unsigned(866, 10), 1672 => to_unsigned(165, 10), 1673 => to_unsigned(740, 10), 1674 => to_unsigned(489, 10), 1675 => to_unsigned(110, 10), 1676 => to_unsigned(548, 10), 1677 => to_unsigned(482, 10), 1678 => to_unsigned(144, 10), 1679 => to_unsigned(612, 10), 1680 => to_unsigned(311, 10), 1681 => to_unsigned(901, 10), 1682 => to_unsigned(345, 10), 1683 => to_unsigned(504, 10), 1684 => to_unsigned(625, 10), 1685 => to_unsigned(769, 10), 1686 => to_unsigned(1023, 10), 1687 => to_unsigned(790, 10), 1688 => to_unsigned(855, 10), 1689 => to_unsigned(204, 10), 1690 => to_unsigned(840, 10), 1691 => to_unsigned(313, 10), 1692 => to_unsigned(420, 10), 1693 => to_unsigned(470, 10), 1694 => to_unsigned(490, 10), 1695 => to_unsigned(433, 10), 1696 => to_unsigned(156, 10), 1697 => to_unsigned(390, 10), 1698 => to_unsigned(142, 10), 1699 => to_unsigned(559, 10), 1700 => to_unsigned(499, 10), 1701 => to_unsigned(220, 10), 1702 => to_unsigned(117, 10), 1703 => to_unsigned(13, 10), 1704 => to_unsigned(482, 10), 1705 => to_unsigned(319, 10), 1706 => to_unsigned(501, 10), 1707 => to_unsigned(326, 10), 1708 => to_unsigned(478, 10), 1709 => to_unsigned(778, 10), 1710 => to_unsigned(640, 10), 1711 => to_unsigned(824, 10), 1712 => to_unsigned(647, 10), 1713 => to_unsigned(770, 10), 1714 => to_unsigned(282, 10), 1715 => to_unsigned(592, 10), 1716 => to_unsigned(869, 10), 1717 => to_unsigned(194, 10), 1718 => to_unsigned(941, 10), 1719 => to_unsigned(95, 10), 1720 => to_unsigned(372, 10), 1721 => to_unsigned(131, 10), 1722 => to_unsigned(741, 10), 1723 => to_unsigned(449, 10), 1724 => to_unsigned(879, 10), 1725 => to_unsigned(37, 10), 1726 => to_unsigned(122, 10), 1727 => to_unsigned(525, 10), 1728 => to_unsigned(700, 10), 1729 => to_unsigned(447, 10), 1730 => to_unsigned(197, 10), 1731 => to_unsigned(274, 10), 1732 => to_unsigned(815, 10), 1733 => to_unsigned(545, 10), 1734 => to_unsigned(215, 10), 1735 => to_unsigned(500, 10), 1736 => to_unsigned(930, 10), 1737 => to_unsigned(490, 10), 1738 => to_unsigned(65, 10), 1739 => to_unsigned(370, 10), 1740 => to_unsigned(47, 10), 1741 => to_unsigned(350, 10), 1742 => to_unsigned(148, 10), 1743 => to_unsigned(152, 10), 1744 => to_unsigned(527, 10), 1745 => to_unsigned(448, 10), 1746 => to_unsigned(403, 10), 1747 => to_unsigned(644, 10), 1748 => to_unsigned(776, 10), 1749 => to_unsigned(258, 10), 1750 => to_unsigned(667, 10), 1751 => to_unsigned(129, 10), 1752 => to_unsigned(60, 10), 1753 => to_unsigned(383, 10), 1754 => to_unsigned(291, 10), 1755 => to_unsigned(156, 10), 1756 => to_unsigned(1004, 10), 1757 => to_unsigned(39, 10), 1758 => to_unsigned(784, 10), 1759 => to_unsigned(551, 10), 1760 => to_unsigned(117, 10), 1761 => to_unsigned(938, 10), 1762 => to_unsigned(305, 10), 1763 => to_unsigned(773, 10), 1764 => to_unsigned(65, 10), 1765 => to_unsigned(1002, 10), 1766 => to_unsigned(605, 10), 1767 => to_unsigned(591, 10), 1768 => to_unsigned(498, 10), 1769 => to_unsigned(349, 10), 1770 => to_unsigned(218, 10), 1771 => to_unsigned(354, 10), 1772 => to_unsigned(500, 10), 1773 => to_unsigned(754, 10), 1774 => to_unsigned(725, 10), 1775 => to_unsigned(84, 10), 1776 => to_unsigned(567, 10), 1777 => to_unsigned(346, 10), 1778 => to_unsigned(357, 10), 1779 => to_unsigned(664, 10), 1780 => to_unsigned(29, 10), 1781 => to_unsigned(305, 10), 1782 => to_unsigned(188, 10), 1783 => to_unsigned(948, 10), 1784 => to_unsigned(606, 10), 1785 => to_unsigned(767, 10), 1786 => to_unsigned(208, 10), 1787 => to_unsigned(204, 10), 1788 => to_unsigned(619, 10), 1789 => to_unsigned(587, 10), 1790 => to_unsigned(146, 10), 1791 => to_unsigned(830, 10), 1792 => to_unsigned(486, 10), 1793 => to_unsigned(738, 10), 1794 => to_unsigned(659, 10), 1795 => to_unsigned(585, 10), 1796 => to_unsigned(544, 10), 1797 => to_unsigned(12, 10), 1798 => to_unsigned(555, 10), 1799 => to_unsigned(18, 10), 1800 => to_unsigned(323, 10), 1801 => to_unsigned(875, 10), 1802 => to_unsigned(174, 10), 1803 => to_unsigned(628, 10), 1804 => to_unsigned(516, 10), 1805 => to_unsigned(779, 10), 1806 => to_unsigned(644, 10), 1807 => to_unsigned(663, 10), 1808 => to_unsigned(697, 10), 1809 => to_unsigned(217, 10), 1810 => to_unsigned(557, 10), 1811 => to_unsigned(26, 10), 1812 => to_unsigned(449, 10), 1813 => to_unsigned(390, 10), 1814 => to_unsigned(725, 10), 1815 => to_unsigned(724, 10), 1816 => to_unsigned(990, 10), 1817 => to_unsigned(483, 10), 1818 => to_unsigned(350, 10), 1819 => to_unsigned(520, 10), 1820 => to_unsigned(824, 10), 1821 => to_unsigned(267, 10), 1822 => to_unsigned(189, 10), 1823 => to_unsigned(420, 10), 1824 => to_unsigned(626, 10), 1825 => to_unsigned(702, 10), 1826 => to_unsigned(130, 10), 1827 => to_unsigned(619, 10), 1828 => to_unsigned(719, 10), 1829 => to_unsigned(750, 10), 1830 => to_unsigned(329, 10), 1831 => to_unsigned(584, 10), 1832 => to_unsigned(963, 10), 1833 => to_unsigned(852, 10), 1834 => to_unsigned(665, 10), 1835 => to_unsigned(53, 10), 1836 => to_unsigned(384, 10), 1837 => to_unsigned(329, 10), 1838 => to_unsigned(562, 10), 1839 => to_unsigned(644, 10), 1840 => to_unsigned(70, 10), 1841 => to_unsigned(586, 10), 1842 => to_unsigned(650, 10), 1843 => to_unsigned(800, 10), 1844 => to_unsigned(114, 10), 1845 => to_unsigned(423, 10), 1846 => to_unsigned(382, 10), 1847 => to_unsigned(259, 10), 1848 => to_unsigned(981, 10), 1849 => to_unsigned(636, 10), 1850 => to_unsigned(211, 10), 1851 => to_unsigned(653, 10), 1852 => to_unsigned(789, 10), 1853 => to_unsigned(628, 10), 1854 => to_unsigned(776, 10), 1855 => to_unsigned(252, 10), 1856 => to_unsigned(970, 10), 1857 => to_unsigned(314, 10), 1858 => to_unsigned(298, 10), 1859 => to_unsigned(541, 10), 1860 => to_unsigned(605, 10), 1861 => to_unsigned(231, 10), 1862 => to_unsigned(514, 10), 1863 => to_unsigned(512, 10), 1864 => to_unsigned(652, 10), 1865 => to_unsigned(698, 10), 1866 => to_unsigned(524, 10), 1867 => to_unsigned(970, 10), 1868 => to_unsigned(528, 10), 1869 => to_unsigned(742, 10), 1870 => to_unsigned(857, 10), 1871 => to_unsigned(923, 10), 1872 => to_unsigned(733, 10), 1873 => to_unsigned(321, 10), 1874 => to_unsigned(496, 10), 1875 => to_unsigned(5, 10), 1876 => to_unsigned(604, 10), 1877 => to_unsigned(530, 10), 1878 => to_unsigned(348, 10), 1879 => to_unsigned(450, 10), 1880 => to_unsigned(141, 10), 1881 => to_unsigned(722, 10), 1882 => to_unsigned(707, 10), 1883 => to_unsigned(716, 10), 1884 => to_unsigned(533, 10), 1885 => to_unsigned(137, 10), 1886 => to_unsigned(477, 10), 1887 => to_unsigned(124, 10), 1888 => to_unsigned(727, 10), 1889 => to_unsigned(801, 10), 1890 => to_unsigned(328, 10), 1891 => to_unsigned(7, 10), 1892 => to_unsigned(349, 10), 1893 => to_unsigned(137, 10), 1894 => to_unsigned(243, 10), 1895 => to_unsigned(688, 10), 1896 => to_unsigned(243, 10), 1897 => to_unsigned(415, 10), 1898 => to_unsigned(795, 10), 1899 => to_unsigned(761, 10), 1900 => to_unsigned(878, 10), 1901 => to_unsigned(36, 10), 1902 => to_unsigned(830, 10), 1903 => to_unsigned(689, 10), 1904 => to_unsigned(843, 10), 1905 => to_unsigned(878, 10), 1906 => to_unsigned(710, 10), 1907 => to_unsigned(925, 10), 1908 => to_unsigned(637, 10), 1909 => to_unsigned(265, 10), 1910 => to_unsigned(14, 10), 1911 => to_unsigned(948, 10), 1912 => to_unsigned(94, 10), 1913 => to_unsigned(630, 10), 1914 => to_unsigned(699, 10), 1915 => to_unsigned(857, 10), 1916 => to_unsigned(4, 10), 1917 => to_unsigned(62, 10), 1918 => to_unsigned(25, 10), 1919 => to_unsigned(62, 10), 1920 => to_unsigned(209, 10), 1921 => to_unsigned(787, 10), 1922 => to_unsigned(623, 10), 1923 => to_unsigned(43, 10), 1924 => to_unsigned(1005, 10), 1925 => to_unsigned(528, 10), 1926 => to_unsigned(480, 10), 1927 => to_unsigned(254, 10), 1928 => to_unsigned(663, 10), 1929 => to_unsigned(929, 10), 1930 => to_unsigned(616, 10), 1931 => to_unsigned(151, 10), 1932 => to_unsigned(127, 10), 1933 => to_unsigned(658, 10), 1934 => to_unsigned(189, 10), 1935 => to_unsigned(109, 10), 1936 => to_unsigned(109, 10), 1937 => to_unsigned(737, 10), 1938 => to_unsigned(676, 10), 1939 => to_unsigned(977, 10), 1940 => to_unsigned(132, 10), 1941 => to_unsigned(153, 10), 1942 => to_unsigned(340, 10), 1943 => to_unsigned(440, 10), 1944 => to_unsigned(486, 10), 1945 => to_unsigned(359, 10), 1946 => to_unsigned(1022, 10), 1947 => to_unsigned(968, 10), 1948 => to_unsigned(1022, 10), 1949 => to_unsigned(419, 10), 1950 => to_unsigned(653, 10), 1951 => to_unsigned(629, 10), 1952 => to_unsigned(422, 10), 1953 => to_unsigned(791, 10), 1954 => to_unsigned(282, 10), 1955 => to_unsigned(456, 10), 1956 => to_unsigned(467, 10), 1957 => to_unsigned(480, 10), 1958 => to_unsigned(757, 10), 1959 => to_unsigned(772, 10), 1960 => to_unsigned(545, 10), 1961 => to_unsigned(471, 10), 1962 => to_unsigned(433, 10), 1963 => to_unsigned(935, 10), 1964 => to_unsigned(724, 10), 1965 => to_unsigned(400, 10), 1966 => to_unsigned(1000, 10), 1967 => to_unsigned(671, 10), 1968 => to_unsigned(505, 10), 1969 => to_unsigned(823, 10), 1970 => to_unsigned(15, 10), 1971 => to_unsigned(227, 10), 1972 => to_unsigned(377, 10), 1973 => to_unsigned(900, 10), 1974 => to_unsigned(654, 10), 1975 => to_unsigned(68, 10), 1976 => to_unsigned(819, 10), 1977 => to_unsigned(672, 10), 1978 => to_unsigned(387, 10), 1979 => to_unsigned(935, 10), 1980 => to_unsigned(181, 10), 1981 => to_unsigned(455, 10), 1982 => to_unsigned(566, 10), 1983 => to_unsigned(920, 10), 1984 => to_unsigned(827, 10), 1985 => to_unsigned(1018, 10), 1986 => to_unsigned(818, 10), 1987 => to_unsigned(993, 10), 1988 => to_unsigned(681, 10), 1989 => to_unsigned(587, 10), 1990 => to_unsigned(978, 10), 1991 => to_unsigned(710, 10), 1992 => to_unsigned(4, 10), 1993 => to_unsigned(61, 10), 1994 => to_unsigned(343, 10), 1995 => to_unsigned(215, 10), 1996 => to_unsigned(156, 10), 1997 => to_unsigned(518, 10), 1998 => to_unsigned(658, 10), 1999 => to_unsigned(450, 10), 2000 => to_unsigned(822, 10), 2001 => to_unsigned(2, 10), 2002 => to_unsigned(868, 10), 2003 => to_unsigned(115, 10), 2004 => to_unsigned(425, 10), 2005 => to_unsigned(764, 10), 2006 => to_unsigned(100, 10), 2007 => to_unsigned(95, 10), 2008 => to_unsigned(448, 10), 2009 => to_unsigned(381, 10), 2010 => to_unsigned(732, 10), 2011 => to_unsigned(42, 10), 2012 => to_unsigned(265, 10), 2013 => to_unsigned(813, 10), 2014 => to_unsigned(595, 10), 2015 => to_unsigned(431, 10), 2016 => to_unsigned(649, 10), 2017 => to_unsigned(238, 10), 2018 => to_unsigned(15, 10), 2019 => to_unsigned(125, 10), 2020 => to_unsigned(615, 10), 2021 => to_unsigned(828, 10), 2022 => to_unsigned(392, 10), 2023 => to_unsigned(121, 10), 2024 => to_unsigned(741, 10), 2025 => to_unsigned(957, 10), 2026 => to_unsigned(743, 10), 2027 => to_unsigned(100, 10), 2028 => to_unsigned(260, 10), 2029 => to_unsigned(780, 10), 2030 => to_unsigned(48, 10), 2031 => to_unsigned(542, 10), 2032 => to_unsigned(758, 10), 2033 => to_unsigned(446, 10), 2034 => to_unsigned(300, 10), 2035 => to_unsigned(833, 10), 2036 => to_unsigned(712, 10), 2037 => to_unsigned(497, 10), 2038 => to_unsigned(955, 10), 2039 => to_unsigned(106, 10), 2040 => to_unsigned(859, 10), 2041 => to_unsigned(506, 10), 2042 => to_unsigned(923, 10), 2043 => to_unsigned(544, 10), 2044 => to_unsigned(983, 10), 2045 => to_unsigned(562, 10), 2046 => to_unsigned(872, 10), 2047 => to_unsigned(741, 10)),
            7 => (0 => to_unsigned(143, 10), 1 => to_unsigned(142, 10), 2 => to_unsigned(82, 10), 3 => to_unsigned(977, 10), 4 => to_unsigned(480, 10), 5 => to_unsigned(675, 10), 6 => to_unsigned(557, 10), 7 => to_unsigned(286, 10), 8 => to_unsigned(381, 10), 9 => to_unsigned(985, 10), 10 => to_unsigned(11, 10), 11 => to_unsigned(583, 10), 12 => to_unsigned(833, 10), 13 => to_unsigned(229, 10), 14 => to_unsigned(466, 10), 15 => to_unsigned(562, 10), 16 => to_unsigned(432, 10), 17 => to_unsigned(612, 10), 18 => to_unsigned(934, 10), 19 => to_unsigned(731, 10), 20 => to_unsigned(507, 10), 21 => to_unsigned(160, 10), 22 => to_unsigned(155, 10), 23 => to_unsigned(27, 10), 24 => to_unsigned(230, 10), 25 => to_unsigned(878, 10), 26 => to_unsigned(634, 10), 27 => to_unsigned(979, 10), 28 => to_unsigned(644, 10), 29 => to_unsigned(239, 10), 30 => to_unsigned(440, 10), 31 => to_unsigned(812, 10), 32 => to_unsigned(872, 10), 33 => to_unsigned(76, 10), 34 => to_unsigned(551, 10), 35 => to_unsigned(1006, 10), 36 => to_unsigned(616, 10), 37 => to_unsigned(227, 10), 38 => to_unsigned(771, 10), 39 => to_unsigned(4, 10), 40 => to_unsigned(748, 10), 41 => to_unsigned(39, 10), 42 => to_unsigned(557, 10), 43 => to_unsigned(815, 10), 44 => to_unsigned(1014, 10), 45 => to_unsigned(499, 10), 46 => to_unsigned(666, 10), 47 => to_unsigned(195, 10), 48 => to_unsigned(535, 10), 49 => to_unsigned(892, 10), 50 => to_unsigned(995, 10), 51 => to_unsigned(979, 10), 52 => to_unsigned(30, 10), 53 => to_unsigned(701, 10), 54 => to_unsigned(111, 10), 55 => to_unsigned(646, 10), 56 => to_unsigned(493, 10), 57 => to_unsigned(171, 10), 58 => to_unsigned(736, 10), 59 => to_unsigned(735, 10), 60 => to_unsigned(832, 10), 61 => to_unsigned(317, 10), 62 => to_unsigned(305, 10), 63 => to_unsigned(892, 10), 64 => to_unsigned(741, 10), 65 => to_unsigned(433, 10), 66 => to_unsigned(183, 10), 67 => to_unsigned(261, 10), 68 => to_unsigned(314, 10), 69 => to_unsigned(906, 10), 70 => to_unsigned(273, 10), 71 => to_unsigned(249, 10), 72 => to_unsigned(185, 10), 73 => to_unsigned(122, 10), 74 => to_unsigned(873, 10), 75 => to_unsigned(450, 10), 76 => to_unsigned(832, 10), 77 => to_unsigned(514, 10), 78 => to_unsigned(152, 10), 79 => to_unsigned(1004, 10), 80 => to_unsigned(856, 10), 81 => to_unsigned(489, 10), 82 => to_unsigned(311, 10), 83 => to_unsigned(682, 10), 84 => to_unsigned(952, 10), 85 => to_unsigned(503, 10), 86 => to_unsigned(218, 10), 87 => to_unsigned(755, 10), 88 => to_unsigned(736, 10), 89 => to_unsigned(878, 10), 90 => to_unsigned(953, 10), 91 => to_unsigned(442, 10), 92 => to_unsigned(664, 10), 93 => to_unsigned(849, 10), 94 => to_unsigned(430, 10), 95 => to_unsigned(1013, 10), 96 => to_unsigned(530, 10), 97 => to_unsigned(143, 10), 98 => to_unsigned(323, 10), 99 => to_unsigned(709, 10), 100 => to_unsigned(458, 10), 101 => to_unsigned(867, 10), 102 => to_unsigned(225, 10), 103 => to_unsigned(642, 10), 104 => to_unsigned(881, 10), 105 => to_unsigned(160, 10), 106 => to_unsigned(473, 10), 107 => to_unsigned(245, 10), 108 => to_unsigned(536, 10), 109 => to_unsigned(900, 10), 110 => to_unsigned(517, 10), 111 => to_unsigned(769, 10), 112 => to_unsigned(733, 10), 113 => to_unsigned(1018, 10), 114 => to_unsigned(987, 10), 115 => to_unsigned(181, 10), 116 => to_unsigned(265, 10), 117 => to_unsigned(737, 10), 118 => to_unsigned(976, 10), 119 => to_unsigned(914, 10), 120 => to_unsigned(215, 10), 121 => to_unsigned(639, 10), 122 => to_unsigned(17, 10), 123 => to_unsigned(208, 10), 124 => to_unsigned(890, 10), 125 => to_unsigned(613, 10), 126 => to_unsigned(558, 10), 127 => to_unsigned(64, 10), 128 => to_unsigned(397, 10), 129 => to_unsigned(538, 10), 130 => to_unsigned(315, 10), 131 => to_unsigned(565, 10), 132 => to_unsigned(970, 10), 133 => to_unsigned(554, 10), 134 => to_unsigned(861, 10), 135 => to_unsigned(281, 10), 136 => to_unsigned(65, 10), 137 => to_unsigned(167, 10), 138 => to_unsigned(251, 10), 139 => to_unsigned(198, 10), 140 => to_unsigned(157, 10), 141 => to_unsigned(687, 10), 142 => to_unsigned(411, 10), 143 => to_unsigned(741, 10), 144 => to_unsigned(832, 10), 145 => to_unsigned(409, 10), 146 => to_unsigned(860, 10), 147 => to_unsigned(343, 10), 148 => to_unsigned(130, 10), 149 => to_unsigned(898, 10), 150 => to_unsigned(975, 10), 151 => to_unsigned(283, 10), 152 => to_unsigned(326, 10), 153 => to_unsigned(737, 10), 154 => to_unsigned(73, 10), 155 => to_unsigned(169, 10), 156 => to_unsigned(192, 10), 157 => to_unsigned(347, 10), 158 => to_unsigned(1013, 10), 159 => to_unsigned(669, 10), 160 => to_unsigned(77, 10), 161 => to_unsigned(1013, 10), 162 => to_unsigned(209, 10), 163 => to_unsigned(922, 10), 164 => to_unsigned(576, 10), 165 => to_unsigned(130, 10), 166 => to_unsigned(1004, 10), 167 => to_unsigned(412, 10), 168 => to_unsigned(886, 10), 169 => to_unsigned(320, 10), 170 => to_unsigned(647, 10), 171 => to_unsigned(468, 10), 172 => to_unsigned(896, 10), 173 => to_unsigned(21, 10), 174 => to_unsigned(1004, 10), 175 => to_unsigned(162, 10), 176 => to_unsigned(573, 10), 177 => to_unsigned(252, 10), 178 => to_unsigned(670, 10), 179 => to_unsigned(730, 10), 180 => to_unsigned(147, 10), 181 => to_unsigned(821, 10), 182 => to_unsigned(933, 10), 183 => to_unsigned(808, 10), 184 => to_unsigned(1011, 10), 185 => to_unsigned(849, 10), 186 => to_unsigned(236, 10), 187 => to_unsigned(964, 10), 188 => to_unsigned(784, 10), 189 => to_unsigned(146, 10), 190 => to_unsigned(440, 10), 191 => to_unsigned(654, 10), 192 => to_unsigned(979, 10), 193 => to_unsigned(890, 10), 194 => to_unsigned(367, 10), 195 => to_unsigned(759, 10), 196 => to_unsigned(845, 10), 197 => to_unsigned(520, 10), 198 => to_unsigned(167, 10), 199 => to_unsigned(622, 10), 200 => to_unsigned(240, 10), 201 => to_unsigned(138, 10), 202 => to_unsigned(165, 10), 203 => to_unsigned(599, 10), 204 => to_unsigned(983, 10), 205 => to_unsigned(494, 10), 206 => to_unsigned(185, 10), 207 => to_unsigned(189, 10), 208 => to_unsigned(507, 10), 209 => to_unsigned(175, 10), 210 => to_unsigned(383, 10), 211 => to_unsigned(65, 10), 212 => to_unsigned(598, 10), 213 => to_unsigned(732, 10), 214 => to_unsigned(605, 10), 215 => to_unsigned(521, 10), 216 => to_unsigned(336, 10), 217 => to_unsigned(910, 10), 218 => to_unsigned(475, 10), 219 => to_unsigned(252, 10), 220 => to_unsigned(767, 10), 221 => to_unsigned(183, 10), 222 => to_unsigned(574, 10), 223 => to_unsigned(716, 10), 224 => to_unsigned(706, 10), 225 => to_unsigned(976, 10), 226 => to_unsigned(1001, 10), 227 => to_unsigned(424, 10), 228 => to_unsigned(807, 10), 229 => to_unsigned(641, 10), 230 => to_unsigned(303, 10), 231 => to_unsigned(745, 10), 232 => to_unsigned(858, 10), 233 => to_unsigned(939, 10), 234 => to_unsigned(171, 10), 235 => to_unsigned(24, 10), 236 => to_unsigned(925, 10), 237 => to_unsigned(145, 10), 238 => to_unsigned(639, 10), 239 => to_unsigned(684, 10), 240 => to_unsigned(484, 10), 241 => to_unsigned(231, 10), 242 => to_unsigned(690, 10), 243 => to_unsigned(805, 10), 244 => to_unsigned(467, 10), 245 => to_unsigned(955, 10), 246 => to_unsigned(1001, 10), 247 => to_unsigned(438, 10), 248 => to_unsigned(121, 10), 249 => to_unsigned(445, 10), 250 => to_unsigned(910, 10), 251 => to_unsigned(38, 10), 252 => to_unsigned(826, 10), 253 => to_unsigned(621, 10), 254 => to_unsigned(393, 10), 255 => to_unsigned(472, 10), 256 => to_unsigned(523, 10), 257 => to_unsigned(272, 10), 258 => to_unsigned(751, 10), 259 => to_unsigned(597, 10), 260 => to_unsigned(126, 10), 261 => to_unsigned(939, 10), 262 => to_unsigned(781, 10), 263 => to_unsigned(406, 10), 264 => to_unsigned(1013, 10), 265 => to_unsigned(536, 10), 266 => to_unsigned(907, 10), 267 => to_unsigned(339, 10), 268 => to_unsigned(349, 10), 269 => to_unsigned(175, 10), 270 => to_unsigned(604, 10), 271 => to_unsigned(380, 10), 272 => to_unsigned(344, 10), 273 => to_unsigned(564, 10), 274 => to_unsigned(182, 10), 275 => to_unsigned(98, 10), 276 => to_unsigned(74, 10), 277 => to_unsigned(414, 10), 278 => to_unsigned(1003, 10), 279 => to_unsigned(753, 10), 280 => to_unsigned(434, 10), 281 => to_unsigned(323, 10), 282 => to_unsigned(169, 10), 283 => to_unsigned(243, 10), 284 => to_unsigned(329, 10), 285 => to_unsigned(306, 10), 286 => to_unsigned(870, 10), 287 => to_unsigned(503, 10), 288 => to_unsigned(566, 10), 289 => to_unsigned(603, 10), 290 => to_unsigned(894, 10), 291 => to_unsigned(4, 10), 292 => to_unsigned(129, 10), 293 => to_unsigned(990, 10), 294 => to_unsigned(764, 10), 295 => to_unsigned(113, 10), 296 => to_unsigned(859, 10), 297 => to_unsigned(791, 10), 298 => to_unsigned(729, 10), 299 => to_unsigned(658, 10), 300 => to_unsigned(922, 10), 301 => to_unsigned(340, 10), 302 => to_unsigned(325, 10), 303 => to_unsigned(952, 10), 304 => to_unsigned(268, 10), 305 => to_unsigned(236, 10), 306 => to_unsigned(15, 10), 307 => to_unsigned(782, 10), 308 => to_unsigned(414, 10), 309 => to_unsigned(968, 10), 310 => to_unsigned(307, 10), 311 => to_unsigned(737, 10), 312 => to_unsigned(410, 10), 313 => to_unsigned(110, 10), 314 => to_unsigned(204, 10), 315 => to_unsigned(371, 10), 316 => to_unsigned(559, 10), 317 => to_unsigned(66, 10), 318 => to_unsigned(112, 10), 319 => to_unsigned(915, 10), 320 => to_unsigned(132, 10), 321 => to_unsigned(699, 10), 322 => to_unsigned(654, 10), 323 => to_unsigned(698, 10), 324 => to_unsigned(291, 10), 325 => to_unsigned(263, 10), 326 => to_unsigned(397, 10), 327 => to_unsigned(448, 10), 328 => to_unsigned(295, 10), 329 => to_unsigned(903, 10), 330 => to_unsigned(249, 10), 331 => to_unsigned(483, 10), 332 => to_unsigned(319, 10), 333 => to_unsigned(386, 10), 334 => to_unsigned(743, 10), 335 => to_unsigned(138, 10), 336 => to_unsigned(854, 10), 337 => to_unsigned(925, 10), 338 => to_unsigned(430, 10), 339 => to_unsigned(136, 10), 340 => to_unsigned(675, 10), 341 => to_unsigned(824, 10), 342 => to_unsigned(640, 10), 343 => to_unsigned(95, 10), 344 => to_unsigned(198, 10), 345 => to_unsigned(869, 10), 346 => to_unsigned(16, 10), 347 => to_unsigned(713, 10), 348 => to_unsigned(191, 10), 349 => to_unsigned(862, 10), 350 => to_unsigned(21, 10), 351 => to_unsigned(446, 10), 352 => to_unsigned(348, 10), 353 => to_unsigned(33, 10), 354 => to_unsigned(1021, 10), 355 => to_unsigned(263, 10), 356 => to_unsigned(398, 10), 357 => to_unsigned(1008, 10), 358 => to_unsigned(694, 10), 359 => to_unsigned(143, 10), 360 => to_unsigned(410, 10), 361 => to_unsigned(523, 10), 362 => to_unsigned(718, 10), 363 => to_unsigned(553, 10), 364 => to_unsigned(312, 10), 365 => to_unsigned(720, 10), 366 => to_unsigned(1002, 10), 367 => to_unsigned(280, 10), 368 => to_unsigned(386, 10), 369 => to_unsigned(959, 10), 370 => to_unsigned(863, 10), 371 => to_unsigned(1010, 10), 372 => to_unsigned(836, 10), 373 => to_unsigned(43, 10), 374 => to_unsigned(115, 10), 375 => to_unsigned(649, 10), 376 => to_unsigned(857, 10), 377 => to_unsigned(187, 10), 378 => to_unsigned(289, 10), 379 => to_unsigned(283, 10), 380 => to_unsigned(778, 10), 381 => to_unsigned(370, 10), 382 => to_unsigned(487, 10), 383 => to_unsigned(222, 10), 384 => to_unsigned(1006, 10), 385 => to_unsigned(829, 10), 386 => to_unsigned(154, 10), 387 => to_unsigned(800, 10), 388 => to_unsigned(81, 10), 389 => to_unsigned(669, 10), 390 => to_unsigned(748, 10), 391 => to_unsigned(477, 10), 392 => to_unsigned(440, 10), 393 => to_unsigned(294, 10), 394 => to_unsigned(232, 10), 395 => to_unsigned(901, 10), 396 => to_unsigned(289, 10), 397 => to_unsigned(288, 10), 398 => to_unsigned(714, 10), 399 => to_unsigned(114, 10), 400 => to_unsigned(425, 10), 401 => to_unsigned(638, 10), 402 => to_unsigned(554, 10), 403 => to_unsigned(635, 10), 404 => to_unsigned(690, 10), 405 => to_unsigned(502, 10), 406 => to_unsigned(590, 10), 407 => to_unsigned(283, 10), 408 => to_unsigned(304, 10), 409 => to_unsigned(779, 10), 410 => to_unsigned(563, 10), 411 => to_unsigned(455, 10), 412 => to_unsigned(12, 10), 413 => to_unsigned(96, 10), 414 => to_unsigned(566, 10), 415 => to_unsigned(183, 10), 416 => to_unsigned(11, 10), 417 => to_unsigned(443, 10), 418 => to_unsigned(90, 10), 419 => to_unsigned(883, 10), 420 => to_unsigned(5, 10), 421 => to_unsigned(1021, 10), 422 => to_unsigned(170, 10), 423 => to_unsigned(503, 10), 424 => to_unsigned(815, 10), 425 => to_unsigned(264, 10), 426 => to_unsigned(533, 10), 427 => to_unsigned(710, 10), 428 => to_unsigned(728, 10), 429 => to_unsigned(744, 10), 430 => to_unsigned(229, 10), 431 => to_unsigned(541, 10), 432 => to_unsigned(781, 10), 433 => to_unsigned(547, 10), 434 => to_unsigned(5, 10), 435 => to_unsigned(1012, 10), 436 => to_unsigned(117, 10), 437 => to_unsigned(205, 10), 438 => to_unsigned(677, 10), 439 => to_unsigned(542, 10), 440 => to_unsigned(608, 10), 441 => to_unsigned(450, 10), 442 => to_unsigned(52, 10), 443 => to_unsigned(77, 10), 444 => to_unsigned(118, 10), 445 => to_unsigned(955, 10), 446 => to_unsigned(381, 10), 447 => to_unsigned(990, 10), 448 => to_unsigned(896, 10), 449 => to_unsigned(649, 10), 450 => to_unsigned(402, 10), 451 => to_unsigned(431, 10), 452 => to_unsigned(400, 10), 453 => to_unsigned(43, 10), 454 => to_unsigned(553, 10), 455 => to_unsigned(207, 10), 456 => to_unsigned(533, 10), 457 => to_unsigned(21, 10), 458 => to_unsigned(246, 10), 459 => to_unsigned(619, 10), 460 => to_unsigned(667, 10), 461 => to_unsigned(958, 10), 462 => to_unsigned(494, 10), 463 => to_unsigned(153, 10), 464 => to_unsigned(772, 10), 465 => to_unsigned(728, 10), 466 => to_unsigned(648, 10), 467 => to_unsigned(309, 10), 468 => to_unsigned(215, 10), 469 => to_unsigned(347, 10), 470 => to_unsigned(872, 10), 471 => to_unsigned(101, 10), 472 => to_unsigned(156, 10), 473 => to_unsigned(490, 10), 474 => to_unsigned(879, 10), 475 => to_unsigned(798, 10), 476 => to_unsigned(737, 10), 477 => to_unsigned(973, 10), 478 => to_unsigned(307, 10), 479 => to_unsigned(232, 10), 480 => to_unsigned(982, 10), 481 => to_unsigned(465, 10), 482 => to_unsigned(938, 10), 483 => to_unsigned(579, 10), 484 => to_unsigned(551, 10), 485 => to_unsigned(724, 10), 486 => to_unsigned(770, 10), 487 => to_unsigned(799, 10), 488 => to_unsigned(719, 10), 489 => to_unsigned(510, 10), 490 => to_unsigned(777, 10), 491 => to_unsigned(338, 10), 492 => to_unsigned(484, 10), 493 => to_unsigned(599, 10), 494 => to_unsigned(337, 10), 495 => to_unsigned(83, 10), 496 => to_unsigned(579, 10), 497 => to_unsigned(997, 10), 498 => to_unsigned(393, 10), 499 => to_unsigned(195, 10), 500 => to_unsigned(502, 10), 501 => to_unsigned(454, 10), 502 => to_unsigned(80, 10), 503 => to_unsigned(360, 10), 504 => to_unsigned(235, 10), 505 => to_unsigned(983, 10), 506 => to_unsigned(990, 10), 507 => to_unsigned(100, 10), 508 => to_unsigned(474, 10), 509 => to_unsigned(25, 10), 510 => to_unsigned(739, 10), 511 => to_unsigned(44, 10), 512 => to_unsigned(225, 10), 513 => to_unsigned(560, 10), 514 => to_unsigned(992, 10), 515 => to_unsigned(68, 10), 516 => to_unsigned(353, 10), 517 => to_unsigned(14, 10), 518 => to_unsigned(216, 10), 519 => to_unsigned(1009, 10), 520 => to_unsigned(135, 10), 521 => to_unsigned(45, 10), 522 => to_unsigned(242, 10), 523 => to_unsigned(740, 10), 524 => to_unsigned(769, 10), 525 => to_unsigned(611, 10), 526 => to_unsigned(80, 10), 527 => to_unsigned(994, 10), 528 => to_unsigned(368, 10), 529 => to_unsigned(888, 10), 530 => to_unsigned(262, 10), 531 => to_unsigned(968, 10), 532 => to_unsigned(109, 10), 533 => to_unsigned(502, 10), 534 => to_unsigned(670, 10), 535 => to_unsigned(137, 10), 536 => to_unsigned(265, 10), 537 => to_unsigned(237, 10), 538 => to_unsigned(398, 10), 539 => to_unsigned(240, 10), 540 => to_unsigned(70, 10), 541 => to_unsigned(10, 10), 542 => to_unsigned(907, 10), 543 => to_unsigned(694, 10), 544 => to_unsigned(866, 10), 545 => to_unsigned(748, 10), 546 => to_unsigned(453, 10), 547 => to_unsigned(879, 10), 548 => to_unsigned(408, 10), 549 => to_unsigned(470, 10), 550 => to_unsigned(282, 10), 551 => to_unsigned(114, 10), 552 => to_unsigned(448, 10), 553 => to_unsigned(186, 10), 554 => to_unsigned(291, 10), 555 => to_unsigned(619, 10), 556 => to_unsigned(770, 10), 557 => to_unsigned(51, 10), 558 => to_unsigned(65, 10), 559 => to_unsigned(826, 10), 560 => to_unsigned(135, 10), 561 => to_unsigned(338, 10), 562 => to_unsigned(748, 10), 563 => to_unsigned(613, 10), 564 => to_unsigned(368, 10), 565 => to_unsigned(16, 10), 566 => to_unsigned(728, 10), 567 => to_unsigned(53, 10), 568 => to_unsigned(212, 10), 569 => to_unsigned(740, 10), 570 => to_unsigned(641, 10), 571 => to_unsigned(687, 10), 572 => to_unsigned(522, 10), 573 => to_unsigned(517, 10), 574 => to_unsigned(349, 10), 575 => to_unsigned(142, 10), 576 => to_unsigned(145, 10), 577 => to_unsigned(94, 10), 578 => to_unsigned(15, 10), 579 => to_unsigned(766, 10), 580 => to_unsigned(430, 10), 581 => to_unsigned(175, 10), 582 => to_unsigned(659, 10), 583 => to_unsigned(767, 10), 584 => to_unsigned(565, 10), 585 => to_unsigned(950, 10), 586 => to_unsigned(936, 10), 587 => to_unsigned(381, 10), 588 => to_unsigned(430, 10), 589 => to_unsigned(664, 10), 590 => to_unsigned(49, 10), 591 => to_unsigned(464, 10), 592 => to_unsigned(536, 10), 593 => to_unsigned(716, 10), 594 => to_unsigned(993, 10), 595 => to_unsigned(243, 10), 596 => to_unsigned(444, 10), 597 => to_unsigned(1021, 10), 598 => to_unsigned(452, 10), 599 => to_unsigned(148, 10), 600 => to_unsigned(309, 10), 601 => to_unsigned(597, 10), 602 => to_unsigned(441, 10), 603 => to_unsigned(69, 10), 604 => to_unsigned(935, 10), 605 => to_unsigned(863, 10), 606 => to_unsigned(128, 10), 607 => to_unsigned(652, 10), 608 => to_unsigned(101, 10), 609 => to_unsigned(982, 10), 610 => to_unsigned(174, 10), 611 => to_unsigned(985, 10), 612 => to_unsigned(87, 10), 613 => to_unsigned(748, 10), 614 => to_unsigned(727, 10), 615 => to_unsigned(732, 10), 616 => to_unsigned(487, 10), 617 => to_unsigned(28, 10), 618 => to_unsigned(935, 10), 619 => to_unsigned(392, 10), 620 => to_unsigned(357, 10), 621 => to_unsigned(740, 10), 622 => to_unsigned(785, 10), 623 => to_unsigned(207, 10), 624 => to_unsigned(437, 10), 625 => to_unsigned(340, 10), 626 => to_unsigned(321, 10), 627 => to_unsigned(244, 10), 628 => to_unsigned(15, 10), 629 => to_unsigned(242, 10), 630 => to_unsigned(613, 10), 631 => to_unsigned(316, 10), 632 => to_unsigned(634, 10), 633 => to_unsigned(776, 10), 634 => to_unsigned(700, 10), 635 => to_unsigned(577, 10), 636 => to_unsigned(182, 10), 637 => to_unsigned(464, 10), 638 => to_unsigned(207, 10), 639 => to_unsigned(425, 10), 640 => to_unsigned(641, 10), 641 => to_unsigned(232, 10), 642 => to_unsigned(639, 10), 643 => to_unsigned(959, 10), 644 => to_unsigned(638, 10), 645 => to_unsigned(142, 10), 646 => to_unsigned(276, 10), 647 => to_unsigned(771, 10), 648 => to_unsigned(156, 10), 649 => to_unsigned(352, 10), 650 => to_unsigned(696, 10), 651 => to_unsigned(863, 10), 652 => to_unsigned(161, 10), 653 => to_unsigned(414, 10), 654 => to_unsigned(347, 10), 655 => to_unsigned(23, 10), 656 => to_unsigned(561, 10), 657 => to_unsigned(701, 10), 658 => to_unsigned(254, 10), 659 => to_unsigned(453, 10), 660 => to_unsigned(875, 10), 661 => to_unsigned(117, 10), 662 => to_unsigned(671, 10), 663 => to_unsigned(3, 10), 664 => to_unsigned(38, 10), 665 => to_unsigned(823, 10), 666 => to_unsigned(114, 10), 667 => to_unsigned(614, 10), 668 => to_unsigned(49, 10), 669 => to_unsigned(78, 10), 670 => to_unsigned(258, 10), 671 => to_unsigned(99, 10), 672 => to_unsigned(237, 10), 673 => to_unsigned(983, 10), 674 => to_unsigned(12, 10), 675 => to_unsigned(841, 10), 676 => to_unsigned(310, 10), 677 => to_unsigned(607, 10), 678 => to_unsigned(726, 10), 679 => to_unsigned(512, 10), 680 => to_unsigned(801, 10), 681 => to_unsigned(355, 10), 682 => to_unsigned(994, 10), 683 => to_unsigned(35, 10), 684 => to_unsigned(960, 10), 685 => to_unsigned(172, 10), 686 => to_unsigned(349, 10), 687 => to_unsigned(44, 10), 688 => to_unsigned(638, 10), 689 => to_unsigned(784, 10), 690 => to_unsigned(450, 10), 691 => to_unsigned(387, 10), 692 => to_unsigned(929, 10), 693 => to_unsigned(47, 10), 694 => to_unsigned(21, 10), 695 => to_unsigned(482, 10), 696 => to_unsigned(157, 10), 697 => to_unsigned(251, 10), 698 => to_unsigned(185, 10), 699 => to_unsigned(881, 10), 700 => to_unsigned(686, 10), 701 => to_unsigned(464, 10), 702 => to_unsigned(769, 10), 703 => to_unsigned(29, 10), 704 => to_unsigned(795, 10), 705 => to_unsigned(146, 10), 706 => to_unsigned(551, 10), 707 => to_unsigned(246, 10), 708 => to_unsigned(172, 10), 709 => to_unsigned(852, 10), 710 => to_unsigned(778, 10), 711 => to_unsigned(320, 10), 712 => to_unsigned(442, 10), 713 => to_unsigned(417, 10), 714 => to_unsigned(812, 10), 715 => to_unsigned(589, 10), 716 => to_unsigned(659, 10), 717 => to_unsigned(636, 10), 718 => to_unsigned(590, 10), 719 => to_unsigned(430, 10), 720 => to_unsigned(849, 10), 721 => to_unsigned(981, 10), 722 => to_unsigned(589, 10), 723 => to_unsigned(924, 10), 724 => to_unsigned(270, 10), 725 => to_unsigned(962, 10), 726 => to_unsigned(627, 10), 727 => to_unsigned(559, 10), 728 => to_unsigned(798, 10), 729 => to_unsigned(946, 10), 730 => to_unsigned(830, 10), 731 => to_unsigned(247, 10), 732 => to_unsigned(383, 10), 733 => to_unsigned(33, 10), 734 => to_unsigned(714, 10), 735 => to_unsigned(127, 10), 736 => to_unsigned(762, 10), 737 => to_unsigned(616, 10), 738 => to_unsigned(229, 10), 739 => to_unsigned(217, 10), 740 => to_unsigned(47, 10), 741 => to_unsigned(620, 10), 742 => to_unsigned(1003, 10), 743 => to_unsigned(937, 10), 744 => to_unsigned(631, 10), 745 => to_unsigned(545, 10), 746 => to_unsigned(512, 10), 747 => to_unsigned(261, 10), 748 => to_unsigned(618, 10), 749 => to_unsigned(574, 10), 750 => to_unsigned(171, 10), 751 => to_unsigned(794, 10), 752 => to_unsigned(831, 10), 753 => to_unsigned(553, 10), 754 => to_unsigned(795, 10), 755 => to_unsigned(526, 10), 756 => to_unsigned(495, 10), 757 => to_unsigned(624, 10), 758 => to_unsigned(258, 10), 759 => to_unsigned(19, 10), 760 => to_unsigned(140, 10), 761 => to_unsigned(880, 10), 762 => to_unsigned(287, 10), 763 => to_unsigned(689, 10), 764 => to_unsigned(550, 10), 765 => to_unsigned(478, 10), 766 => to_unsigned(566, 10), 767 => to_unsigned(747, 10), 768 => to_unsigned(769, 10), 769 => to_unsigned(634, 10), 770 => to_unsigned(801, 10), 771 => to_unsigned(575, 10), 772 => to_unsigned(487, 10), 773 => to_unsigned(433, 10), 774 => to_unsigned(848, 10), 775 => to_unsigned(1018, 10), 776 => to_unsigned(812, 10), 777 => to_unsigned(114, 10), 778 => to_unsigned(12, 10), 779 => to_unsigned(155, 10), 780 => to_unsigned(86, 10), 781 => to_unsigned(110, 10), 782 => to_unsigned(750, 10), 783 => to_unsigned(716, 10), 784 => to_unsigned(613, 10), 785 => to_unsigned(115, 10), 786 => to_unsigned(141, 10), 787 => to_unsigned(630, 10), 788 => to_unsigned(839, 10), 789 => to_unsigned(931, 10), 790 => to_unsigned(748, 10), 791 => to_unsigned(958, 10), 792 => to_unsigned(61, 10), 793 => to_unsigned(214, 10), 794 => to_unsigned(235, 10), 795 => to_unsigned(468, 10), 796 => to_unsigned(800, 10), 797 => to_unsigned(829, 10), 798 => to_unsigned(1022, 10), 799 => to_unsigned(243, 10), 800 => to_unsigned(690, 10), 801 => to_unsigned(415, 10), 802 => to_unsigned(181, 10), 803 => to_unsigned(338, 10), 804 => to_unsigned(231, 10), 805 => to_unsigned(443, 10), 806 => to_unsigned(563, 10), 807 => to_unsigned(906, 10), 808 => to_unsigned(970, 10), 809 => to_unsigned(230, 10), 810 => to_unsigned(92, 10), 811 => to_unsigned(314, 10), 812 => to_unsigned(929, 10), 813 => to_unsigned(607, 10), 814 => to_unsigned(572, 10), 815 => to_unsigned(284, 10), 816 => to_unsigned(592, 10), 817 => to_unsigned(361, 10), 818 => to_unsigned(764, 10), 819 => to_unsigned(625, 10), 820 => to_unsigned(273, 10), 821 => to_unsigned(336, 10), 822 => to_unsigned(218, 10), 823 => to_unsigned(845, 10), 824 => to_unsigned(963, 10), 825 => to_unsigned(454, 10), 826 => to_unsigned(145, 10), 827 => to_unsigned(264, 10), 828 => to_unsigned(732, 10), 829 => to_unsigned(471, 10), 830 => to_unsigned(551, 10), 831 => to_unsigned(282, 10), 832 => to_unsigned(91, 10), 833 => to_unsigned(162, 10), 834 => to_unsigned(287, 10), 835 => to_unsigned(190, 10), 836 => to_unsigned(350, 10), 837 => to_unsigned(425, 10), 838 => to_unsigned(223, 10), 839 => to_unsigned(342, 10), 840 => to_unsigned(701, 10), 841 => to_unsigned(11, 10), 842 => to_unsigned(356, 10), 843 => to_unsigned(83, 10), 844 => to_unsigned(999, 10), 845 => to_unsigned(563, 10), 846 => to_unsigned(798, 10), 847 => to_unsigned(23, 10), 848 => to_unsigned(643, 10), 849 => to_unsigned(59, 10), 850 => to_unsigned(511, 10), 851 => to_unsigned(339, 10), 852 => to_unsigned(885, 10), 853 => to_unsigned(609, 10), 854 => to_unsigned(827, 10), 855 => to_unsigned(5, 10), 856 => to_unsigned(171, 10), 857 => to_unsigned(26, 10), 858 => to_unsigned(1011, 10), 859 => to_unsigned(370, 10), 860 => to_unsigned(45, 10), 861 => to_unsigned(661, 10), 862 => to_unsigned(186, 10), 863 => to_unsigned(239, 10), 864 => to_unsigned(577, 10), 865 => to_unsigned(963, 10), 866 => to_unsigned(555, 10), 867 => to_unsigned(977, 10), 868 => to_unsigned(461, 10), 869 => to_unsigned(432, 10), 870 => to_unsigned(482, 10), 871 => to_unsigned(326, 10), 872 => to_unsigned(976, 10), 873 => to_unsigned(590, 10), 874 => to_unsigned(44, 10), 875 => to_unsigned(828, 10), 876 => to_unsigned(479, 10), 877 => to_unsigned(37, 10), 878 => to_unsigned(601, 10), 879 => to_unsigned(734, 10), 880 => to_unsigned(225, 10), 881 => to_unsigned(318, 10), 882 => to_unsigned(658, 10), 883 => to_unsigned(576, 10), 884 => to_unsigned(939, 10), 885 => to_unsigned(86, 10), 886 => to_unsigned(627, 10), 887 => to_unsigned(487, 10), 888 => to_unsigned(932, 10), 889 => to_unsigned(322, 10), 890 => to_unsigned(465, 10), 891 => to_unsigned(434, 10), 892 => to_unsigned(715, 10), 893 => to_unsigned(257, 10), 894 => to_unsigned(650, 10), 895 => to_unsigned(328, 10), 896 => to_unsigned(175, 10), 897 => to_unsigned(481, 10), 898 => to_unsigned(51, 10), 899 => to_unsigned(291, 10), 900 => to_unsigned(865, 10), 901 => to_unsigned(461, 10), 902 => to_unsigned(71, 10), 903 => to_unsigned(242, 10), 904 => to_unsigned(426, 10), 905 => to_unsigned(558, 10), 906 => to_unsigned(619, 10), 907 => to_unsigned(620, 10), 908 => to_unsigned(671, 10), 909 => to_unsigned(426, 10), 910 => to_unsigned(126, 10), 911 => to_unsigned(568, 10), 912 => to_unsigned(468, 10), 913 => to_unsigned(985, 10), 914 => to_unsigned(116, 10), 915 => to_unsigned(736, 10), 916 => to_unsigned(0, 10), 917 => to_unsigned(637, 10), 918 => to_unsigned(193, 10), 919 => to_unsigned(430, 10), 920 => to_unsigned(892, 10), 921 => to_unsigned(451, 10), 922 => to_unsigned(578, 10), 923 => to_unsigned(203, 10), 924 => to_unsigned(942, 10), 925 => to_unsigned(760, 10), 926 => to_unsigned(612, 10), 927 => to_unsigned(345, 10), 928 => to_unsigned(536, 10), 929 => to_unsigned(318, 10), 930 => to_unsigned(838, 10), 931 => to_unsigned(746, 10), 932 => to_unsigned(885, 10), 933 => to_unsigned(254, 10), 934 => to_unsigned(691, 10), 935 => to_unsigned(228, 10), 936 => to_unsigned(760, 10), 937 => to_unsigned(349, 10), 938 => to_unsigned(470, 10), 939 => to_unsigned(366, 10), 940 => to_unsigned(934, 10), 941 => to_unsigned(356, 10), 942 => to_unsigned(397, 10), 943 => to_unsigned(552, 10), 944 => to_unsigned(603, 10), 945 => to_unsigned(237, 10), 946 => to_unsigned(555, 10), 947 => to_unsigned(529, 10), 948 => to_unsigned(310, 10), 949 => to_unsigned(237, 10), 950 => to_unsigned(712, 10), 951 => to_unsigned(655, 10), 952 => to_unsigned(840, 10), 953 => to_unsigned(578, 10), 954 => to_unsigned(152, 10), 955 => to_unsigned(974, 10), 956 => to_unsigned(975, 10), 957 => to_unsigned(810, 10), 958 => to_unsigned(371, 10), 959 => to_unsigned(206, 10), 960 => to_unsigned(11, 10), 961 => to_unsigned(560, 10), 962 => to_unsigned(632, 10), 963 => to_unsigned(446, 10), 964 => to_unsigned(238, 10), 965 => to_unsigned(426, 10), 966 => to_unsigned(93, 10), 967 => to_unsigned(603, 10), 968 => to_unsigned(988, 10), 969 => to_unsigned(729, 10), 970 => to_unsigned(237, 10), 971 => to_unsigned(516, 10), 972 => to_unsigned(809, 10), 973 => to_unsigned(848, 10), 974 => to_unsigned(304, 10), 975 => to_unsigned(117, 10), 976 => to_unsigned(330, 10), 977 => to_unsigned(380, 10), 978 => to_unsigned(76, 10), 979 => to_unsigned(230, 10), 980 => to_unsigned(243, 10), 981 => to_unsigned(332, 10), 982 => to_unsigned(568, 10), 983 => to_unsigned(392, 10), 984 => to_unsigned(344, 10), 985 => to_unsigned(951, 10), 986 => to_unsigned(442, 10), 987 => to_unsigned(605, 10), 988 => to_unsigned(619, 10), 989 => to_unsigned(490, 10), 990 => to_unsigned(556, 10), 991 => to_unsigned(884, 10), 992 => to_unsigned(614, 10), 993 => to_unsigned(572, 10), 994 => to_unsigned(702, 10), 995 => to_unsigned(818, 10), 996 => to_unsigned(854, 10), 997 => to_unsigned(348, 10), 998 => to_unsigned(603, 10), 999 => to_unsigned(819, 10), 1000 => to_unsigned(592, 10), 1001 => to_unsigned(769, 10), 1002 => to_unsigned(280, 10), 1003 => to_unsigned(53, 10), 1004 => to_unsigned(997, 10), 1005 => to_unsigned(536, 10), 1006 => to_unsigned(963, 10), 1007 => to_unsigned(55, 10), 1008 => to_unsigned(870, 10), 1009 => to_unsigned(939, 10), 1010 => to_unsigned(991, 10), 1011 => to_unsigned(159, 10), 1012 => to_unsigned(166, 10), 1013 => to_unsigned(850, 10), 1014 => to_unsigned(461, 10), 1015 => to_unsigned(350, 10), 1016 => to_unsigned(708, 10), 1017 => to_unsigned(777, 10), 1018 => to_unsigned(93, 10), 1019 => to_unsigned(794, 10), 1020 => to_unsigned(1010, 10), 1021 => to_unsigned(483, 10), 1022 => to_unsigned(291, 10), 1023 => to_unsigned(671, 10), 1024 => to_unsigned(716, 10), 1025 => to_unsigned(273, 10), 1026 => to_unsigned(968, 10), 1027 => to_unsigned(732, 10), 1028 => to_unsigned(527, 10), 1029 => to_unsigned(860, 10), 1030 => to_unsigned(40, 10), 1031 => to_unsigned(893, 10), 1032 => to_unsigned(180, 10), 1033 => to_unsigned(1023, 10), 1034 => to_unsigned(994, 10), 1035 => to_unsigned(447, 10), 1036 => to_unsigned(660, 10), 1037 => to_unsigned(210, 10), 1038 => to_unsigned(943, 10), 1039 => to_unsigned(128, 10), 1040 => to_unsigned(111, 10), 1041 => to_unsigned(979, 10), 1042 => to_unsigned(140, 10), 1043 => to_unsigned(917, 10), 1044 => to_unsigned(21, 10), 1045 => to_unsigned(562, 10), 1046 => to_unsigned(826, 10), 1047 => to_unsigned(327, 10), 1048 => to_unsigned(890, 10), 1049 => to_unsigned(370, 10), 1050 => to_unsigned(662, 10), 1051 => to_unsigned(521, 10), 1052 => to_unsigned(192, 10), 1053 => to_unsigned(721, 10), 1054 => to_unsigned(389, 10), 1055 => to_unsigned(588, 10), 1056 => to_unsigned(304, 10), 1057 => to_unsigned(257, 10), 1058 => to_unsigned(701, 10), 1059 => to_unsigned(903, 10), 1060 => to_unsigned(995, 10), 1061 => to_unsigned(92, 10), 1062 => to_unsigned(825, 10), 1063 => to_unsigned(848, 10), 1064 => to_unsigned(157, 10), 1065 => to_unsigned(610, 10), 1066 => to_unsigned(193, 10), 1067 => to_unsigned(804, 10), 1068 => to_unsigned(272, 10), 1069 => to_unsigned(940, 10), 1070 => to_unsigned(220, 10), 1071 => to_unsigned(898, 10), 1072 => to_unsigned(128, 10), 1073 => to_unsigned(147, 10), 1074 => to_unsigned(746, 10), 1075 => to_unsigned(279, 10), 1076 => to_unsigned(617, 10), 1077 => to_unsigned(146, 10), 1078 => to_unsigned(388, 10), 1079 => to_unsigned(771, 10), 1080 => to_unsigned(900, 10), 1081 => to_unsigned(109, 10), 1082 => to_unsigned(253, 10), 1083 => to_unsigned(346, 10), 1084 => to_unsigned(231, 10), 1085 => to_unsigned(335, 10), 1086 => to_unsigned(902, 10), 1087 => to_unsigned(756, 10), 1088 => to_unsigned(127, 10), 1089 => to_unsigned(602, 10), 1090 => to_unsigned(513, 10), 1091 => to_unsigned(756, 10), 1092 => to_unsigned(956, 10), 1093 => to_unsigned(70, 10), 1094 => to_unsigned(800, 10), 1095 => to_unsigned(173, 10), 1096 => to_unsigned(597, 10), 1097 => to_unsigned(709, 10), 1098 => to_unsigned(13, 10), 1099 => to_unsigned(999, 10), 1100 => to_unsigned(126, 10), 1101 => to_unsigned(154, 10), 1102 => to_unsigned(26, 10), 1103 => to_unsigned(790, 10), 1104 => to_unsigned(589, 10), 1105 => to_unsigned(52, 10), 1106 => to_unsigned(360, 10), 1107 => to_unsigned(884, 10), 1108 => to_unsigned(790, 10), 1109 => to_unsigned(656, 10), 1110 => to_unsigned(24, 10), 1111 => to_unsigned(748, 10), 1112 => to_unsigned(524, 10), 1113 => to_unsigned(77, 10), 1114 => to_unsigned(939, 10), 1115 => to_unsigned(868, 10), 1116 => to_unsigned(216, 10), 1117 => to_unsigned(167, 10), 1118 => to_unsigned(1021, 10), 1119 => to_unsigned(548, 10), 1120 => to_unsigned(378, 10), 1121 => to_unsigned(874, 10), 1122 => to_unsigned(237, 10), 1123 => to_unsigned(581, 10), 1124 => to_unsigned(196, 10), 1125 => to_unsigned(360, 10), 1126 => to_unsigned(631, 10), 1127 => to_unsigned(274, 10), 1128 => to_unsigned(547, 10), 1129 => to_unsigned(1, 10), 1130 => to_unsigned(250, 10), 1131 => to_unsigned(674, 10), 1132 => to_unsigned(708, 10), 1133 => to_unsigned(236, 10), 1134 => to_unsigned(216, 10), 1135 => to_unsigned(579, 10), 1136 => to_unsigned(51, 10), 1137 => to_unsigned(752, 10), 1138 => to_unsigned(729, 10), 1139 => to_unsigned(764, 10), 1140 => to_unsigned(491, 10), 1141 => to_unsigned(713, 10), 1142 => to_unsigned(533, 10), 1143 => to_unsigned(247, 10), 1144 => to_unsigned(401, 10), 1145 => to_unsigned(527, 10), 1146 => to_unsigned(799, 10), 1147 => to_unsigned(495, 10), 1148 => to_unsigned(790, 10), 1149 => to_unsigned(149, 10), 1150 => to_unsigned(576, 10), 1151 => to_unsigned(877, 10), 1152 => to_unsigned(745, 10), 1153 => to_unsigned(1023, 10), 1154 => to_unsigned(88, 10), 1155 => to_unsigned(147, 10), 1156 => to_unsigned(739, 10), 1157 => to_unsigned(868, 10), 1158 => to_unsigned(385, 10), 1159 => to_unsigned(558, 10), 1160 => to_unsigned(822, 10), 1161 => to_unsigned(123, 10), 1162 => to_unsigned(299, 10), 1163 => to_unsigned(925, 10), 1164 => to_unsigned(697, 10), 1165 => to_unsigned(278, 10), 1166 => to_unsigned(412, 10), 1167 => to_unsigned(596, 10), 1168 => to_unsigned(339, 10), 1169 => to_unsigned(305, 10), 1170 => to_unsigned(562, 10), 1171 => to_unsigned(9, 10), 1172 => to_unsigned(995, 10), 1173 => to_unsigned(802, 10), 1174 => to_unsigned(82, 10), 1175 => to_unsigned(105, 10), 1176 => to_unsigned(932, 10), 1177 => to_unsigned(756, 10), 1178 => to_unsigned(681, 10), 1179 => to_unsigned(75, 10), 1180 => to_unsigned(949, 10), 1181 => to_unsigned(599, 10), 1182 => to_unsigned(975, 10), 1183 => to_unsigned(462, 10), 1184 => to_unsigned(143, 10), 1185 => to_unsigned(241, 10), 1186 => to_unsigned(854, 10), 1187 => to_unsigned(517, 10), 1188 => to_unsigned(935, 10), 1189 => to_unsigned(801, 10), 1190 => to_unsigned(677, 10), 1191 => to_unsigned(921, 10), 1192 => to_unsigned(842, 10), 1193 => to_unsigned(726, 10), 1194 => to_unsigned(156, 10), 1195 => to_unsigned(538, 10), 1196 => to_unsigned(532, 10), 1197 => to_unsigned(869, 10), 1198 => to_unsigned(903, 10), 1199 => to_unsigned(251, 10), 1200 => to_unsigned(374, 10), 1201 => to_unsigned(736, 10), 1202 => to_unsigned(386, 10), 1203 => to_unsigned(501, 10), 1204 => to_unsigned(557, 10), 1205 => to_unsigned(109, 10), 1206 => to_unsigned(590, 10), 1207 => to_unsigned(392, 10), 1208 => to_unsigned(809, 10), 1209 => to_unsigned(910, 10), 1210 => to_unsigned(132, 10), 1211 => to_unsigned(162, 10), 1212 => to_unsigned(199, 10), 1213 => to_unsigned(145, 10), 1214 => to_unsigned(134, 10), 1215 => to_unsigned(122, 10), 1216 => to_unsigned(148, 10), 1217 => to_unsigned(711, 10), 1218 => to_unsigned(272, 10), 1219 => to_unsigned(1021, 10), 1220 => to_unsigned(340, 10), 1221 => to_unsigned(330, 10), 1222 => to_unsigned(797, 10), 1223 => to_unsigned(218, 10), 1224 => to_unsigned(473, 10), 1225 => to_unsigned(553, 10), 1226 => to_unsigned(988, 10), 1227 => to_unsigned(333, 10), 1228 => to_unsigned(980, 10), 1229 => to_unsigned(857, 10), 1230 => to_unsigned(534, 10), 1231 => to_unsigned(784, 10), 1232 => to_unsigned(761, 10), 1233 => to_unsigned(773, 10), 1234 => to_unsigned(482, 10), 1235 => to_unsigned(621, 10), 1236 => to_unsigned(605, 10), 1237 => to_unsigned(538, 10), 1238 => to_unsigned(1010, 10), 1239 => to_unsigned(36, 10), 1240 => to_unsigned(613, 10), 1241 => to_unsigned(935, 10), 1242 => to_unsigned(12, 10), 1243 => to_unsigned(550, 10), 1244 => to_unsigned(867, 10), 1245 => to_unsigned(452, 10), 1246 => to_unsigned(431, 10), 1247 => to_unsigned(350, 10), 1248 => to_unsigned(115, 10), 1249 => to_unsigned(403, 10), 1250 => to_unsigned(823, 10), 1251 => to_unsigned(206, 10), 1252 => to_unsigned(502, 10), 1253 => to_unsigned(325, 10), 1254 => to_unsigned(251, 10), 1255 => to_unsigned(850, 10), 1256 => to_unsigned(190, 10), 1257 => to_unsigned(653, 10), 1258 => to_unsigned(186, 10), 1259 => to_unsigned(30, 10), 1260 => to_unsigned(738, 10), 1261 => to_unsigned(913, 10), 1262 => to_unsigned(636, 10), 1263 => to_unsigned(237, 10), 1264 => to_unsigned(120, 10), 1265 => to_unsigned(925, 10), 1266 => to_unsigned(840, 10), 1267 => to_unsigned(929, 10), 1268 => to_unsigned(62, 10), 1269 => to_unsigned(576, 10), 1270 => to_unsigned(322, 10), 1271 => to_unsigned(421, 10), 1272 => to_unsigned(227, 10), 1273 => to_unsigned(454, 10), 1274 => to_unsigned(756, 10), 1275 => to_unsigned(224, 10), 1276 => to_unsigned(900, 10), 1277 => to_unsigned(882, 10), 1278 => to_unsigned(138, 10), 1279 => to_unsigned(176, 10), 1280 => to_unsigned(324, 10), 1281 => to_unsigned(531, 10), 1282 => to_unsigned(485, 10), 1283 => to_unsigned(223, 10), 1284 => to_unsigned(881, 10), 1285 => to_unsigned(983, 10), 1286 => to_unsigned(1011, 10), 1287 => to_unsigned(438, 10), 1288 => to_unsigned(843, 10), 1289 => to_unsigned(49, 10), 1290 => to_unsigned(450, 10), 1291 => to_unsigned(332, 10), 1292 => to_unsigned(24, 10), 1293 => to_unsigned(577, 10), 1294 => to_unsigned(454, 10), 1295 => to_unsigned(653, 10), 1296 => to_unsigned(481, 10), 1297 => to_unsigned(701, 10), 1298 => to_unsigned(550, 10), 1299 => to_unsigned(383, 10), 1300 => to_unsigned(710, 10), 1301 => to_unsigned(999, 10), 1302 => to_unsigned(105, 10), 1303 => to_unsigned(113, 10), 1304 => to_unsigned(247, 10), 1305 => to_unsigned(998, 10), 1306 => to_unsigned(430, 10), 1307 => to_unsigned(1019, 10), 1308 => to_unsigned(641, 10), 1309 => to_unsigned(1000, 10), 1310 => to_unsigned(231, 10), 1311 => to_unsigned(580, 10), 1312 => to_unsigned(89, 10), 1313 => to_unsigned(350, 10), 1314 => to_unsigned(32, 10), 1315 => to_unsigned(441, 10), 1316 => to_unsigned(1, 10), 1317 => to_unsigned(754, 10), 1318 => to_unsigned(475, 10), 1319 => to_unsigned(316, 10), 1320 => to_unsigned(29, 10), 1321 => to_unsigned(925, 10), 1322 => to_unsigned(782, 10), 1323 => to_unsigned(224, 10), 1324 => to_unsigned(701, 10), 1325 => to_unsigned(137, 10), 1326 => to_unsigned(862, 10), 1327 => to_unsigned(841, 10), 1328 => to_unsigned(666, 10), 1329 => to_unsigned(112, 10), 1330 => to_unsigned(461, 10), 1331 => to_unsigned(517, 10), 1332 => to_unsigned(592, 10), 1333 => to_unsigned(395, 10), 1334 => to_unsigned(778, 10), 1335 => to_unsigned(922, 10), 1336 => to_unsigned(389, 10), 1337 => to_unsigned(576, 10), 1338 => to_unsigned(529, 10), 1339 => to_unsigned(996, 10), 1340 => to_unsigned(309, 10), 1341 => to_unsigned(675, 10), 1342 => to_unsigned(481, 10), 1343 => to_unsigned(842, 10), 1344 => to_unsigned(120, 10), 1345 => to_unsigned(512, 10), 1346 => to_unsigned(856, 10), 1347 => to_unsigned(462, 10), 1348 => to_unsigned(821, 10), 1349 => to_unsigned(115, 10), 1350 => to_unsigned(422, 10), 1351 => to_unsigned(38, 10), 1352 => to_unsigned(256, 10), 1353 => to_unsigned(69, 10), 1354 => to_unsigned(502, 10), 1355 => to_unsigned(531, 10), 1356 => to_unsigned(689, 10), 1357 => to_unsigned(645, 10), 1358 => to_unsigned(694, 10), 1359 => to_unsigned(458, 10), 1360 => to_unsigned(407, 10), 1361 => to_unsigned(866, 10), 1362 => to_unsigned(569, 10), 1363 => to_unsigned(777, 10), 1364 => to_unsigned(497, 10), 1365 => to_unsigned(367, 10), 1366 => to_unsigned(599, 10), 1367 => to_unsigned(144, 10), 1368 => to_unsigned(737, 10), 1369 => to_unsigned(660, 10), 1370 => to_unsigned(695, 10), 1371 => to_unsigned(106, 10), 1372 => to_unsigned(206, 10), 1373 => to_unsigned(445, 10), 1374 => to_unsigned(803, 10), 1375 => to_unsigned(479, 10), 1376 => to_unsigned(586, 10), 1377 => to_unsigned(947, 10), 1378 => to_unsigned(597, 10), 1379 => to_unsigned(53, 10), 1380 => to_unsigned(944, 10), 1381 => to_unsigned(273, 10), 1382 => to_unsigned(141, 10), 1383 => to_unsigned(696, 10), 1384 => to_unsigned(977, 10), 1385 => to_unsigned(450, 10), 1386 => to_unsigned(1003, 10), 1387 => to_unsigned(668, 10), 1388 => to_unsigned(591, 10), 1389 => to_unsigned(346, 10), 1390 => to_unsigned(516, 10), 1391 => to_unsigned(85, 10), 1392 => to_unsigned(393, 10), 1393 => to_unsigned(493, 10), 1394 => to_unsigned(997, 10), 1395 => to_unsigned(246, 10), 1396 => to_unsigned(618, 10), 1397 => to_unsigned(56, 10), 1398 => to_unsigned(457, 10), 1399 => to_unsigned(813, 10), 1400 => to_unsigned(241, 10), 1401 => to_unsigned(243, 10), 1402 => to_unsigned(276, 10), 1403 => to_unsigned(49, 10), 1404 => to_unsigned(649, 10), 1405 => to_unsigned(167, 10), 1406 => to_unsigned(485, 10), 1407 => to_unsigned(427, 10), 1408 => to_unsigned(603, 10), 1409 => to_unsigned(903, 10), 1410 => to_unsigned(90, 10), 1411 => to_unsigned(205, 10), 1412 => to_unsigned(985, 10), 1413 => to_unsigned(94, 10), 1414 => to_unsigned(492, 10), 1415 => to_unsigned(69, 10), 1416 => to_unsigned(287, 10), 1417 => to_unsigned(882, 10), 1418 => to_unsigned(630, 10), 1419 => to_unsigned(218, 10), 1420 => to_unsigned(821, 10), 1421 => to_unsigned(976, 10), 1422 => to_unsigned(972, 10), 1423 => to_unsigned(121, 10), 1424 => to_unsigned(538, 10), 1425 => to_unsigned(442, 10), 1426 => to_unsigned(972, 10), 1427 => to_unsigned(792, 10), 1428 => to_unsigned(524, 10), 1429 => to_unsigned(289, 10), 1430 => to_unsigned(917, 10), 1431 => to_unsigned(175, 10), 1432 => to_unsigned(1012, 10), 1433 => to_unsigned(381, 10), 1434 => to_unsigned(37, 10), 1435 => to_unsigned(97, 10), 1436 => to_unsigned(907, 10), 1437 => to_unsigned(893, 10), 1438 => to_unsigned(683, 10), 1439 => to_unsigned(43, 10), 1440 => to_unsigned(766, 10), 1441 => to_unsigned(348, 10), 1442 => to_unsigned(836, 10), 1443 => to_unsigned(42, 10), 1444 => to_unsigned(584, 10), 1445 => to_unsigned(197, 10), 1446 => to_unsigned(272, 10), 1447 => to_unsigned(971, 10), 1448 => to_unsigned(493, 10), 1449 => to_unsigned(916, 10), 1450 => to_unsigned(248, 10), 1451 => to_unsigned(977, 10), 1452 => to_unsigned(299, 10), 1453 => to_unsigned(2, 10), 1454 => to_unsigned(392, 10), 1455 => to_unsigned(693, 10), 1456 => to_unsigned(227, 10), 1457 => to_unsigned(182, 10), 1458 => to_unsigned(261, 10), 1459 => to_unsigned(823, 10), 1460 => to_unsigned(708, 10), 1461 => to_unsigned(643, 10), 1462 => to_unsigned(580, 10), 1463 => to_unsigned(425, 10), 1464 => to_unsigned(122, 10), 1465 => to_unsigned(370, 10), 1466 => to_unsigned(784, 10), 1467 => to_unsigned(1010, 10), 1468 => to_unsigned(224, 10), 1469 => to_unsigned(883, 10), 1470 => to_unsigned(892, 10), 1471 => to_unsigned(850, 10), 1472 => to_unsigned(795, 10), 1473 => to_unsigned(1013, 10), 1474 => to_unsigned(742, 10), 1475 => to_unsigned(826, 10), 1476 => to_unsigned(405, 10), 1477 => to_unsigned(425, 10), 1478 => to_unsigned(316, 10), 1479 => to_unsigned(811, 10), 1480 => to_unsigned(528, 10), 1481 => to_unsigned(899, 10), 1482 => to_unsigned(115, 10), 1483 => to_unsigned(311, 10), 1484 => to_unsigned(717, 10), 1485 => to_unsigned(949, 10), 1486 => to_unsigned(260, 10), 1487 => to_unsigned(877, 10), 1488 => to_unsigned(88, 10), 1489 => to_unsigned(695, 10), 1490 => to_unsigned(983, 10), 1491 => to_unsigned(406, 10), 1492 => to_unsigned(877, 10), 1493 => to_unsigned(438, 10), 1494 => to_unsigned(178, 10), 1495 => to_unsigned(280, 10), 1496 => to_unsigned(515, 10), 1497 => to_unsigned(66, 10), 1498 => to_unsigned(32, 10), 1499 => to_unsigned(851, 10), 1500 => to_unsigned(447, 10), 1501 => to_unsigned(343, 10), 1502 => to_unsigned(148, 10), 1503 => to_unsigned(498, 10), 1504 => to_unsigned(653, 10), 1505 => to_unsigned(676, 10), 1506 => to_unsigned(211, 10), 1507 => to_unsigned(532, 10), 1508 => to_unsigned(697, 10), 1509 => to_unsigned(290, 10), 1510 => to_unsigned(999, 10), 1511 => to_unsigned(3, 10), 1512 => to_unsigned(727, 10), 1513 => to_unsigned(828, 10), 1514 => to_unsigned(437, 10), 1515 => to_unsigned(226, 10), 1516 => to_unsigned(313, 10), 1517 => to_unsigned(91, 10), 1518 => to_unsigned(513, 10), 1519 => to_unsigned(937, 10), 1520 => to_unsigned(473, 10), 1521 => to_unsigned(19, 10), 1522 => to_unsigned(815, 10), 1523 => to_unsigned(618, 10), 1524 => to_unsigned(958, 10), 1525 => to_unsigned(720, 10), 1526 => to_unsigned(299, 10), 1527 => to_unsigned(313, 10), 1528 => to_unsigned(267, 10), 1529 => to_unsigned(685, 10), 1530 => to_unsigned(916, 10), 1531 => to_unsigned(925, 10), 1532 => to_unsigned(938, 10), 1533 => to_unsigned(583, 10), 1534 => to_unsigned(562, 10), 1535 => to_unsigned(139, 10), 1536 => to_unsigned(588, 10), 1537 => to_unsigned(763, 10), 1538 => to_unsigned(530, 10), 1539 => to_unsigned(966, 10), 1540 => to_unsigned(111, 10), 1541 => to_unsigned(72, 10), 1542 => to_unsigned(972, 10), 1543 => to_unsigned(18, 10), 1544 => to_unsigned(531, 10), 1545 => to_unsigned(576, 10), 1546 => to_unsigned(1012, 10), 1547 => to_unsigned(906, 10), 1548 => to_unsigned(358, 10), 1549 => to_unsigned(219, 10), 1550 => to_unsigned(348, 10), 1551 => to_unsigned(271, 10), 1552 => to_unsigned(360, 10), 1553 => to_unsigned(931, 10), 1554 => to_unsigned(980, 10), 1555 => to_unsigned(1004, 10), 1556 => to_unsigned(659, 10), 1557 => to_unsigned(623, 10), 1558 => to_unsigned(790, 10), 1559 => to_unsigned(831, 10), 1560 => to_unsigned(397, 10), 1561 => to_unsigned(381, 10), 1562 => to_unsigned(140, 10), 1563 => to_unsigned(451, 10), 1564 => to_unsigned(1, 10), 1565 => to_unsigned(471, 10), 1566 => to_unsigned(964, 10), 1567 => to_unsigned(896, 10), 1568 => to_unsigned(585, 10), 1569 => to_unsigned(725, 10), 1570 => to_unsigned(402, 10), 1571 => to_unsigned(28, 10), 1572 => to_unsigned(412, 10), 1573 => to_unsigned(144, 10), 1574 => to_unsigned(601, 10), 1575 => to_unsigned(134, 10), 1576 => to_unsigned(683, 10), 1577 => to_unsigned(718, 10), 1578 => to_unsigned(932, 10), 1579 => to_unsigned(716, 10), 1580 => to_unsigned(109, 10), 1581 => to_unsigned(392, 10), 1582 => to_unsigned(904, 10), 1583 => to_unsigned(685, 10), 1584 => to_unsigned(50, 10), 1585 => to_unsigned(44, 10), 1586 => to_unsigned(36, 10), 1587 => to_unsigned(923, 10), 1588 => to_unsigned(281, 10), 1589 => to_unsigned(196, 10), 1590 => to_unsigned(696, 10), 1591 => to_unsigned(925, 10), 1592 => to_unsigned(286, 10), 1593 => to_unsigned(293, 10), 1594 => to_unsigned(101, 10), 1595 => to_unsigned(204, 10), 1596 => to_unsigned(65, 10), 1597 => to_unsigned(550, 10), 1598 => to_unsigned(398, 10), 1599 => to_unsigned(38, 10), 1600 => to_unsigned(1002, 10), 1601 => to_unsigned(909, 10), 1602 => to_unsigned(677, 10), 1603 => to_unsigned(733, 10), 1604 => to_unsigned(222, 10), 1605 => to_unsigned(295, 10), 1606 => to_unsigned(507, 10), 1607 => to_unsigned(11, 10), 1608 => to_unsigned(255, 10), 1609 => to_unsigned(33, 10), 1610 => to_unsigned(955, 10), 1611 => to_unsigned(373, 10), 1612 => to_unsigned(828, 10), 1613 => to_unsigned(175, 10), 1614 => to_unsigned(632, 10), 1615 => to_unsigned(295, 10), 1616 => to_unsigned(111, 10), 1617 => to_unsigned(495, 10), 1618 => to_unsigned(489, 10), 1619 => to_unsigned(23, 10), 1620 => to_unsigned(0, 10), 1621 => to_unsigned(368, 10), 1622 => to_unsigned(117, 10), 1623 => to_unsigned(122, 10), 1624 => to_unsigned(1014, 10), 1625 => to_unsigned(770, 10), 1626 => to_unsigned(43, 10), 1627 => to_unsigned(335, 10), 1628 => to_unsigned(774, 10), 1629 => to_unsigned(201, 10), 1630 => to_unsigned(893, 10), 1631 => to_unsigned(524, 10), 1632 => to_unsigned(567, 10), 1633 => to_unsigned(943, 10), 1634 => to_unsigned(738, 10), 1635 => to_unsigned(835, 10), 1636 => to_unsigned(969, 10), 1637 => to_unsigned(282, 10), 1638 => to_unsigned(431, 10), 1639 => to_unsigned(497, 10), 1640 => to_unsigned(343, 10), 1641 => to_unsigned(877, 10), 1642 => to_unsigned(958, 10), 1643 => to_unsigned(784, 10), 1644 => to_unsigned(652, 10), 1645 => to_unsigned(76, 10), 1646 => to_unsigned(312, 10), 1647 => to_unsigned(734, 10), 1648 => to_unsigned(556, 10), 1649 => to_unsigned(400, 10), 1650 => to_unsigned(698, 10), 1651 => to_unsigned(288, 10), 1652 => to_unsigned(569, 10), 1653 => to_unsigned(487, 10), 1654 => to_unsigned(322, 10), 1655 => to_unsigned(135, 10), 1656 => to_unsigned(680, 10), 1657 => to_unsigned(228, 10), 1658 => to_unsigned(440, 10), 1659 => to_unsigned(34, 10), 1660 => to_unsigned(902, 10), 1661 => to_unsigned(882, 10), 1662 => to_unsigned(502, 10), 1663 => to_unsigned(717, 10), 1664 => to_unsigned(559, 10), 1665 => to_unsigned(371, 10), 1666 => to_unsigned(630, 10), 1667 => to_unsigned(486, 10), 1668 => to_unsigned(696, 10), 1669 => to_unsigned(775, 10), 1670 => to_unsigned(618, 10), 1671 => to_unsigned(174, 10), 1672 => to_unsigned(435, 10), 1673 => to_unsigned(913, 10), 1674 => to_unsigned(16, 10), 1675 => to_unsigned(928, 10), 1676 => to_unsigned(918, 10), 1677 => to_unsigned(277, 10), 1678 => to_unsigned(972, 10), 1679 => to_unsigned(429, 10), 1680 => to_unsigned(530, 10), 1681 => to_unsigned(656, 10), 1682 => to_unsigned(553, 10), 1683 => to_unsigned(831, 10), 1684 => to_unsigned(68, 10), 1685 => to_unsigned(481, 10), 1686 => to_unsigned(831, 10), 1687 => to_unsigned(879, 10), 1688 => to_unsigned(166, 10), 1689 => to_unsigned(235, 10), 1690 => to_unsigned(742, 10), 1691 => to_unsigned(10, 10), 1692 => to_unsigned(391, 10), 1693 => to_unsigned(598, 10), 1694 => to_unsigned(966, 10), 1695 => to_unsigned(798, 10), 1696 => to_unsigned(470, 10), 1697 => to_unsigned(308, 10), 1698 => to_unsigned(690, 10), 1699 => to_unsigned(322, 10), 1700 => to_unsigned(12, 10), 1701 => to_unsigned(285, 10), 1702 => to_unsigned(571, 10), 1703 => to_unsigned(610, 10), 1704 => to_unsigned(275, 10), 1705 => to_unsigned(280, 10), 1706 => to_unsigned(717, 10), 1707 => to_unsigned(573, 10), 1708 => to_unsigned(729, 10), 1709 => to_unsigned(852, 10), 1710 => to_unsigned(372, 10), 1711 => to_unsigned(759, 10), 1712 => to_unsigned(276, 10), 1713 => to_unsigned(572, 10), 1714 => to_unsigned(568, 10), 1715 => to_unsigned(425, 10), 1716 => to_unsigned(929, 10), 1717 => to_unsigned(798, 10), 1718 => to_unsigned(751, 10), 1719 => to_unsigned(523, 10), 1720 => to_unsigned(999, 10), 1721 => to_unsigned(665, 10), 1722 => to_unsigned(22, 10), 1723 => to_unsigned(437, 10), 1724 => to_unsigned(956, 10), 1725 => to_unsigned(335, 10), 1726 => to_unsigned(185, 10), 1727 => to_unsigned(640, 10), 1728 => to_unsigned(197, 10), 1729 => to_unsigned(629, 10), 1730 => to_unsigned(234, 10), 1731 => to_unsigned(549, 10), 1732 => to_unsigned(296, 10), 1733 => to_unsigned(170, 10), 1734 => to_unsigned(636, 10), 1735 => to_unsigned(950, 10), 1736 => to_unsigned(770, 10), 1737 => to_unsigned(680, 10), 1738 => to_unsigned(760, 10), 1739 => to_unsigned(708, 10), 1740 => to_unsigned(126, 10), 1741 => to_unsigned(57, 10), 1742 => to_unsigned(41, 10), 1743 => to_unsigned(715, 10), 1744 => to_unsigned(497, 10), 1745 => to_unsigned(182, 10), 1746 => to_unsigned(164, 10), 1747 => to_unsigned(796, 10), 1748 => to_unsigned(948, 10), 1749 => to_unsigned(353, 10), 1750 => to_unsigned(521, 10), 1751 => to_unsigned(127, 10), 1752 => to_unsigned(771, 10), 1753 => to_unsigned(606, 10), 1754 => to_unsigned(971, 10), 1755 => to_unsigned(861, 10), 1756 => to_unsigned(550, 10), 1757 => to_unsigned(623, 10), 1758 => to_unsigned(784, 10), 1759 => to_unsigned(622, 10), 1760 => to_unsigned(272, 10), 1761 => to_unsigned(671, 10), 1762 => to_unsigned(569, 10), 1763 => to_unsigned(299, 10), 1764 => to_unsigned(811, 10), 1765 => to_unsigned(385, 10), 1766 => to_unsigned(305, 10), 1767 => to_unsigned(207, 10), 1768 => to_unsigned(837, 10), 1769 => to_unsigned(305, 10), 1770 => to_unsigned(955, 10), 1771 => to_unsigned(517, 10), 1772 => to_unsigned(2, 10), 1773 => to_unsigned(480, 10), 1774 => to_unsigned(2, 10), 1775 => to_unsigned(785, 10), 1776 => to_unsigned(710, 10), 1777 => to_unsigned(671, 10), 1778 => to_unsigned(776, 10), 1779 => to_unsigned(89, 10), 1780 => to_unsigned(887, 10), 1781 => to_unsigned(90, 10), 1782 => to_unsigned(422, 10), 1783 => to_unsigned(257, 10), 1784 => to_unsigned(956, 10), 1785 => to_unsigned(791, 10), 1786 => to_unsigned(620, 10), 1787 => to_unsigned(783, 10), 1788 => to_unsigned(583, 10), 1789 => to_unsigned(507, 10), 1790 => to_unsigned(714, 10), 1791 => to_unsigned(180, 10), 1792 => to_unsigned(443, 10), 1793 => to_unsigned(171, 10), 1794 => to_unsigned(364, 10), 1795 => to_unsigned(37, 10), 1796 => to_unsigned(459, 10), 1797 => to_unsigned(873, 10), 1798 => to_unsigned(197, 10), 1799 => to_unsigned(378, 10), 1800 => to_unsigned(176, 10), 1801 => to_unsigned(991, 10), 1802 => to_unsigned(800, 10), 1803 => to_unsigned(849, 10), 1804 => to_unsigned(100, 10), 1805 => to_unsigned(459, 10), 1806 => to_unsigned(345, 10), 1807 => to_unsigned(119, 10), 1808 => to_unsigned(138, 10), 1809 => to_unsigned(819, 10), 1810 => to_unsigned(336, 10), 1811 => to_unsigned(78, 10), 1812 => to_unsigned(814, 10), 1813 => to_unsigned(162, 10), 1814 => to_unsigned(892, 10), 1815 => to_unsigned(192, 10), 1816 => to_unsigned(360, 10), 1817 => to_unsigned(398, 10), 1818 => to_unsigned(540, 10), 1819 => to_unsigned(94, 10), 1820 => to_unsigned(284, 10), 1821 => to_unsigned(625, 10), 1822 => to_unsigned(575, 10), 1823 => to_unsigned(364, 10), 1824 => to_unsigned(585, 10), 1825 => to_unsigned(411, 10), 1826 => to_unsigned(153, 10), 1827 => to_unsigned(92, 10), 1828 => to_unsigned(636, 10), 1829 => to_unsigned(381, 10), 1830 => to_unsigned(948, 10), 1831 => to_unsigned(885, 10), 1832 => to_unsigned(222, 10), 1833 => to_unsigned(334, 10), 1834 => to_unsigned(586, 10), 1835 => to_unsigned(817, 10), 1836 => to_unsigned(768, 10), 1837 => to_unsigned(555, 10), 1838 => to_unsigned(535, 10), 1839 => to_unsigned(352, 10), 1840 => to_unsigned(1019, 10), 1841 => to_unsigned(498, 10), 1842 => to_unsigned(355, 10), 1843 => to_unsigned(99, 10), 1844 => to_unsigned(246, 10), 1845 => to_unsigned(225, 10), 1846 => to_unsigned(383, 10), 1847 => to_unsigned(342, 10), 1848 => to_unsigned(920, 10), 1849 => to_unsigned(898, 10), 1850 => to_unsigned(693, 10), 1851 => to_unsigned(855, 10), 1852 => to_unsigned(525, 10), 1853 => to_unsigned(828, 10), 1854 => to_unsigned(515, 10), 1855 => to_unsigned(679, 10), 1856 => to_unsigned(903, 10), 1857 => to_unsigned(558, 10), 1858 => to_unsigned(613, 10), 1859 => to_unsigned(150, 10), 1860 => to_unsigned(200, 10), 1861 => to_unsigned(900, 10), 1862 => to_unsigned(546, 10), 1863 => to_unsigned(703, 10), 1864 => to_unsigned(391, 10), 1865 => to_unsigned(691, 10), 1866 => to_unsigned(278, 10), 1867 => to_unsigned(945, 10), 1868 => to_unsigned(547, 10), 1869 => to_unsigned(196, 10), 1870 => to_unsigned(324, 10), 1871 => to_unsigned(793, 10), 1872 => to_unsigned(620, 10), 1873 => to_unsigned(481, 10), 1874 => to_unsigned(501, 10), 1875 => to_unsigned(964, 10), 1876 => to_unsigned(381, 10), 1877 => to_unsigned(521, 10), 1878 => to_unsigned(157, 10), 1879 => to_unsigned(868, 10), 1880 => to_unsigned(931, 10), 1881 => to_unsigned(182, 10), 1882 => to_unsigned(27, 10), 1883 => to_unsigned(513, 10), 1884 => to_unsigned(406, 10), 1885 => to_unsigned(712, 10), 1886 => to_unsigned(830, 10), 1887 => to_unsigned(488, 10), 1888 => to_unsigned(616, 10), 1889 => to_unsigned(696, 10), 1890 => to_unsigned(338, 10), 1891 => to_unsigned(623, 10), 1892 => to_unsigned(33, 10), 1893 => to_unsigned(17, 10), 1894 => to_unsigned(758, 10), 1895 => to_unsigned(757, 10), 1896 => to_unsigned(1001, 10), 1897 => to_unsigned(294, 10), 1898 => to_unsigned(236, 10), 1899 => to_unsigned(316, 10), 1900 => to_unsigned(1012, 10), 1901 => to_unsigned(181, 10), 1902 => to_unsigned(590, 10), 1903 => to_unsigned(797, 10), 1904 => to_unsigned(319, 10), 1905 => to_unsigned(765, 10), 1906 => to_unsigned(1016, 10), 1907 => to_unsigned(939, 10), 1908 => to_unsigned(581, 10), 1909 => to_unsigned(112, 10), 1910 => to_unsigned(434, 10), 1911 => to_unsigned(425, 10), 1912 => to_unsigned(461, 10), 1913 => to_unsigned(428, 10), 1914 => to_unsigned(566, 10), 1915 => to_unsigned(956, 10), 1916 => to_unsigned(516, 10), 1917 => to_unsigned(538, 10), 1918 => to_unsigned(669, 10), 1919 => to_unsigned(163, 10), 1920 => to_unsigned(858, 10), 1921 => to_unsigned(969, 10), 1922 => to_unsigned(708, 10), 1923 => to_unsigned(358, 10), 1924 => to_unsigned(798, 10), 1925 => to_unsigned(1000, 10), 1926 => to_unsigned(507, 10), 1927 => to_unsigned(765, 10), 1928 => to_unsigned(82, 10), 1929 => to_unsigned(970, 10), 1930 => to_unsigned(597, 10), 1931 => to_unsigned(206, 10), 1932 => to_unsigned(957, 10), 1933 => to_unsigned(176, 10), 1934 => to_unsigned(444, 10), 1935 => to_unsigned(526, 10), 1936 => to_unsigned(356, 10), 1937 => to_unsigned(265, 10), 1938 => to_unsigned(219, 10), 1939 => to_unsigned(660, 10), 1940 => to_unsigned(271, 10), 1941 => to_unsigned(322, 10), 1942 => to_unsigned(147, 10), 1943 => to_unsigned(790, 10), 1944 => to_unsigned(118, 10), 1945 => to_unsigned(384, 10), 1946 => to_unsigned(629, 10), 1947 => to_unsigned(218, 10), 1948 => to_unsigned(836, 10), 1949 => to_unsigned(37, 10), 1950 => to_unsigned(569, 10), 1951 => to_unsigned(246, 10), 1952 => to_unsigned(1007, 10), 1953 => to_unsigned(534, 10), 1954 => to_unsigned(57, 10), 1955 => to_unsigned(683, 10), 1956 => to_unsigned(572, 10), 1957 => to_unsigned(547, 10), 1958 => to_unsigned(460, 10), 1959 => to_unsigned(211, 10), 1960 => to_unsigned(633, 10), 1961 => to_unsigned(599, 10), 1962 => to_unsigned(27, 10), 1963 => to_unsigned(404, 10), 1964 => to_unsigned(171, 10), 1965 => to_unsigned(681, 10), 1966 => to_unsigned(112, 10), 1967 => to_unsigned(895, 10), 1968 => to_unsigned(573, 10), 1969 => to_unsigned(950, 10), 1970 => to_unsigned(310, 10), 1971 => to_unsigned(635, 10), 1972 => to_unsigned(276, 10), 1973 => to_unsigned(880, 10), 1974 => to_unsigned(258, 10), 1975 => to_unsigned(878, 10), 1976 => to_unsigned(249, 10), 1977 => to_unsigned(279, 10), 1978 => to_unsigned(162, 10), 1979 => to_unsigned(442, 10), 1980 => to_unsigned(724, 10), 1981 => to_unsigned(512, 10), 1982 => to_unsigned(139, 10), 1983 => to_unsigned(256, 10), 1984 => to_unsigned(193, 10), 1985 => to_unsigned(83, 10), 1986 => to_unsigned(519, 10), 1987 => to_unsigned(57, 10), 1988 => to_unsigned(827, 10), 1989 => to_unsigned(660, 10), 1990 => to_unsigned(443, 10), 1991 => to_unsigned(442, 10), 1992 => to_unsigned(48, 10), 1993 => to_unsigned(843, 10), 1994 => to_unsigned(375, 10), 1995 => to_unsigned(200, 10), 1996 => to_unsigned(880, 10), 1997 => to_unsigned(804, 10), 1998 => to_unsigned(313, 10), 1999 => to_unsigned(484, 10), 2000 => to_unsigned(928, 10), 2001 => to_unsigned(683, 10), 2002 => to_unsigned(585, 10), 2003 => to_unsigned(821, 10), 2004 => to_unsigned(197, 10), 2005 => to_unsigned(277, 10), 2006 => to_unsigned(902, 10), 2007 => to_unsigned(150, 10), 2008 => to_unsigned(909, 10), 2009 => to_unsigned(877, 10), 2010 => to_unsigned(452, 10), 2011 => to_unsigned(104, 10), 2012 => to_unsigned(807, 10), 2013 => to_unsigned(488, 10), 2014 => to_unsigned(940, 10), 2015 => to_unsigned(404, 10), 2016 => to_unsigned(987, 10), 2017 => to_unsigned(69, 10), 2018 => to_unsigned(1009, 10), 2019 => to_unsigned(863, 10), 2020 => to_unsigned(626, 10), 2021 => to_unsigned(838, 10), 2022 => to_unsigned(329, 10), 2023 => to_unsigned(978, 10), 2024 => to_unsigned(124, 10), 2025 => to_unsigned(216, 10), 2026 => to_unsigned(267, 10), 2027 => to_unsigned(369, 10), 2028 => to_unsigned(82, 10), 2029 => to_unsigned(110, 10), 2030 => to_unsigned(261, 10), 2031 => to_unsigned(673, 10), 2032 => to_unsigned(638, 10), 2033 => to_unsigned(500, 10), 2034 => to_unsigned(681, 10), 2035 => to_unsigned(1021, 10), 2036 => to_unsigned(678, 10), 2037 => to_unsigned(22, 10), 2038 => to_unsigned(900, 10), 2039 => to_unsigned(352, 10), 2040 => to_unsigned(874, 10), 2041 => to_unsigned(293, 10), 2042 => to_unsigned(596, 10), 2043 => to_unsigned(1021, 10), 2044 => to_unsigned(63, 10), 2045 => to_unsigned(774, 10), 2046 => to_unsigned(368, 10), 2047 => to_unsigned(413, 10)),
            8 => (0 => to_unsigned(619, 10), 1 => to_unsigned(159, 10), 2 => to_unsigned(164, 10), 3 => to_unsigned(59, 10), 4 => to_unsigned(547, 10), 5 => to_unsigned(302, 10), 6 => to_unsigned(565, 10), 7 => to_unsigned(765, 10), 8 => to_unsigned(128, 10), 9 => to_unsigned(753, 10), 10 => to_unsigned(847, 10), 11 => to_unsigned(121, 10), 12 => to_unsigned(665, 10), 13 => to_unsigned(931, 10), 14 => to_unsigned(363, 10), 15 => to_unsigned(834, 10), 16 => to_unsigned(836, 10), 17 => to_unsigned(298, 10), 18 => to_unsigned(21, 10), 19 => to_unsigned(399, 10), 20 => to_unsigned(911, 10), 21 => to_unsigned(778, 10), 22 => to_unsigned(436, 10), 23 => to_unsigned(945, 10), 24 => to_unsigned(339, 10), 25 => to_unsigned(582, 10), 26 => to_unsigned(155, 10), 27 => to_unsigned(493, 10), 28 => to_unsigned(851, 10), 29 => to_unsigned(111, 10), 30 => to_unsigned(561, 10), 31 => to_unsigned(93, 10), 32 => to_unsigned(40, 10), 33 => to_unsigned(280, 10), 34 => to_unsigned(583, 10), 35 => to_unsigned(166, 10), 36 => to_unsigned(153, 10), 37 => to_unsigned(236, 10), 38 => to_unsigned(162, 10), 39 => to_unsigned(391, 10), 40 => to_unsigned(786, 10), 41 => to_unsigned(904, 10), 42 => to_unsigned(937, 10), 43 => to_unsigned(726, 10), 44 => to_unsigned(958, 10), 45 => to_unsigned(831, 10), 46 => to_unsigned(523, 10), 47 => to_unsigned(235, 10), 48 => to_unsigned(339, 10), 49 => to_unsigned(334, 10), 50 => to_unsigned(671, 10), 51 => to_unsigned(390, 10), 52 => to_unsigned(40, 10), 53 => to_unsigned(230, 10), 54 => to_unsigned(981, 10), 55 => to_unsigned(377, 10), 56 => to_unsigned(970, 10), 57 => to_unsigned(233, 10), 58 => to_unsigned(51, 10), 59 => to_unsigned(402, 10), 60 => to_unsigned(177, 10), 61 => to_unsigned(827, 10), 62 => to_unsigned(241, 10), 63 => to_unsigned(561, 10), 64 => to_unsigned(468, 10), 65 => to_unsigned(511, 10), 66 => to_unsigned(108, 10), 67 => to_unsigned(229, 10), 68 => to_unsigned(182, 10), 69 => to_unsigned(905, 10), 70 => to_unsigned(889, 10), 71 => to_unsigned(939, 10), 72 => to_unsigned(579, 10), 73 => to_unsigned(441, 10), 74 => to_unsigned(511, 10), 75 => to_unsigned(952, 10), 76 => to_unsigned(643, 10), 77 => to_unsigned(503, 10), 78 => to_unsigned(962, 10), 79 => to_unsigned(257, 10), 80 => to_unsigned(599, 10), 81 => to_unsigned(572, 10), 82 => to_unsigned(671, 10), 83 => to_unsigned(498, 10), 84 => to_unsigned(447, 10), 85 => to_unsigned(567, 10), 86 => to_unsigned(419, 10), 87 => to_unsigned(480, 10), 88 => to_unsigned(372, 10), 89 => to_unsigned(939, 10), 90 => to_unsigned(773, 10), 91 => to_unsigned(166, 10), 92 => to_unsigned(513, 10), 93 => to_unsigned(473, 10), 94 => to_unsigned(617, 10), 95 => to_unsigned(483, 10), 96 => to_unsigned(168, 10), 97 => to_unsigned(801, 10), 98 => to_unsigned(429, 10), 99 => to_unsigned(562, 10), 100 => to_unsigned(719, 10), 101 => to_unsigned(17, 10), 102 => to_unsigned(26, 10), 103 => to_unsigned(843, 10), 104 => to_unsigned(664, 10), 105 => to_unsigned(625, 10), 106 => to_unsigned(116, 10), 107 => to_unsigned(306, 10), 108 => to_unsigned(828, 10), 109 => to_unsigned(264, 10), 110 => to_unsigned(433, 10), 111 => to_unsigned(156, 10), 112 => to_unsigned(301, 10), 113 => to_unsigned(870, 10), 114 => to_unsigned(166, 10), 115 => to_unsigned(272, 10), 116 => to_unsigned(15, 10), 117 => to_unsigned(491, 10), 118 => to_unsigned(882, 10), 119 => to_unsigned(811, 10), 120 => to_unsigned(730, 10), 121 => to_unsigned(37, 10), 122 => to_unsigned(690, 10), 123 => to_unsigned(517, 10), 124 => to_unsigned(643, 10), 125 => to_unsigned(624, 10), 126 => to_unsigned(37, 10), 127 => to_unsigned(727, 10), 128 => to_unsigned(766, 10), 129 => to_unsigned(691, 10), 130 => to_unsigned(639, 10), 131 => to_unsigned(376, 10), 132 => to_unsigned(426, 10), 133 => to_unsigned(776, 10), 134 => to_unsigned(873, 10), 135 => to_unsigned(967, 10), 136 => to_unsigned(699, 10), 137 => to_unsigned(865, 10), 138 => to_unsigned(61, 10), 139 => to_unsigned(633, 10), 140 => to_unsigned(58, 10), 141 => to_unsigned(779, 10), 142 => to_unsigned(112, 10), 143 => to_unsigned(118, 10), 144 => to_unsigned(565, 10), 145 => to_unsigned(847, 10), 146 => to_unsigned(922, 10), 147 => to_unsigned(734, 10), 148 => to_unsigned(669, 10), 149 => to_unsigned(210, 10), 150 => to_unsigned(232, 10), 151 => to_unsigned(105, 10), 152 => to_unsigned(473, 10), 153 => to_unsigned(32, 10), 154 => to_unsigned(136, 10), 155 => to_unsigned(224, 10), 156 => to_unsigned(50, 10), 157 => to_unsigned(765, 10), 158 => to_unsigned(460, 10), 159 => to_unsigned(896, 10), 160 => to_unsigned(24, 10), 161 => to_unsigned(255, 10), 162 => to_unsigned(918, 10), 163 => to_unsigned(477, 10), 164 => to_unsigned(114, 10), 165 => to_unsigned(913, 10), 166 => to_unsigned(444, 10), 167 => to_unsigned(1003, 10), 168 => to_unsigned(312, 10), 169 => to_unsigned(927, 10), 170 => to_unsigned(464, 10), 171 => to_unsigned(471, 10), 172 => to_unsigned(738, 10), 173 => to_unsigned(217, 10), 174 => to_unsigned(729, 10), 175 => to_unsigned(840, 10), 176 => to_unsigned(794, 10), 177 => to_unsigned(71, 10), 178 => to_unsigned(979, 10), 179 => to_unsigned(612, 10), 180 => to_unsigned(883, 10), 181 => to_unsigned(891, 10), 182 => to_unsigned(729, 10), 183 => to_unsigned(291, 10), 184 => to_unsigned(117, 10), 185 => to_unsigned(973, 10), 186 => to_unsigned(530, 10), 187 => to_unsigned(889, 10), 188 => to_unsigned(346, 10), 189 => to_unsigned(679, 10), 190 => to_unsigned(243, 10), 191 => to_unsigned(690, 10), 192 => to_unsigned(973, 10), 193 => to_unsigned(258, 10), 194 => to_unsigned(723, 10), 195 => to_unsigned(589, 10), 196 => to_unsigned(980, 10), 197 => to_unsigned(172, 10), 198 => to_unsigned(681, 10), 199 => to_unsigned(47, 10), 200 => to_unsigned(196, 10), 201 => to_unsigned(339, 10), 202 => to_unsigned(185, 10), 203 => to_unsigned(554, 10), 204 => to_unsigned(545, 10), 205 => to_unsigned(619, 10), 206 => to_unsigned(570, 10), 207 => to_unsigned(529, 10), 208 => to_unsigned(237, 10), 209 => to_unsigned(615, 10), 210 => to_unsigned(193, 10), 211 => to_unsigned(481, 10), 212 => to_unsigned(324, 10), 213 => to_unsigned(1006, 10), 214 => to_unsigned(334, 10), 215 => to_unsigned(579, 10), 216 => to_unsigned(396, 10), 217 => to_unsigned(959, 10), 218 => to_unsigned(818, 10), 219 => to_unsigned(968, 10), 220 => to_unsigned(5, 10), 221 => to_unsigned(121, 10), 222 => to_unsigned(479, 10), 223 => to_unsigned(38, 10), 224 => to_unsigned(148, 10), 225 => to_unsigned(507, 10), 226 => to_unsigned(171, 10), 227 => to_unsigned(286, 10), 228 => to_unsigned(755, 10), 229 => to_unsigned(850, 10), 230 => to_unsigned(753, 10), 231 => to_unsigned(325, 10), 232 => to_unsigned(505, 10), 233 => to_unsigned(478, 10), 234 => to_unsigned(527, 10), 235 => to_unsigned(45, 10), 236 => to_unsigned(852, 10), 237 => to_unsigned(742, 10), 238 => to_unsigned(370, 10), 239 => to_unsigned(424, 10), 240 => to_unsigned(794, 10), 241 => to_unsigned(947, 10), 242 => to_unsigned(507, 10), 243 => to_unsigned(818, 10), 244 => to_unsigned(61, 10), 245 => to_unsigned(561, 10), 246 => to_unsigned(479, 10), 247 => to_unsigned(575, 10), 248 => to_unsigned(836, 10), 249 => to_unsigned(244, 10), 250 => to_unsigned(658, 10), 251 => to_unsigned(596, 10), 252 => to_unsigned(112, 10), 253 => to_unsigned(413, 10), 254 => to_unsigned(606, 10), 255 => to_unsigned(204, 10), 256 => to_unsigned(219, 10), 257 => to_unsigned(597, 10), 258 => to_unsigned(572, 10), 259 => to_unsigned(306, 10), 260 => to_unsigned(208, 10), 261 => to_unsigned(626, 10), 262 => to_unsigned(178, 10), 263 => to_unsigned(191, 10), 264 => to_unsigned(329, 10), 265 => to_unsigned(331, 10), 266 => to_unsigned(870, 10), 267 => to_unsigned(932, 10), 268 => to_unsigned(511, 10), 269 => to_unsigned(555, 10), 270 => to_unsigned(374, 10), 271 => to_unsigned(599, 10), 272 => to_unsigned(770, 10), 273 => to_unsigned(126, 10), 274 => to_unsigned(201, 10), 275 => to_unsigned(217, 10), 276 => to_unsigned(872, 10), 277 => to_unsigned(872, 10), 278 => to_unsigned(733, 10), 279 => to_unsigned(221, 10), 280 => to_unsigned(557, 10), 281 => to_unsigned(89, 10), 282 => to_unsigned(298, 10), 283 => to_unsigned(903, 10), 284 => to_unsigned(441, 10), 285 => to_unsigned(569, 10), 286 => to_unsigned(678, 10), 287 => to_unsigned(763, 10), 288 => to_unsigned(484, 10), 289 => to_unsigned(955, 10), 290 => to_unsigned(582, 10), 291 => to_unsigned(529, 10), 292 => to_unsigned(813, 10), 293 => to_unsigned(378, 10), 294 => to_unsigned(331, 10), 295 => to_unsigned(370, 10), 296 => to_unsigned(511, 10), 297 => to_unsigned(330, 10), 298 => to_unsigned(882, 10), 299 => to_unsigned(1001, 10), 300 => to_unsigned(651, 10), 301 => to_unsigned(143, 10), 302 => to_unsigned(209, 10), 303 => to_unsigned(684, 10), 304 => to_unsigned(855, 10), 305 => to_unsigned(446, 10), 306 => to_unsigned(289, 10), 307 => to_unsigned(905, 10), 308 => to_unsigned(456, 10), 309 => to_unsigned(276, 10), 310 => to_unsigned(623, 10), 311 => to_unsigned(812, 10), 312 => to_unsigned(125, 10), 313 => to_unsigned(60, 10), 314 => to_unsigned(77, 10), 315 => to_unsigned(427, 10), 316 => to_unsigned(598, 10), 317 => to_unsigned(122, 10), 318 => to_unsigned(1007, 10), 319 => to_unsigned(693, 10), 320 => to_unsigned(31, 10), 321 => to_unsigned(358, 10), 322 => to_unsigned(648, 10), 323 => to_unsigned(935, 10), 324 => to_unsigned(270, 10), 325 => to_unsigned(317, 10), 326 => to_unsigned(455, 10), 327 => to_unsigned(658, 10), 328 => to_unsigned(93, 10), 329 => to_unsigned(521, 10), 330 => to_unsigned(386, 10), 331 => to_unsigned(214, 10), 332 => to_unsigned(922, 10), 333 => to_unsigned(786, 10), 334 => to_unsigned(200, 10), 335 => to_unsigned(788, 10), 336 => to_unsigned(448, 10), 337 => to_unsigned(763, 10), 338 => to_unsigned(694, 10), 339 => to_unsigned(778, 10), 340 => to_unsigned(678, 10), 341 => to_unsigned(94, 10), 342 => to_unsigned(948, 10), 343 => to_unsigned(676, 10), 344 => to_unsigned(698, 10), 345 => to_unsigned(112, 10), 346 => to_unsigned(493, 10), 347 => to_unsigned(279, 10), 348 => to_unsigned(573, 10), 349 => to_unsigned(445, 10), 350 => to_unsigned(989, 10), 351 => to_unsigned(158, 10), 352 => to_unsigned(434, 10), 353 => to_unsigned(193, 10), 354 => to_unsigned(27, 10), 355 => to_unsigned(408, 10), 356 => to_unsigned(46, 10), 357 => to_unsigned(804, 10), 358 => to_unsigned(179, 10), 359 => to_unsigned(293, 10), 360 => to_unsigned(664, 10), 361 => to_unsigned(585, 10), 362 => to_unsigned(579, 10), 363 => to_unsigned(201, 10), 364 => to_unsigned(526, 10), 365 => to_unsigned(927, 10), 366 => to_unsigned(948, 10), 367 => to_unsigned(379, 10), 368 => to_unsigned(751, 10), 369 => to_unsigned(69, 10), 370 => to_unsigned(547, 10), 371 => to_unsigned(90, 10), 372 => to_unsigned(684, 10), 373 => to_unsigned(589, 10), 374 => to_unsigned(212, 10), 375 => to_unsigned(474, 10), 376 => to_unsigned(288, 10), 377 => to_unsigned(689, 10), 378 => to_unsigned(117, 10), 379 => to_unsigned(823, 10), 380 => to_unsigned(426, 10), 381 => to_unsigned(623, 10), 382 => to_unsigned(98, 10), 383 => to_unsigned(463, 10), 384 => to_unsigned(212, 10), 385 => to_unsigned(223, 10), 386 => to_unsigned(259, 10), 387 => to_unsigned(785, 10), 388 => to_unsigned(152, 10), 389 => to_unsigned(377, 10), 390 => to_unsigned(739, 10), 391 => to_unsigned(454, 10), 392 => to_unsigned(612, 10), 393 => to_unsigned(308, 10), 394 => to_unsigned(109, 10), 395 => to_unsigned(981, 10), 396 => to_unsigned(898, 10), 397 => to_unsigned(419, 10), 398 => to_unsigned(273, 10), 399 => to_unsigned(141, 10), 400 => to_unsigned(785, 10), 401 => to_unsigned(504, 10), 402 => to_unsigned(100, 10), 403 => to_unsigned(819, 10), 404 => to_unsigned(311, 10), 405 => to_unsigned(517, 10), 406 => to_unsigned(997, 10), 407 => to_unsigned(462, 10), 408 => to_unsigned(234, 10), 409 => to_unsigned(804, 10), 410 => to_unsigned(655, 10), 411 => to_unsigned(582, 10), 412 => to_unsigned(454, 10), 413 => to_unsigned(634, 10), 414 => to_unsigned(900, 10), 415 => to_unsigned(899, 10), 416 => to_unsigned(238, 10), 417 => to_unsigned(429, 10), 418 => to_unsigned(956, 10), 419 => to_unsigned(30, 10), 420 => to_unsigned(943, 10), 421 => to_unsigned(289, 10), 422 => to_unsigned(476, 10), 423 => to_unsigned(825, 10), 424 => to_unsigned(575, 10), 425 => to_unsigned(831, 10), 426 => to_unsigned(855, 10), 427 => to_unsigned(54, 10), 428 => to_unsigned(766, 10), 429 => to_unsigned(847, 10), 430 => to_unsigned(283, 10), 431 => to_unsigned(753, 10), 432 => to_unsigned(693, 10), 433 => to_unsigned(285, 10), 434 => to_unsigned(798, 10), 435 => to_unsigned(655, 10), 436 => to_unsigned(252, 10), 437 => to_unsigned(87, 10), 438 => to_unsigned(942, 10), 439 => to_unsigned(368, 10), 440 => to_unsigned(159, 10), 441 => to_unsigned(677, 10), 442 => to_unsigned(864, 10), 443 => to_unsigned(767, 10), 444 => to_unsigned(986, 10), 445 => to_unsigned(722, 10), 446 => to_unsigned(612, 10), 447 => to_unsigned(565, 10), 448 => to_unsigned(789, 10), 449 => to_unsigned(731, 10), 450 => to_unsigned(462, 10), 451 => to_unsigned(257, 10), 452 => to_unsigned(227, 10), 453 => to_unsigned(591, 10), 454 => to_unsigned(57, 10), 455 => to_unsigned(351, 10), 456 => to_unsigned(918, 10), 457 => to_unsigned(803, 10), 458 => to_unsigned(861, 10), 459 => to_unsigned(643, 10), 460 => to_unsigned(435, 10), 461 => to_unsigned(379, 10), 462 => to_unsigned(54, 10), 463 => to_unsigned(160, 10), 464 => to_unsigned(759, 10), 465 => to_unsigned(949, 10), 466 => to_unsigned(360, 10), 467 => to_unsigned(601, 10), 468 => to_unsigned(319, 10), 469 => to_unsigned(754, 10), 470 => to_unsigned(277, 10), 471 => to_unsigned(627, 10), 472 => to_unsigned(308, 10), 473 => to_unsigned(130, 10), 474 => to_unsigned(907, 10), 475 => to_unsigned(750, 10), 476 => to_unsigned(965, 10), 477 => to_unsigned(510, 10), 478 => to_unsigned(31, 10), 479 => to_unsigned(746, 10), 480 => to_unsigned(1011, 10), 481 => to_unsigned(669, 10), 482 => to_unsigned(445, 10), 483 => to_unsigned(250, 10), 484 => to_unsigned(902, 10), 485 => to_unsigned(677, 10), 486 => to_unsigned(0, 10), 487 => to_unsigned(263, 10), 488 => to_unsigned(670, 10), 489 => to_unsigned(969, 10), 490 => to_unsigned(866, 10), 491 => to_unsigned(695, 10), 492 => to_unsigned(980, 10), 493 => to_unsigned(721, 10), 494 => to_unsigned(380, 10), 495 => to_unsigned(789, 10), 496 => to_unsigned(665, 10), 497 => to_unsigned(790, 10), 498 => to_unsigned(940, 10), 499 => to_unsigned(265, 10), 500 => to_unsigned(237, 10), 501 => to_unsigned(1003, 10), 502 => to_unsigned(790, 10), 503 => to_unsigned(437, 10), 504 => to_unsigned(633, 10), 505 => to_unsigned(638, 10), 506 => to_unsigned(292, 10), 507 => to_unsigned(472, 10), 508 => to_unsigned(826, 10), 509 => to_unsigned(896, 10), 510 => to_unsigned(345, 10), 511 => to_unsigned(712, 10), 512 => to_unsigned(694, 10), 513 => to_unsigned(527, 10), 514 => to_unsigned(864, 10), 515 => to_unsigned(496, 10), 516 => to_unsigned(203, 10), 517 => to_unsigned(622, 10), 518 => to_unsigned(764, 10), 519 => to_unsigned(974, 10), 520 => to_unsigned(444, 10), 521 => to_unsigned(743, 10), 522 => to_unsigned(682, 10), 523 => to_unsigned(880, 10), 524 => to_unsigned(422, 10), 525 => to_unsigned(686, 10), 526 => to_unsigned(365, 10), 527 => to_unsigned(80, 10), 528 => to_unsigned(722, 10), 529 => to_unsigned(573, 10), 530 => to_unsigned(540, 10), 531 => to_unsigned(704, 10), 532 => to_unsigned(736, 10), 533 => to_unsigned(194, 10), 534 => to_unsigned(48, 10), 535 => to_unsigned(575, 10), 536 => to_unsigned(914, 10), 537 => to_unsigned(485, 10), 538 => to_unsigned(687, 10), 539 => to_unsigned(208, 10), 540 => to_unsigned(933, 10), 541 => to_unsigned(90, 10), 542 => to_unsigned(646, 10), 543 => to_unsigned(179, 10), 544 => to_unsigned(587, 10), 545 => to_unsigned(641, 10), 546 => to_unsigned(755, 10), 547 => to_unsigned(897, 10), 548 => to_unsigned(25, 10), 549 => to_unsigned(492, 10), 550 => to_unsigned(701, 10), 551 => to_unsigned(573, 10), 552 => to_unsigned(340, 10), 553 => to_unsigned(358, 10), 554 => to_unsigned(588, 10), 555 => to_unsigned(581, 10), 556 => to_unsigned(742, 10), 557 => to_unsigned(947, 10), 558 => to_unsigned(338, 10), 559 => to_unsigned(920, 10), 560 => to_unsigned(995, 10), 561 => to_unsigned(420, 10), 562 => to_unsigned(680, 10), 563 => to_unsigned(845, 10), 564 => to_unsigned(686, 10), 565 => to_unsigned(676, 10), 566 => to_unsigned(155, 10), 567 => to_unsigned(659, 10), 568 => to_unsigned(449, 10), 569 => to_unsigned(485, 10), 570 => to_unsigned(295, 10), 571 => to_unsigned(246, 10), 572 => to_unsigned(542, 10), 573 => to_unsigned(219, 10), 574 => to_unsigned(38, 10), 575 => to_unsigned(496, 10), 576 => to_unsigned(758, 10), 577 => to_unsigned(754, 10), 578 => to_unsigned(74, 10), 579 => to_unsigned(305, 10), 580 => to_unsigned(771, 10), 581 => to_unsigned(469, 10), 582 => to_unsigned(514, 10), 583 => to_unsigned(933, 10), 584 => to_unsigned(132, 10), 585 => to_unsigned(169, 10), 586 => to_unsigned(580, 10), 587 => to_unsigned(285, 10), 588 => to_unsigned(189, 10), 589 => to_unsigned(477, 10), 590 => to_unsigned(540, 10), 591 => to_unsigned(332, 10), 592 => to_unsigned(19, 10), 593 => to_unsigned(649, 10), 594 => to_unsigned(461, 10), 595 => to_unsigned(52, 10), 596 => to_unsigned(470, 10), 597 => to_unsigned(294, 10), 598 => to_unsigned(804, 10), 599 => to_unsigned(27, 10), 600 => to_unsigned(814, 10), 601 => to_unsigned(729, 10), 602 => to_unsigned(591, 10), 603 => to_unsigned(73, 10), 604 => to_unsigned(615, 10), 605 => to_unsigned(800, 10), 606 => to_unsigned(324, 10), 607 => to_unsigned(514, 10), 608 => to_unsigned(675, 10), 609 => to_unsigned(913, 10), 610 => to_unsigned(138, 10), 611 => to_unsigned(638, 10), 612 => to_unsigned(959, 10), 613 => to_unsigned(456, 10), 614 => to_unsigned(722, 10), 615 => to_unsigned(293, 10), 616 => to_unsigned(1006, 10), 617 => to_unsigned(459, 10), 618 => to_unsigned(415, 10), 619 => to_unsigned(1013, 10), 620 => to_unsigned(613, 10), 621 => to_unsigned(993, 10), 622 => to_unsigned(976, 10), 623 => to_unsigned(631, 10), 624 => to_unsigned(942, 10), 625 => to_unsigned(633, 10), 626 => to_unsigned(946, 10), 627 => to_unsigned(931, 10), 628 => to_unsigned(332, 10), 629 => to_unsigned(452, 10), 630 => to_unsigned(997, 10), 631 => to_unsigned(871, 10), 632 => to_unsigned(250, 10), 633 => to_unsigned(737, 10), 634 => to_unsigned(385, 10), 635 => to_unsigned(256, 10), 636 => to_unsigned(262, 10), 637 => to_unsigned(810, 10), 638 => to_unsigned(40, 10), 639 => to_unsigned(669, 10), 640 => to_unsigned(567, 10), 641 => to_unsigned(101, 10), 642 => to_unsigned(897, 10), 643 => to_unsigned(404, 10), 644 => to_unsigned(387, 10), 645 => to_unsigned(198, 10), 646 => to_unsigned(935, 10), 647 => to_unsigned(886, 10), 648 => to_unsigned(141, 10), 649 => to_unsigned(789, 10), 650 => to_unsigned(424, 10), 651 => to_unsigned(616, 10), 652 => to_unsigned(70, 10), 653 => to_unsigned(137, 10), 654 => to_unsigned(489, 10), 655 => to_unsigned(341, 10), 656 => to_unsigned(636, 10), 657 => to_unsigned(1001, 10), 658 => to_unsigned(858, 10), 659 => to_unsigned(283, 10), 660 => to_unsigned(419, 10), 661 => to_unsigned(656, 10), 662 => to_unsigned(421, 10), 663 => to_unsigned(380, 10), 664 => to_unsigned(835, 10), 665 => to_unsigned(1020, 10), 666 => to_unsigned(508, 10), 667 => to_unsigned(328, 10), 668 => to_unsigned(99, 10), 669 => to_unsigned(593, 10), 670 => to_unsigned(380, 10), 671 => to_unsigned(826, 10), 672 => to_unsigned(117, 10), 673 => to_unsigned(582, 10), 674 => to_unsigned(8, 10), 675 => to_unsigned(629, 10), 676 => to_unsigned(996, 10), 677 => to_unsigned(973, 10), 678 => to_unsigned(344, 10), 679 => to_unsigned(760, 10), 680 => to_unsigned(686, 10), 681 => to_unsigned(818, 10), 682 => to_unsigned(997, 10), 683 => to_unsigned(124, 10), 684 => to_unsigned(93, 10), 685 => to_unsigned(499, 10), 686 => to_unsigned(907, 10), 687 => to_unsigned(367, 10), 688 => to_unsigned(540, 10), 689 => to_unsigned(200, 10), 690 => to_unsigned(889, 10), 691 => to_unsigned(751, 10), 692 => to_unsigned(277, 10), 693 => to_unsigned(932, 10), 694 => to_unsigned(296, 10), 695 => to_unsigned(417, 10), 696 => to_unsigned(614, 10), 697 => to_unsigned(60, 10), 698 => to_unsigned(881, 10), 699 => to_unsigned(446, 10), 700 => to_unsigned(131, 10), 701 => to_unsigned(847, 10), 702 => to_unsigned(253, 10), 703 => to_unsigned(164, 10), 704 => to_unsigned(217, 10), 705 => to_unsigned(711, 10), 706 => to_unsigned(594, 10), 707 => to_unsigned(661, 10), 708 => to_unsigned(703, 10), 709 => to_unsigned(126, 10), 710 => to_unsigned(953, 10), 711 => to_unsigned(3, 10), 712 => to_unsigned(47, 10), 713 => to_unsigned(722, 10), 714 => to_unsigned(343, 10), 715 => to_unsigned(612, 10), 716 => to_unsigned(431, 10), 717 => to_unsigned(864, 10), 718 => to_unsigned(919, 10), 719 => to_unsigned(186, 10), 720 => to_unsigned(223, 10), 721 => to_unsigned(493, 10), 722 => to_unsigned(426, 10), 723 => to_unsigned(477, 10), 724 => to_unsigned(720, 10), 725 => to_unsigned(356, 10), 726 => to_unsigned(942, 10), 727 => to_unsigned(452, 10), 728 => to_unsigned(518, 10), 729 => to_unsigned(177, 10), 730 => to_unsigned(725, 10), 731 => to_unsigned(112, 10), 732 => to_unsigned(963, 10), 733 => to_unsigned(131, 10), 734 => to_unsigned(480, 10), 735 => to_unsigned(958, 10), 736 => to_unsigned(465, 10), 737 => to_unsigned(21, 10), 738 => to_unsigned(365, 10), 739 => to_unsigned(134, 10), 740 => to_unsigned(809, 10), 741 => to_unsigned(980, 10), 742 => to_unsigned(860, 10), 743 => to_unsigned(512, 10), 744 => to_unsigned(133, 10), 745 => to_unsigned(562, 10), 746 => to_unsigned(29, 10), 747 => to_unsigned(241, 10), 748 => to_unsigned(67, 10), 749 => to_unsigned(1010, 10), 750 => to_unsigned(988, 10), 751 => to_unsigned(1003, 10), 752 => to_unsigned(568, 10), 753 => to_unsigned(147, 10), 754 => to_unsigned(386, 10), 755 => to_unsigned(970, 10), 756 => to_unsigned(18, 10), 757 => to_unsigned(203, 10), 758 => to_unsigned(562, 10), 759 => to_unsigned(43, 10), 760 => to_unsigned(62, 10), 761 => to_unsigned(640, 10), 762 => to_unsigned(138, 10), 763 => to_unsigned(687, 10), 764 => to_unsigned(912, 10), 765 => to_unsigned(476, 10), 766 => to_unsigned(811, 10), 767 => to_unsigned(908, 10), 768 => to_unsigned(221, 10), 769 => to_unsigned(465, 10), 770 => to_unsigned(906, 10), 771 => to_unsigned(449, 10), 772 => to_unsigned(645, 10), 773 => to_unsigned(679, 10), 774 => to_unsigned(732, 10), 775 => to_unsigned(125, 10), 776 => to_unsigned(648, 10), 777 => to_unsigned(992, 10), 778 => to_unsigned(808, 10), 779 => to_unsigned(527, 10), 780 => to_unsigned(257, 10), 781 => to_unsigned(934, 10), 782 => to_unsigned(929, 10), 783 => to_unsigned(687, 10), 784 => to_unsigned(958, 10), 785 => to_unsigned(367, 10), 786 => to_unsigned(695, 10), 787 => to_unsigned(717, 10), 788 => to_unsigned(811, 10), 789 => to_unsigned(1017, 10), 790 => to_unsigned(670, 10), 791 => to_unsigned(969, 10), 792 => to_unsigned(43, 10), 793 => to_unsigned(500, 10), 794 => to_unsigned(285, 10), 795 => to_unsigned(646, 10), 796 => to_unsigned(19, 10), 797 => to_unsigned(790, 10), 798 => to_unsigned(790, 10), 799 => to_unsigned(680, 10), 800 => to_unsigned(342, 10), 801 => to_unsigned(203, 10), 802 => to_unsigned(1013, 10), 803 => to_unsigned(836, 10), 804 => to_unsigned(270, 10), 805 => to_unsigned(36, 10), 806 => to_unsigned(329, 10), 807 => to_unsigned(525, 10), 808 => to_unsigned(975, 10), 809 => to_unsigned(650, 10), 810 => to_unsigned(343, 10), 811 => to_unsigned(810, 10), 812 => to_unsigned(636, 10), 813 => to_unsigned(723, 10), 814 => to_unsigned(88, 10), 815 => to_unsigned(729, 10), 816 => to_unsigned(938, 10), 817 => to_unsigned(964, 10), 818 => to_unsigned(128, 10), 819 => to_unsigned(956, 10), 820 => to_unsigned(613, 10), 821 => to_unsigned(87, 10), 822 => to_unsigned(638, 10), 823 => to_unsigned(838, 10), 824 => to_unsigned(859, 10), 825 => to_unsigned(246, 10), 826 => to_unsigned(584, 10), 827 => to_unsigned(199, 10), 828 => to_unsigned(45, 10), 829 => to_unsigned(238, 10), 830 => to_unsigned(341, 10), 831 => to_unsigned(138, 10), 832 => to_unsigned(5, 10), 833 => to_unsigned(104, 10), 834 => to_unsigned(149, 10), 835 => to_unsigned(441, 10), 836 => to_unsigned(512, 10), 837 => to_unsigned(380, 10), 838 => to_unsigned(55, 10), 839 => to_unsigned(702, 10), 840 => to_unsigned(493, 10), 841 => to_unsigned(57, 10), 842 => to_unsigned(42, 10), 843 => to_unsigned(73, 10), 844 => to_unsigned(443, 10), 845 => to_unsigned(867, 10), 846 => to_unsigned(340, 10), 847 => to_unsigned(936, 10), 848 => to_unsigned(1, 10), 849 => to_unsigned(608, 10), 850 => to_unsigned(52, 10), 851 => to_unsigned(356, 10), 852 => to_unsigned(124, 10), 853 => to_unsigned(932, 10), 854 => to_unsigned(982, 10), 855 => to_unsigned(593, 10), 856 => to_unsigned(920, 10), 857 => to_unsigned(874, 10), 858 => to_unsigned(43, 10), 859 => to_unsigned(170, 10), 860 => to_unsigned(780, 10), 861 => to_unsigned(807, 10), 862 => to_unsigned(226, 10), 863 => to_unsigned(95, 10), 864 => to_unsigned(255, 10), 865 => to_unsigned(853, 10), 866 => to_unsigned(425, 10), 867 => to_unsigned(832, 10), 868 => to_unsigned(287, 10), 869 => to_unsigned(87, 10), 870 => to_unsigned(861, 10), 871 => to_unsigned(351, 10), 872 => to_unsigned(66, 10), 873 => to_unsigned(677, 10), 874 => to_unsigned(302, 10), 875 => to_unsigned(16, 10), 876 => to_unsigned(831, 10), 877 => to_unsigned(1016, 10), 878 => to_unsigned(970, 10), 879 => to_unsigned(282, 10), 880 => to_unsigned(596, 10), 881 => to_unsigned(917, 10), 882 => to_unsigned(704, 10), 883 => to_unsigned(935, 10), 884 => to_unsigned(514, 10), 885 => to_unsigned(805, 10), 886 => to_unsigned(846, 10), 887 => to_unsigned(602, 10), 888 => to_unsigned(459, 10), 889 => to_unsigned(657, 10), 890 => to_unsigned(772, 10), 891 => to_unsigned(121, 10), 892 => to_unsigned(680, 10), 893 => to_unsigned(898, 10), 894 => to_unsigned(254, 10), 895 => to_unsigned(284, 10), 896 => to_unsigned(640, 10), 897 => to_unsigned(691, 10), 898 => to_unsigned(837, 10), 899 => to_unsigned(435, 10), 900 => to_unsigned(254, 10), 901 => to_unsigned(172, 10), 902 => to_unsigned(287, 10), 903 => to_unsigned(176, 10), 904 => to_unsigned(895, 10), 905 => to_unsigned(570, 10), 906 => to_unsigned(921, 10), 907 => to_unsigned(50, 10), 908 => to_unsigned(535, 10), 909 => to_unsigned(774, 10), 910 => to_unsigned(426, 10), 911 => to_unsigned(815, 10), 912 => to_unsigned(268, 10), 913 => to_unsigned(55, 10), 914 => to_unsigned(553, 10), 915 => to_unsigned(234, 10), 916 => to_unsigned(692, 10), 917 => to_unsigned(42, 10), 918 => to_unsigned(667, 10), 919 => to_unsigned(484, 10), 920 => to_unsigned(44, 10), 921 => to_unsigned(958, 10), 922 => to_unsigned(1015, 10), 923 => to_unsigned(928, 10), 924 => to_unsigned(491, 10), 925 => to_unsigned(726, 10), 926 => to_unsigned(513, 10), 927 => to_unsigned(607, 10), 928 => to_unsigned(840, 10), 929 => to_unsigned(915, 10), 930 => to_unsigned(148, 10), 931 => to_unsigned(830, 10), 932 => to_unsigned(0, 10), 933 => to_unsigned(363, 10), 934 => to_unsigned(183, 10), 935 => to_unsigned(529, 10), 936 => to_unsigned(787, 10), 937 => to_unsigned(709, 10), 938 => to_unsigned(610, 10), 939 => to_unsigned(284, 10), 940 => to_unsigned(954, 10), 941 => to_unsigned(797, 10), 942 => to_unsigned(487, 10), 943 => to_unsigned(77, 10), 944 => to_unsigned(685, 10), 945 => to_unsigned(632, 10), 946 => to_unsigned(863, 10), 947 => to_unsigned(751, 10), 948 => to_unsigned(506, 10), 949 => to_unsigned(695, 10), 950 => to_unsigned(154, 10), 951 => to_unsigned(808, 10), 952 => to_unsigned(666, 10), 953 => to_unsigned(341, 10), 954 => to_unsigned(64, 10), 955 => to_unsigned(80, 10), 956 => to_unsigned(153, 10), 957 => to_unsigned(542, 10), 958 => to_unsigned(218, 10), 959 => to_unsigned(195, 10), 960 => to_unsigned(964, 10), 961 => to_unsigned(389, 10), 962 => to_unsigned(866, 10), 963 => to_unsigned(558, 10), 964 => to_unsigned(456, 10), 965 => to_unsigned(74, 10), 966 => to_unsigned(366, 10), 967 => to_unsigned(674, 10), 968 => to_unsigned(880, 10), 969 => to_unsigned(105, 10), 970 => to_unsigned(370, 10), 971 => to_unsigned(638, 10), 972 => to_unsigned(973, 10), 973 => to_unsigned(316, 10), 974 => to_unsigned(338, 10), 975 => to_unsigned(188, 10), 976 => to_unsigned(970, 10), 977 => to_unsigned(830, 10), 978 => to_unsigned(268, 10), 979 => to_unsigned(745, 10), 980 => to_unsigned(163, 10), 981 => to_unsigned(697, 10), 982 => to_unsigned(8, 10), 983 => to_unsigned(114, 10), 984 => to_unsigned(413, 10), 985 => to_unsigned(182, 10), 986 => to_unsigned(388, 10), 987 => to_unsigned(682, 10), 988 => to_unsigned(221, 10), 989 => to_unsigned(944, 10), 990 => to_unsigned(651, 10), 991 => to_unsigned(55, 10), 992 => to_unsigned(182, 10), 993 => to_unsigned(654, 10), 994 => to_unsigned(738, 10), 995 => to_unsigned(871, 10), 996 => to_unsigned(640, 10), 997 => to_unsigned(104, 10), 998 => to_unsigned(844, 10), 999 => to_unsigned(1021, 10), 1000 => to_unsigned(660, 10), 1001 => to_unsigned(312, 10), 1002 => to_unsigned(29, 10), 1003 => to_unsigned(590, 10), 1004 => to_unsigned(748, 10), 1005 => to_unsigned(150, 10), 1006 => to_unsigned(84, 10), 1007 => to_unsigned(641, 10), 1008 => to_unsigned(431, 10), 1009 => to_unsigned(574, 10), 1010 => to_unsigned(291, 10), 1011 => to_unsigned(377, 10), 1012 => to_unsigned(794, 10), 1013 => to_unsigned(501, 10), 1014 => to_unsigned(53, 10), 1015 => to_unsigned(809, 10), 1016 => to_unsigned(499, 10), 1017 => to_unsigned(843, 10), 1018 => to_unsigned(268, 10), 1019 => to_unsigned(615, 10), 1020 => to_unsigned(717, 10), 1021 => to_unsigned(111, 10), 1022 => to_unsigned(580, 10), 1023 => to_unsigned(899, 10), 1024 => to_unsigned(839, 10), 1025 => to_unsigned(234, 10), 1026 => to_unsigned(843, 10), 1027 => to_unsigned(493, 10), 1028 => to_unsigned(171, 10), 1029 => to_unsigned(200, 10), 1030 => to_unsigned(538, 10), 1031 => to_unsigned(192, 10), 1032 => to_unsigned(647, 10), 1033 => to_unsigned(960, 10), 1034 => to_unsigned(246, 10), 1035 => to_unsigned(132, 10), 1036 => to_unsigned(100, 10), 1037 => to_unsigned(559, 10), 1038 => to_unsigned(478, 10), 1039 => to_unsigned(181, 10), 1040 => to_unsigned(972, 10), 1041 => to_unsigned(14, 10), 1042 => to_unsigned(704, 10), 1043 => to_unsigned(47, 10), 1044 => to_unsigned(465, 10), 1045 => to_unsigned(469, 10), 1046 => to_unsigned(973, 10), 1047 => to_unsigned(766, 10), 1048 => to_unsigned(936, 10), 1049 => to_unsigned(283, 10), 1050 => to_unsigned(379, 10), 1051 => to_unsigned(181, 10), 1052 => to_unsigned(382, 10), 1053 => to_unsigned(952, 10), 1054 => to_unsigned(739, 10), 1055 => to_unsigned(346, 10), 1056 => to_unsigned(278, 10), 1057 => to_unsigned(344, 10), 1058 => to_unsigned(793, 10), 1059 => to_unsigned(411, 10), 1060 => to_unsigned(720, 10), 1061 => to_unsigned(325, 10), 1062 => to_unsigned(337, 10), 1063 => to_unsigned(867, 10), 1064 => to_unsigned(480, 10), 1065 => to_unsigned(119, 10), 1066 => to_unsigned(659, 10), 1067 => to_unsigned(480, 10), 1068 => to_unsigned(157, 10), 1069 => to_unsigned(402, 10), 1070 => to_unsigned(662, 10), 1071 => to_unsigned(496, 10), 1072 => to_unsigned(69, 10), 1073 => to_unsigned(147, 10), 1074 => to_unsigned(733, 10), 1075 => to_unsigned(684, 10), 1076 => to_unsigned(166, 10), 1077 => to_unsigned(107, 10), 1078 => to_unsigned(891, 10), 1079 => to_unsigned(54, 10), 1080 => to_unsigned(455, 10), 1081 => to_unsigned(541, 10), 1082 => to_unsigned(1010, 10), 1083 => to_unsigned(390, 10), 1084 => to_unsigned(394, 10), 1085 => to_unsigned(740, 10), 1086 => to_unsigned(942, 10), 1087 => to_unsigned(631, 10), 1088 => to_unsigned(368, 10), 1089 => to_unsigned(714, 10), 1090 => to_unsigned(853, 10), 1091 => to_unsigned(277, 10), 1092 => to_unsigned(510, 10), 1093 => to_unsigned(995, 10), 1094 => to_unsigned(925, 10), 1095 => to_unsigned(34, 10), 1096 => to_unsigned(156, 10), 1097 => to_unsigned(769, 10), 1098 => to_unsigned(688, 10), 1099 => to_unsigned(825, 10), 1100 => to_unsigned(717, 10), 1101 => to_unsigned(167, 10), 1102 => to_unsigned(61, 10), 1103 => to_unsigned(4, 10), 1104 => to_unsigned(322, 10), 1105 => to_unsigned(585, 10), 1106 => to_unsigned(556, 10), 1107 => to_unsigned(683, 10), 1108 => to_unsigned(594, 10), 1109 => to_unsigned(900, 10), 1110 => to_unsigned(380, 10), 1111 => to_unsigned(744, 10), 1112 => to_unsigned(1008, 10), 1113 => to_unsigned(481, 10), 1114 => to_unsigned(228, 10), 1115 => to_unsigned(122, 10), 1116 => to_unsigned(684, 10), 1117 => to_unsigned(740, 10), 1118 => to_unsigned(947, 10), 1119 => to_unsigned(369, 10), 1120 => to_unsigned(357, 10), 1121 => to_unsigned(614, 10), 1122 => to_unsigned(271, 10), 1123 => to_unsigned(703, 10), 1124 => to_unsigned(689, 10), 1125 => to_unsigned(958, 10), 1126 => to_unsigned(524, 10), 1127 => to_unsigned(168, 10), 1128 => to_unsigned(980, 10), 1129 => to_unsigned(16, 10), 1130 => to_unsigned(849, 10), 1131 => to_unsigned(730, 10), 1132 => to_unsigned(869, 10), 1133 => to_unsigned(174, 10), 1134 => to_unsigned(489, 10), 1135 => to_unsigned(631, 10), 1136 => to_unsigned(556, 10), 1137 => to_unsigned(619, 10), 1138 => to_unsigned(619, 10), 1139 => to_unsigned(431, 10), 1140 => to_unsigned(480, 10), 1141 => to_unsigned(277, 10), 1142 => to_unsigned(624, 10), 1143 => to_unsigned(162, 10), 1144 => to_unsigned(841, 10), 1145 => to_unsigned(253, 10), 1146 => to_unsigned(108, 10), 1147 => to_unsigned(40, 10), 1148 => to_unsigned(797, 10), 1149 => to_unsigned(348, 10), 1150 => to_unsigned(647, 10), 1151 => to_unsigned(727, 10), 1152 => to_unsigned(706, 10), 1153 => to_unsigned(394, 10), 1154 => to_unsigned(537, 10), 1155 => to_unsigned(597, 10), 1156 => to_unsigned(296, 10), 1157 => to_unsigned(518, 10), 1158 => to_unsigned(466, 10), 1159 => to_unsigned(144, 10), 1160 => to_unsigned(139, 10), 1161 => to_unsigned(685, 10), 1162 => to_unsigned(664, 10), 1163 => to_unsigned(790, 10), 1164 => to_unsigned(955, 10), 1165 => to_unsigned(67, 10), 1166 => to_unsigned(1003, 10), 1167 => to_unsigned(94, 10), 1168 => to_unsigned(941, 10), 1169 => to_unsigned(104, 10), 1170 => to_unsigned(775, 10), 1171 => to_unsigned(770, 10), 1172 => to_unsigned(797, 10), 1173 => to_unsigned(968, 10), 1174 => to_unsigned(817, 10), 1175 => to_unsigned(632, 10), 1176 => to_unsigned(925, 10), 1177 => to_unsigned(770, 10), 1178 => to_unsigned(262, 10), 1179 => to_unsigned(446, 10), 1180 => to_unsigned(564, 10), 1181 => to_unsigned(90, 10), 1182 => to_unsigned(769, 10), 1183 => to_unsigned(381, 10), 1184 => to_unsigned(607, 10), 1185 => to_unsigned(744, 10), 1186 => to_unsigned(811, 10), 1187 => to_unsigned(618, 10), 1188 => to_unsigned(317, 10), 1189 => to_unsigned(367, 10), 1190 => to_unsigned(845, 10), 1191 => to_unsigned(430, 10), 1192 => to_unsigned(501, 10), 1193 => to_unsigned(712, 10), 1194 => to_unsigned(837, 10), 1195 => to_unsigned(843, 10), 1196 => to_unsigned(287, 10), 1197 => to_unsigned(546, 10), 1198 => to_unsigned(576, 10), 1199 => to_unsigned(510, 10), 1200 => to_unsigned(268, 10), 1201 => to_unsigned(428, 10), 1202 => to_unsigned(852, 10), 1203 => to_unsigned(372, 10), 1204 => to_unsigned(142, 10), 1205 => to_unsigned(610, 10), 1206 => to_unsigned(29, 10), 1207 => to_unsigned(861, 10), 1208 => to_unsigned(822, 10), 1209 => to_unsigned(285, 10), 1210 => to_unsigned(897, 10), 1211 => to_unsigned(210, 10), 1212 => to_unsigned(539, 10), 1213 => to_unsigned(201, 10), 1214 => to_unsigned(555, 10), 1215 => to_unsigned(500, 10), 1216 => to_unsigned(508, 10), 1217 => to_unsigned(88, 10), 1218 => to_unsigned(360, 10), 1219 => to_unsigned(413, 10), 1220 => to_unsigned(268, 10), 1221 => to_unsigned(161, 10), 1222 => to_unsigned(458, 10), 1223 => to_unsigned(63, 10), 1224 => to_unsigned(945, 10), 1225 => to_unsigned(652, 10), 1226 => to_unsigned(134, 10), 1227 => to_unsigned(454, 10), 1228 => to_unsigned(1018, 10), 1229 => to_unsigned(30, 10), 1230 => to_unsigned(618, 10), 1231 => to_unsigned(581, 10), 1232 => to_unsigned(868, 10), 1233 => to_unsigned(29, 10), 1234 => to_unsigned(538, 10), 1235 => to_unsigned(444, 10), 1236 => to_unsigned(797, 10), 1237 => to_unsigned(18, 10), 1238 => to_unsigned(1020, 10), 1239 => to_unsigned(583, 10), 1240 => to_unsigned(660, 10), 1241 => to_unsigned(600, 10), 1242 => to_unsigned(544, 10), 1243 => to_unsigned(191, 10), 1244 => to_unsigned(734, 10), 1245 => to_unsigned(987, 10), 1246 => to_unsigned(24, 10), 1247 => to_unsigned(252, 10), 1248 => to_unsigned(643, 10), 1249 => to_unsigned(645, 10), 1250 => to_unsigned(397, 10), 1251 => to_unsigned(235, 10), 1252 => to_unsigned(325, 10), 1253 => to_unsigned(401, 10), 1254 => to_unsigned(856, 10), 1255 => to_unsigned(595, 10), 1256 => to_unsigned(432, 10), 1257 => to_unsigned(601, 10), 1258 => to_unsigned(377, 10), 1259 => to_unsigned(132, 10), 1260 => to_unsigned(145, 10), 1261 => to_unsigned(510, 10), 1262 => to_unsigned(545, 10), 1263 => to_unsigned(792, 10), 1264 => to_unsigned(356, 10), 1265 => to_unsigned(740, 10), 1266 => to_unsigned(805, 10), 1267 => to_unsigned(543, 10), 1268 => to_unsigned(212, 10), 1269 => to_unsigned(564, 10), 1270 => to_unsigned(467, 10), 1271 => to_unsigned(658, 10), 1272 => to_unsigned(718, 10), 1273 => to_unsigned(668, 10), 1274 => to_unsigned(882, 10), 1275 => to_unsigned(474, 10), 1276 => to_unsigned(632, 10), 1277 => to_unsigned(378, 10), 1278 => to_unsigned(719, 10), 1279 => to_unsigned(744, 10), 1280 => to_unsigned(1, 10), 1281 => to_unsigned(717, 10), 1282 => to_unsigned(894, 10), 1283 => to_unsigned(542, 10), 1284 => to_unsigned(379, 10), 1285 => to_unsigned(977, 10), 1286 => to_unsigned(308, 10), 1287 => to_unsigned(191, 10), 1288 => to_unsigned(165, 10), 1289 => to_unsigned(678, 10), 1290 => to_unsigned(542, 10), 1291 => to_unsigned(42, 10), 1292 => to_unsigned(1009, 10), 1293 => to_unsigned(356, 10), 1294 => to_unsigned(778, 10), 1295 => to_unsigned(1000, 10), 1296 => to_unsigned(465, 10), 1297 => to_unsigned(814, 10), 1298 => to_unsigned(376, 10), 1299 => to_unsigned(949, 10), 1300 => to_unsigned(503, 10), 1301 => to_unsigned(272, 10), 1302 => to_unsigned(570, 10), 1303 => to_unsigned(916, 10), 1304 => to_unsigned(814, 10), 1305 => to_unsigned(206, 10), 1306 => to_unsigned(992, 10), 1307 => to_unsigned(908, 10), 1308 => to_unsigned(459, 10), 1309 => to_unsigned(132, 10), 1310 => to_unsigned(17, 10), 1311 => to_unsigned(531, 10), 1312 => to_unsigned(558, 10), 1313 => to_unsigned(19, 10), 1314 => to_unsigned(521, 10), 1315 => to_unsigned(264, 10), 1316 => to_unsigned(490, 10), 1317 => to_unsigned(20, 10), 1318 => to_unsigned(615, 10), 1319 => to_unsigned(686, 10), 1320 => to_unsigned(495, 10), 1321 => to_unsigned(122, 10), 1322 => to_unsigned(1008, 10), 1323 => to_unsigned(982, 10), 1324 => to_unsigned(134, 10), 1325 => to_unsigned(115, 10), 1326 => to_unsigned(799, 10), 1327 => to_unsigned(89, 10), 1328 => to_unsigned(230, 10), 1329 => to_unsigned(994, 10), 1330 => to_unsigned(569, 10), 1331 => to_unsigned(713, 10), 1332 => to_unsigned(977, 10), 1333 => to_unsigned(19, 10), 1334 => to_unsigned(916, 10), 1335 => to_unsigned(444, 10), 1336 => to_unsigned(719, 10), 1337 => to_unsigned(269, 10), 1338 => to_unsigned(760, 10), 1339 => to_unsigned(304, 10), 1340 => to_unsigned(195, 10), 1341 => to_unsigned(774, 10), 1342 => to_unsigned(779, 10), 1343 => to_unsigned(122, 10), 1344 => to_unsigned(47, 10), 1345 => to_unsigned(527, 10), 1346 => to_unsigned(79, 10), 1347 => to_unsigned(584, 10), 1348 => to_unsigned(805, 10), 1349 => to_unsigned(818, 10), 1350 => to_unsigned(209, 10), 1351 => to_unsigned(156, 10), 1352 => to_unsigned(470, 10), 1353 => to_unsigned(929, 10), 1354 => to_unsigned(636, 10), 1355 => to_unsigned(941, 10), 1356 => to_unsigned(709, 10), 1357 => to_unsigned(66, 10), 1358 => to_unsigned(855, 10), 1359 => to_unsigned(959, 10), 1360 => to_unsigned(928, 10), 1361 => to_unsigned(468, 10), 1362 => to_unsigned(510, 10), 1363 => to_unsigned(791, 10), 1364 => to_unsigned(270, 10), 1365 => to_unsigned(71, 10), 1366 => to_unsigned(709, 10), 1367 => to_unsigned(1012, 10), 1368 => to_unsigned(179, 10), 1369 => to_unsigned(679, 10), 1370 => to_unsigned(393, 10), 1371 => to_unsigned(34, 10), 1372 => to_unsigned(947, 10), 1373 => to_unsigned(447, 10), 1374 => to_unsigned(634, 10), 1375 => to_unsigned(230, 10), 1376 => to_unsigned(569, 10), 1377 => to_unsigned(991, 10), 1378 => to_unsigned(155, 10), 1379 => to_unsigned(441, 10), 1380 => to_unsigned(600, 10), 1381 => to_unsigned(165, 10), 1382 => to_unsigned(303, 10), 1383 => to_unsigned(758, 10), 1384 => to_unsigned(190, 10), 1385 => to_unsigned(300, 10), 1386 => to_unsigned(19, 10), 1387 => to_unsigned(113, 10), 1388 => to_unsigned(750, 10), 1389 => to_unsigned(884, 10), 1390 => to_unsigned(516, 10), 1391 => to_unsigned(904, 10), 1392 => to_unsigned(944, 10), 1393 => to_unsigned(765, 10), 1394 => to_unsigned(303, 10), 1395 => to_unsigned(628, 10), 1396 => to_unsigned(296, 10), 1397 => to_unsigned(778, 10), 1398 => to_unsigned(546, 10), 1399 => to_unsigned(698, 10), 1400 => to_unsigned(438, 10), 1401 => to_unsigned(45, 10), 1402 => to_unsigned(524, 10), 1403 => to_unsigned(574, 10), 1404 => to_unsigned(258, 10), 1405 => to_unsigned(158, 10), 1406 => to_unsigned(943, 10), 1407 => to_unsigned(967, 10), 1408 => to_unsigned(526, 10), 1409 => to_unsigned(644, 10), 1410 => to_unsigned(75, 10), 1411 => to_unsigned(376, 10), 1412 => to_unsigned(345, 10), 1413 => to_unsigned(761, 10), 1414 => to_unsigned(29, 10), 1415 => to_unsigned(563, 10), 1416 => to_unsigned(528, 10), 1417 => to_unsigned(261, 10), 1418 => to_unsigned(714, 10), 1419 => to_unsigned(638, 10), 1420 => to_unsigned(957, 10), 1421 => to_unsigned(285, 10), 1422 => to_unsigned(521, 10), 1423 => to_unsigned(644, 10), 1424 => to_unsigned(353, 10), 1425 => to_unsigned(750, 10), 1426 => to_unsigned(270, 10), 1427 => to_unsigned(851, 10), 1428 => to_unsigned(602, 10), 1429 => to_unsigned(592, 10), 1430 => to_unsigned(220, 10), 1431 => to_unsigned(368, 10), 1432 => to_unsigned(228, 10), 1433 => to_unsigned(478, 10), 1434 => to_unsigned(457, 10), 1435 => to_unsigned(288, 10), 1436 => to_unsigned(976, 10), 1437 => to_unsigned(280, 10), 1438 => to_unsigned(86, 10), 1439 => to_unsigned(870, 10), 1440 => to_unsigned(463, 10), 1441 => to_unsigned(163, 10), 1442 => to_unsigned(560, 10), 1443 => to_unsigned(656, 10), 1444 => to_unsigned(245, 10), 1445 => to_unsigned(779, 10), 1446 => to_unsigned(52, 10), 1447 => to_unsigned(470, 10), 1448 => to_unsigned(209, 10), 1449 => to_unsigned(566, 10), 1450 => to_unsigned(210, 10), 1451 => to_unsigned(228, 10), 1452 => to_unsigned(734, 10), 1453 => to_unsigned(952, 10), 1454 => to_unsigned(511, 10), 1455 => to_unsigned(761, 10), 1456 => to_unsigned(22, 10), 1457 => to_unsigned(168, 10), 1458 => to_unsigned(912, 10), 1459 => to_unsigned(396, 10), 1460 => to_unsigned(167, 10), 1461 => to_unsigned(278, 10), 1462 => to_unsigned(966, 10), 1463 => to_unsigned(213, 10), 1464 => to_unsigned(994, 10), 1465 => to_unsigned(728, 10), 1466 => to_unsigned(1018, 10), 1467 => to_unsigned(969, 10), 1468 => to_unsigned(887, 10), 1469 => to_unsigned(378, 10), 1470 => to_unsigned(447, 10), 1471 => to_unsigned(579, 10), 1472 => to_unsigned(52, 10), 1473 => to_unsigned(590, 10), 1474 => to_unsigned(913, 10), 1475 => to_unsigned(918, 10), 1476 => to_unsigned(302, 10), 1477 => to_unsigned(543, 10), 1478 => to_unsigned(561, 10), 1479 => to_unsigned(797, 10), 1480 => to_unsigned(777, 10), 1481 => to_unsigned(92, 10), 1482 => to_unsigned(948, 10), 1483 => to_unsigned(1, 10), 1484 => to_unsigned(149, 10), 1485 => to_unsigned(227, 10), 1486 => to_unsigned(33, 10), 1487 => to_unsigned(354, 10), 1488 => to_unsigned(395, 10), 1489 => to_unsigned(632, 10), 1490 => to_unsigned(709, 10), 1491 => to_unsigned(170, 10), 1492 => to_unsigned(51, 10), 1493 => to_unsigned(141, 10), 1494 => to_unsigned(166, 10), 1495 => to_unsigned(303, 10), 1496 => to_unsigned(14, 10), 1497 => to_unsigned(159, 10), 1498 => to_unsigned(61, 10), 1499 => to_unsigned(988, 10), 1500 => to_unsigned(220, 10), 1501 => to_unsigned(729, 10), 1502 => to_unsigned(243, 10), 1503 => to_unsigned(501, 10), 1504 => to_unsigned(834, 10), 1505 => to_unsigned(253, 10), 1506 => to_unsigned(211, 10), 1507 => to_unsigned(45, 10), 1508 => to_unsigned(298, 10), 1509 => to_unsigned(150, 10), 1510 => to_unsigned(155, 10), 1511 => to_unsigned(907, 10), 1512 => to_unsigned(377, 10), 1513 => to_unsigned(566, 10), 1514 => to_unsigned(925, 10), 1515 => to_unsigned(624, 10), 1516 => to_unsigned(619, 10), 1517 => to_unsigned(333, 10), 1518 => to_unsigned(165, 10), 1519 => to_unsigned(180, 10), 1520 => to_unsigned(222, 10), 1521 => to_unsigned(611, 10), 1522 => to_unsigned(81, 10), 1523 => to_unsigned(544, 10), 1524 => to_unsigned(686, 10), 1525 => to_unsigned(571, 10), 1526 => to_unsigned(902, 10), 1527 => to_unsigned(921, 10), 1528 => to_unsigned(473, 10), 1529 => to_unsigned(199, 10), 1530 => to_unsigned(615, 10), 1531 => to_unsigned(415, 10), 1532 => to_unsigned(103, 10), 1533 => to_unsigned(653, 10), 1534 => to_unsigned(691, 10), 1535 => to_unsigned(24, 10), 1536 => to_unsigned(209, 10), 1537 => to_unsigned(503, 10), 1538 => to_unsigned(698, 10), 1539 => to_unsigned(861, 10), 1540 => to_unsigned(534, 10), 1541 => to_unsigned(412, 10), 1542 => to_unsigned(872, 10), 1543 => to_unsigned(820, 10), 1544 => to_unsigned(462, 10), 1545 => to_unsigned(360, 10), 1546 => to_unsigned(921, 10), 1547 => to_unsigned(239, 10), 1548 => to_unsigned(491, 10), 1549 => to_unsigned(276, 10), 1550 => to_unsigned(963, 10), 1551 => to_unsigned(203, 10), 1552 => to_unsigned(253, 10), 1553 => to_unsigned(397, 10), 1554 => to_unsigned(0, 10), 1555 => to_unsigned(485, 10), 1556 => to_unsigned(786, 10), 1557 => to_unsigned(297, 10), 1558 => to_unsigned(768, 10), 1559 => to_unsigned(76, 10), 1560 => to_unsigned(161, 10), 1561 => to_unsigned(798, 10), 1562 => to_unsigned(643, 10), 1563 => to_unsigned(419, 10), 1564 => to_unsigned(26, 10), 1565 => to_unsigned(382, 10), 1566 => to_unsigned(848, 10), 1567 => to_unsigned(556, 10), 1568 => to_unsigned(942, 10), 1569 => to_unsigned(643, 10), 1570 => to_unsigned(105, 10), 1571 => to_unsigned(955, 10), 1572 => to_unsigned(960, 10), 1573 => to_unsigned(641, 10), 1574 => to_unsigned(263, 10), 1575 => to_unsigned(606, 10), 1576 => to_unsigned(344, 10), 1577 => to_unsigned(415, 10), 1578 => to_unsigned(707, 10), 1579 => to_unsigned(112, 10), 1580 => to_unsigned(950, 10), 1581 => to_unsigned(763, 10), 1582 => to_unsigned(624, 10), 1583 => to_unsigned(610, 10), 1584 => to_unsigned(582, 10), 1585 => to_unsigned(776, 10), 1586 => to_unsigned(384, 10), 1587 => to_unsigned(919, 10), 1588 => to_unsigned(24, 10), 1589 => to_unsigned(990, 10), 1590 => to_unsigned(103, 10), 1591 => to_unsigned(730, 10), 1592 => to_unsigned(602, 10), 1593 => to_unsigned(37, 10), 1594 => to_unsigned(44, 10), 1595 => to_unsigned(843, 10), 1596 => to_unsigned(142, 10), 1597 => to_unsigned(701, 10), 1598 => to_unsigned(543, 10), 1599 => to_unsigned(109, 10), 1600 => to_unsigned(777, 10), 1601 => to_unsigned(1008, 10), 1602 => to_unsigned(142, 10), 1603 => to_unsigned(234, 10), 1604 => to_unsigned(202, 10), 1605 => to_unsigned(715, 10), 1606 => to_unsigned(927, 10), 1607 => to_unsigned(797, 10), 1608 => to_unsigned(434, 10), 1609 => to_unsigned(13, 10), 1610 => to_unsigned(787, 10), 1611 => to_unsigned(608, 10), 1612 => to_unsigned(627, 10), 1613 => to_unsigned(944, 10), 1614 => to_unsigned(414, 10), 1615 => to_unsigned(613, 10), 1616 => to_unsigned(216, 10), 1617 => to_unsigned(638, 10), 1618 => to_unsigned(399, 10), 1619 => to_unsigned(40, 10), 1620 => to_unsigned(267, 10), 1621 => to_unsigned(484, 10), 1622 => to_unsigned(639, 10), 1623 => to_unsigned(75, 10), 1624 => to_unsigned(73, 10), 1625 => to_unsigned(448, 10), 1626 => to_unsigned(857, 10), 1627 => to_unsigned(209, 10), 1628 => to_unsigned(576, 10), 1629 => to_unsigned(167, 10), 1630 => to_unsigned(886, 10), 1631 => to_unsigned(58, 10), 1632 => to_unsigned(623, 10), 1633 => to_unsigned(711, 10), 1634 => to_unsigned(47, 10), 1635 => to_unsigned(645, 10), 1636 => to_unsigned(964, 10), 1637 => to_unsigned(936, 10), 1638 => to_unsigned(472, 10), 1639 => to_unsigned(26, 10), 1640 => to_unsigned(1006, 10), 1641 => to_unsigned(210, 10), 1642 => to_unsigned(105, 10), 1643 => to_unsigned(588, 10), 1644 => to_unsigned(201, 10), 1645 => to_unsigned(914, 10), 1646 => to_unsigned(777, 10), 1647 => to_unsigned(996, 10), 1648 => to_unsigned(953, 10), 1649 => to_unsigned(1, 10), 1650 => to_unsigned(695, 10), 1651 => to_unsigned(558, 10), 1652 => to_unsigned(59, 10), 1653 => to_unsigned(683, 10), 1654 => to_unsigned(568, 10), 1655 => to_unsigned(308, 10), 1656 => to_unsigned(837, 10), 1657 => to_unsigned(155, 10), 1658 => to_unsigned(669, 10), 1659 => to_unsigned(298, 10), 1660 => to_unsigned(984, 10), 1661 => to_unsigned(636, 10), 1662 => to_unsigned(281, 10), 1663 => to_unsigned(365, 10), 1664 => to_unsigned(309, 10), 1665 => to_unsigned(754, 10), 1666 => to_unsigned(879, 10), 1667 => to_unsigned(594, 10), 1668 => to_unsigned(805, 10), 1669 => to_unsigned(788, 10), 1670 => to_unsigned(478, 10), 1671 => to_unsigned(439, 10), 1672 => to_unsigned(705, 10), 1673 => to_unsigned(270, 10), 1674 => to_unsigned(926, 10), 1675 => to_unsigned(346, 10), 1676 => to_unsigned(487, 10), 1677 => to_unsigned(104, 10), 1678 => to_unsigned(68, 10), 1679 => to_unsigned(696, 10), 1680 => to_unsigned(917, 10), 1681 => to_unsigned(96, 10), 1682 => to_unsigned(759, 10), 1683 => to_unsigned(453, 10), 1684 => to_unsigned(701, 10), 1685 => to_unsigned(946, 10), 1686 => to_unsigned(544, 10), 1687 => to_unsigned(946, 10), 1688 => to_unsigned(961, 10), 1689 => to_unsigned(417, 10), 1690 => to_unsigned(446, 10), 1691 => to_unsigned(281, 10), 1692 => to_unsigned(754, 10), 1693 => to_unsigned(701, 10), 1694 => to_unsigned(609, 10), 1695 => to_unsigned(405, 10), 1696 => to_unsigned(997, 10), 1697 => to_unsigned(950, 10), 1698 => to_unsigned(892, 10), 1699 => to_unsigned(553, 10), 1700 => to_unsigned(802, 10), 1701 => to_unsigned(403, 10), 1702 => to_unsigned(1000, 10), 1703 => to_unsigned(226, 10), 1704 => to_unsigned(942, 10), 1705 => to_unsigned(155, 10), 1706 => to_unsigned(908, 10), 1707 => to_unsigned(242, 10), 1708 => to_unsigned(36, 10), 1709 => to_unsigned(69, 10), 1710 => to_unsigned(163, 10), 1711 => to_unsigned(261, 10), 1712 => to_unsigned(994, 10), 1713 => to_unsigned(30, 10), 1714 => to_unsigned(321, 10), 1715 => to_unsigned(992, 10), 1716 => to_unsigned(131, 10), 1717 => to_unsigned(562, 10), 1718 => to_unsigned(950, 10), 1719 => to_unsigned(966, 10), 1720 => to_unsigned(983, 10), 1721 => to_unsigned(673, 10), 1722 => to_unsigned(683, 10), 1723 => to_unsigned(17, 10), 1724 => to_unsigned(820, 10), 1725 => to_unsigned(470, 10), 1726 => to_unsigned(157, 10), 1727 => to_unsigned(377, 10), 1728 => to_unsigned(346, 10), 1729 => to_unsigned(203, 10), 1730 => to_unsigned(751, 10), 1731 => to_unsigned(599, 10), 1732 => to_unsigned(444, 10), 1733 => to_unsigned(488, 10), 1734 => to_unsigned(426, 10), 1735 => to_unsigned(480, 10), 1736 => to_unsigned(500, 10), 1737 => to_unsigned(450, 10), 1738 => to_unsigned(377, 10), 1739 => to_unsigned(78, 10), 1740 => to_unsigned(269, 10), 1741 => to_unsigned(431, 10), 1742 => to_unsigned(398, 10), 1743 => to_unsigned(451, 10), 1744 => to_unsigned(878, 10), 1745 => to_unsigned(555, 10), 1746 => to_unsigned(635, 10), 1747 => to_unsigned(399, 10), 1748 => to_unsigned(340, 10), 1749 => to_unsigned(17, 10), 1750 => to_unsigned(645, 10), 1751 => to_unsigned(807, 10), 1752 => to_unsigned(944, 10), 1753 => to_unsigned(365, 10), 1754 => to_unsigned(961, 10), 1755 => to_unsigned(657, 10), 1756 => to_unsigned(464, 10), 1757 => to_unsigned(261, 10), 1758 => to_unsigned(170, 10), 1759 => to_unsigned(842, 10), 1760 => to_unsigned(91, 10), 1761 => to_unsigned(534, 10), 1762 => to_unsigned(362, 10), 1763 => to_unsigned(431, 10), 1764 => to_unsigned(847, 10), 1765 => to_unsigned(911, 10), 1766 => to_unsigned(653, 10), 1767 => to_unsigned(133, 10), 1768 => to_unsigned(793, 10), 1769 => to_unsigned(908, 10), 1770 => to_unsigned(660, 10), 1771 => to_unsigned(720, 10), 1772 => to_unsigned(283, 10), 1773 => to_unsigned(894, 10), 1774 => to_unsigned(28, 10), 1775 => to_unsigned(961, 10), 1776 => to_unsigned(859, 10), 1777 => to_unsigned(790, 10), 1778 => to_unsigned(624, 10), 1779 => to_unsigned(241, 10), 1780 => to_unsigned(154, 10), 1781 => to_unsigned(176, 10), 1782 => to_unsigned(938, 10), 1783 => to_unsigned(771, 10), 1784 => to_unsigned(661, 10), 1785 => to_unsigned(593, 10), 1786 => to_unsigned(371, 10), 1787 => to_unsigned(767, 10), 1788 => to_unsigned(221, 10), 1789 => to_unsigned(320, 10), 1790 => to_unsigned(516, 10), 1791 => to_unsigned(743, 10), 1792 => to_unsigned(600, 10), 1793 => to_unsigned(492, 10), 1794 => to_unsigned(479, 10), 1795 => to_unsigned(547, 10), 1796 => to_unsigned(573, 10), 1797 => to_unsigned(113, 10), 1798 => to_unsigned(694, 10), 1799 => to_unsigned(450, 10), 1800 => to_unsigned(89, 10), 1801 => to_unsigned(670, 10), 1802 => to_unsigned(977, 10), 1803 => to_unsigned(688, 10), 1804 => to_unsigned(264, 10), 1805 => to_unsigned(144, 10), 1806 => to_unsigned(120, 10), 1807 => to_unsigned(158, 10), 1808 => to_unsigned(195, 10), 1809 => to_unsigned(366, 10), 1810 => to_unsigned(791, 10), 1811 => to_unsigned(608, 10), 1812 => to_unsigned(47, 10), 1813 => to_unsigned(267, 10), 1814 => to_unsigned(301, 10), 1815 => to_unsigned(91, 10), 1816 => to_unsigned(164, 10), 1817 => to_unsigned(255, 10), 1818 => to_unsigned(284, 10), 1819 => to_unsigned(809, 10), 1820 => to_unsigned(731, 10), 1821 => to_unsigned(775, 10), 1822 => to_unsigned(956, 10), 1823 => to_unsigned(821, 10), 1824 => to_unsigned(376, 10), 1825 => to_unsigned(621, 10), 1826 => to_unsigned(120, 10), 1827 => to_unsigned(991, 10), 1828 => to_unsigned(82, 10), 1829 => to_unsigned(417, 10), 1830 => to_unsigned(942, 10), 1831 => to_unsigned(785, 10), 1832 => to_unsigned(1004, 10), 1833 => to_unsigned(901, 10), 1834 => to_unsigned(349, 10), 1835 => to_unsigned(358, 10), 1836 => to_unsigned(41, 10), 1837 => to_unsigned(442, 10), 1838 => to_unsigned(459, 10), 1839 => to_unsigned(613, 10), 1840 => to_unsigned(744, 10), 1841 => to_unsigned(904, 10), 1842 => to_unsigned(876, 10), 1843 => to_unsigned(484, 10), 1844 => to_unsigned(474, 10), 1845 => to_unsigned(985, 10), 1846 => to_unsigned(668, 10), 1847 => to_unsigned(858, 10), 1848 => to_unsigned(798, 10), 1849 => to_unsigned(730, 10), 1850 => to_unsigned(882, 10), 1851 => to_unsigned(384, 10), 1852 => to_unsigned(552, 10), 1853 => to_unsigned(121, 10), 1854 => to_unsigned(25, 10), 1855 => to_unsigned(679, 10), 1856 => to_unsigned(646, 10), 1857 => to_unsigned(643, 10), 1858 => to_unsigned(556, 10), 1859 => to_unsigned(587, 10), 1860 => to_unsigned(678, 10), 1861 => to_unsigned(170, 10), 1862 => to_unsigned(501, 10), 1863 => to_unsigned(582, 10), 1864 => to_unsigned(352, 10), 1865 => to_unsigned(62, 10), 1866 => to_unsigned(214, 10), 1867 => to_unsigned(407, 10), 1868 => to_unsigned(772, 10), 1869 => to_unsigned(66, 10), 1870 => to_unsigned(940, 10), 1871 => to_unsigned(871, 10), 1872 => to_unsigned(185, 10), 1873 => to_unsigned(319, 10), 1874 => to_unsigned(462, 10), 1875 => to_unsigned(795, 10), 1876 => to_unsigned(641, 10), 1877 => to_unsigned(109, 10), 1878 => to_unsigned(847, 10), 1879 => to_unsigned(302, 10), 1880 => to_unsigned(439, 10), 1881 => to_unsigned(1007, 10), 1882 => to_unsigned(788, 10), 1883 => to_unsigned(904, 10), 1884 => to_unsigned(104, 10), 1885 => to_unsigned(635, 10), 1886 => to_unsigned(272, 10), 1887 => to_unsigned(661, 10), 1888 => to_unsigned(374, 10), 1889 => to_unsigned(34, 10), 1890 => to_unsigned(805, 10), 1891 => to_unsigned(984, 10), 1892 => to_unsigned(899, 10), 1893 => to_unsigned(214, 10), 1894 => to_unsigned(895, 10), 1895 => to_unsigned(866, 10), 1896 => to_unsigned(334, 10), 1897 => to_unsigned(491, 10), 1898 => to_unsigned(267, 10), 1899 => to_unsigned(384, 10), 1900 => to_unsigned(925, 10), 1901 => to_unsigned(244, 10), 1902 => to_unsigned(205, 10), 1903 => to_unsigned(947, 10), 1904 => to_unsigned(278, 10), 1905 => to_unsigned(358, 10), 1906 => to_unsigned(666, 10), 1907 => to_unsigned(890, 10), 1908 => to_unsigned(821, 10), 1909 => to_unsigned(114, 10), 1910 => to_unsigned(413, 10), 1911 => to_unsigned(679, 10), 1912 => to_unsigned(183, 10), 1913 => to_unsigned(114, 10), 1914 => to_unsigned(519, 10), 1915 => to_unsigned(707, 10), 1916 => to_unsigned(940, 10), 1917 => to_unsigned(468, 10), 1918 => to_unsigned(351, 10), 1919 => to_unsigned(239, 10), 1920 => to_unsigned(7, 10), 1921 => to_unsigned(888, 10), 1922 => to_unsigned(206, 10), 1923 => to_unsigned(13, 10), 1924 => to_unsigned(617, 10), 1925 => to_unsigned(734, 10), 1926 => to_unsigned(497, 10), 1927 => to_unsigned(834, 10), 1928 => to_unsigned(889, 10), 1929 => to_unsigned(378, 10), 1930 => to_unsigned(262, 10), 1931 => to_unsigned(219, 10), 1932 => to_unsigned(519, 10), 1933 => to_unsigned(745, 10), 1934 => to_unsigned(133, 10), 1935 => to_unsigned(355, 10), 1936 => to_unsigned(44, 10), 1937 => to_unsigned(614, 10), 1938 => to_unsigned(971, 10), 1939 => to_unsigned(501, 10), 1940 => to_unsigned(932, 10), 1941 => to_unsigned(673, 10), 1942 => to_unsigned(875, 10), 1943 => to_unsigned(437, 10), 1944 => to_unsigned(858, 10), 1945 => to_unsigned(793, 10), 1946 => to_unsigned(908, 10), 1947 => to_unsigned(988, 10), 1948 => to_unsigned(951, 10), 1949 => to_unsigned(456, 10), 1950 => to_unsigned(556, 10), 1951 => to_unsigned(843, 10), 1952 => to_unsigned(1002, 10), 1953 => to_unsigned(513, 10), 1954 => to_unsigned(828, 10), 1955 => to_unsigned(682, 10), 1956 => to_unsigned(437, 10), 1957 => to_unsigned(530, 10), 1958 => to_unsigned(323, 10), 1959 => to_unsigned(130, 10), 1960 => to_unsigned(1017, 10), 1961 => to_unsigned(38, 10), 1962 => to_unsigned(904, 10), 1963 => to_unsigned(470, 10), 1964 => to_unsigned(611, 10), 1965 => to_unsigned(196, 10), 1966 => to_unsigned(682, 10), 1967 => to_unsigned(207, 10), 1968 => to_unsigned(926, 10), 1969 => to_unsigned(785, 10), 1970 => to_unsigned(702, 10), 1971 => to_unsigned(357, 10), 1972 => to_unsigned(196, 10), 1973 => to_unsigned(790, 10), 1974 => to_unsigned(627, 10), 1975 => to_unsigned(430, 10), 1976 => to_unsigned(754, 10), 1977 => to_unsigned(134, 10), 1978 => to_unsigned(665, 10), 1979 => to_unsigned(982, 10), 1980 => to_unsigned(627, 10), 1981 => to_unsigned(184, 10), 1982 => to_unsigned(611, 10), 1983 => to_unsigned(828, 10), 1984 => to_unsigned(965, 10), 1985 => to_unsigned(188, 10), 1986 => to_unsigned(298, 10), 1987 => to_unsigned(986, 10), 1988 => to_unsigned(262, 10), 1989 => to_unsigned(484, 10), 1990 => to_unsigned(42, 10), 1991 => to_unsigned(291, 10), 1992 => to_unsigned(692, 10), 1993 => to_unsigned(536, 10), 1994 => to_unsigned(528, 10), 1995 => to_unsigned(847, 10), 1996 => to_unsigned(851, 10), 1997 => to_unsigned(669, 10), 1998 => to_unsigned(193, 10), 1999 => to_unsigned(414, 10), 2000 => to_unsigned(324, 10), 2001 => to_unsigned(1002, 10), 2002 => to_unsigned(633, 10), 2003 => to_unsigned(312, 10), 2004 => to_unsigned(96, 10), 2005 => to_unsigned(696, 10), 2006 => to_unsigned(531, 10), 2007 => to_unsigned(88, 10), 2008 => to_unsigned(1008, 10), 2009 => to_unsigned(441, 10), 2010 => to_unsigned(690, 10), 2011 => to_unsigned(755, 10), 2012 => to_unsigned(370, 10), 2013 => to_unsigned(435, 10), 2014 => to_unsigned(747, 10), 2015 => to_unsigned(2, 10), 2016 => to_unsigned(173, 10), 2017 => to_unsigned(285, 10), 2018 => to_unsigned(781, 10), 2019 => to_unsigned(770, 10), 2020 => to_unsigned(300, 10), 2021 => to_unsigned(112, 10), 2022 => to_unsigned(385, 10), 2023 => to_unsigned(688, 10), 2024 => to_unsigned(655, 10), 2025 => to_unsigned(68, 10), 2026 => to_unsigned(227, 10), 2027 => to_unsigned(50, 10), 2028 => to_unsigned(591, 10), 2029 => to_unsigned(702, 10), 2030 => to_unsigned(918, 10), 2031 => to_unsigned(148, 10), 2032 => to_unsigned(481, 10), 2033 => to_unsigned(546, 10), 2034 => to_unsigned(194, 10), 2035 => to_unsigned(799, 10), 2036 => to_unsigned(638, 10), 2037 => to_unsigned(387, 10), 2038 => to_unsigned(261, 10), 2039 => to_unsigned(213, 10), 2040 => to_unsigned(621, 10), 2041 => to_unsigned(575, 10), 2042 => to_unsigned(895, 10), 2043 => to_unsigned(684, 10), 2044 => to_unsigned(810, 10), 2045 => to_unsigned(651, 10), 2046 => to_unsigned(257, 10), 2047 => to_unsigned(595, 10)),
            9 => (0 => to_unsigned(597, 10), 1 => to_unsigned(874, 10), 2 => to_unsigned(536, 10), 3 => to_unsigned(785, 10), 4 => to_unsigned(743, 10), 5 => to_unsigned(483, 10), 6 => to_unsigned(1010, 10), 7 => to_unsigned(43, 10), 8 => to_unsigned(248, 10), 9 => to_unsigned(524, 10), 10 => to_unsigned(251, 10), 11 => to_unsigned(429, 10), 12 => to_unsigned(429, 10), 13 => to_unsigned(191, 10), 14 => to_unsigned(897, 10), 15 => to_unsigned(601, 10), 16 => to_unsigned(508, 10), 17 => to_unsigned(90, 10), 18 => to_unsigned(991, 10), 19 => to_unsigned(616, 10), 20 => to_unsigned(831, 10), 21 => to_unsigned(896, 10), 22 => to_unsigned(138, 10), 23 => to_unsigned(689, 10), 24 => to_unsigned(679, 10), 25 => to_unsigned(149, 10), 26 => to_unsigned(972, 10), 27 => to_unsigned(559, 10), 28 => to_unsigned(98, 10), 29 => to_unsigned(396, 10), 30 => to_unsigned(247, 10), 31 => to_unsigned(683, 10), 32 => to_unsigned(423, 10), 33 => to_unsigned(339, 10), 34 => to_unsigned(46, 10), 35 => to_unsigned(558, 10), 36 => to_unsigned(998, 10), 37 => to_unsigned(312, 10), 38 => to_unsigned(833, 10), 39 => to_unsigned(580, 10), 40 => to_unsigned(432, 10), 41 => to_unsigned(98, 10), 42 => to_unsigned(610, 10), 43 => to_unsigned(856, 10), 44 => to_unsigned(680, 10), 45 => to_unsigned(340, 10), 46 => to_unsigned(648, 10), 47 => to_unsigned(30, 10), 48 => to_unsigned(915, 10), 49 => to_unsigned(28, 10), 50 => to_unsigned(359, 10), 51 => to_unsigned(301, 10), 52 => to_unsigned(598, 10), 53 => to_unsigned(392, 10), 54 => to_unsigned(910, 10), 55 => to_unsigned(777, 10), 56 => to_unsigned(767, 10), 57 => to_unsigned(237, 10), 58 => to_unsigned(278, 10), 59 => to_unsigned(309, 10), 60 => to_unsigned(949, 10), 61 => to_unsigned(398, 10), 62 => to_unsigned(911, 10), 63 => to_unsigned(818, 10), 64 => to_unsigned(1019, 10), 65 => to_unsigned(816, 10), 66 => to_unsigned(579, 10), 67 => to_unsigned(66, 10), 68 => to_unsigned(646, 10), 69 => to_unsigned(158, 10), 70 => to_unsigned(289, 10), 71 => to_unsigned(886, 10), 72 => to_unsigned(797, 10), 73 => to_unsigned(880, 10), 74 => to_unsigned(243, 10), 75 => to_unsigned(596, 10), 76 => to_unsigned(331, 10), 77 => to_unsigned(91, 10), 78 => to_unsigned(372, 10), 79 => to_unsigned(616, 10), 80 => to_unsigned(576, 10), 81 => to_unsigned(552, 10), 82 => to_unsigned(858, 10), 83 => to_unsigned(471, 10), 84 => to_unsigned(932, 10), 85 => to_unsigned(857, 10), 86 => to_unsigned(93, 10), 87 => to_unsigned(87, 10), 88 => to_unsigned(700, 10), 89 => to_unsigned(966, 10), 90 => to_unsigned(540, 10), 91 => to_unsigned(228, 10), 92 => to_unsigned(635, 10), 93 => to_unsigned(138, 10), 94 => to_unsigned(796, 10), 95 => to_unsigned(643, 10), 96 => to_unsigned(180, 10), 97 => to_unsigned(602, 10), 98 => to_unsigned(767, 10), 99 => to_unsigned(795, 10), 100 => to_unsigned(631, 10), 101 => to_unsigned(726, 10), 102 => to_unsigned(725, 10), 103 => to_unsigned(409, 10), 104 => to_unsigned(129, 10), 105 => to_unsigned(766, 10), 106 => to_unsigned(879, 10), 107 => to_unsigned(58, 10), 108 => to_unsigned(548, 10), 109 => to_unsigned(960, 10), 110 => to_unsigned(221, 10), 111 => to_unsigned(1021, 10), 112 => to_unsigned(223, 10), 113 => to_unsigned(620, 10), 114 => to_unsigned(278, 10), 115 => to_unsigned(237, 10), 116 => to_unsigned(715, 10), 117 => to_unsigned(641, 10), 118 => to_unsigned(309, 10), 119 => to_unsigned(256, 10), 120 => to_unsigned(527, 10), 121 => to_unsigned(69, 10), 122 => to_unsigned(811, 10), 123 => to_unsigned(160, 10), 124 => to_unsigned(119, 10), 125 => to_unsigned(484, 10), 126 => to_unsigned(1021, 10), 127 => to_unsigned(730, 10), 128 => to_unsigned(528, 10), 129 => to_unsigned(792, 10), 130 => to_unsigned(546, 10), 131 => to_unsigned(893, 10), 132 => to_unsigned(1000, 10), 133 => to_unsigned(580, 10), 134 => to_unsigned(829, 10), 135 => to_unsigned(600, 10), 136 => to_unsigned(881, 10), 137 => to_unsigned(436, 10), 138 => to_unsigned(451, 10), 139 => to_unsigned(519, 10), 140 => to_unsigned(247, 10), 141 => to_unsigned(729, 10), 142 => to_unsigned(672, 10), 143 => to_unsigned(180, 10), 144 => to_unsigned(34, 10), 145 => to_unsigned(473, 10), 146 => to_unsigned(78, 10), 147 => to_unsigned(268, 10), 148 => to_unsigned(643, 10), 149 => to_unsigned(718, 10), 150 => to_unsigned(703, 10), 151 => to_unsigned(45, 10), 152 => to_unsigned(753, 10), 153 => to_unsigned(253, 10), 154 => to_unsigned(329, 10), 155 => to_unsigned(502, 10), 156 => to_unsigned(779, 10), 157 => to_unsigned(569, 10), 158 => to_unsigned(671, 10), 159 => to_unsigned(770, 10), 160 => to_unsigned(855, 10), 161 => to_unsigned(842, 10), 162 => to_unsigned(599, 10), 163 => to_unsigned(655, 10), 164 => to_unsigned(660, 10), 165 => to_unsigned(200, 10), 166 => to_unsigned(823, 10), 167 => to_unsigned(7, 10), 168 => to_unsigned(642, 10), 169 => to_unsigned(486, 10), 170 => to_unsigned(749, 10), 171 => to_unsigned(926, 10), 172 => to_unsigned(563, 10), 173 => to_unsigned(241, 10), 174 => to_unsigned(628, 10), 175 => to_unsigned(846, 10), 176 => to_unsigned(764, 10), 177 => to_unsigned(289, 10), 178 => to_unsigned(112, 10), 179 => to_unsigned(778, 10), 180 => to_unsigned(283, 10), 181 => to_unsigned(224, 10), 182 => to_unsigned(921, 10), 183 => to_unsigned(868, 10), 184 => to_unsigned(287, 10), 185 => to_unsigned(739, 10), 186 => to_unsigned(115, 10), 187 => to_unsigned(654, 10), 188 => to_unsigned(244, 10), 189 => to_unsigned(522, 10), 190 => to_unsigned(856, 10), 191 => to_unsigned(612, 10), 192 => to_unsigned(477, 10), 193 => to_unsigned(7, 10), 194 => to_unsigned(433, 10), 195 => to_unsigned(95, 10), 196 => to_unsigned(371, 10), 197 => to_unsigned(336, 10), 198 => to_unsigned(637, 10), 199 => to_unsigned(339, 10), 200 => to_unsigned(264, 10), 201 => to_unsigned(614, 10), 202 => to_unsigned(371, 10), 203 => to_unsigned(295, 10), 204 => to_unsigned(998, 10), 205 => to_unsigned(172, 10), 206 => to_unsigned(230, 10), 207 => to_unsigned(112, 10), 208 => to_unsigned(378, 10), 209 => to_unsigned(623, 10), 210 => to_unsigned(1, 10), 211 => to_unsigned(409, 10), 212 => to_unsigned(64, 10), 213 => to_unsigned(85, 10), 214 => to_unsigned(172, 10), 215 => to_unsigned(777, 10), 216 => to_unsigned(114, 10), 217 => to_unsigned(96, 10), 218 => to_unsigned(750, 10), 219 => to_unsigned(985, 10), 220 => to_unsigned(643, 10), 221 => to_unsigned(881, 10), 222 => to_unsigned(522, 10), 223 => to_unsigned(332, 10), 224 => to_unsigned(74, 10), 225 => to_unsigned(613, 10), 226 => to_unsigned(430, 10), 227 => to_unsigned(300, 10), 228 => to_unsigned(560, 10), 229 => to_unsigned(635, 10), 230 => to_unsigned(79, 10), 231 => to_unsigned(150, 10), 232 => to_unsigned(489, 10), 233 => to_unsigned(136, 10), 234 => to_unsigned(996, 10), 235 => to_unsigned(1000, 10), 236 => to_unsigned(56, 10), 237 => to_unsigned(362, 10), 238 => to_unsigned(705, 10), 239 => to_unsigned(485, 10), 240 => to_unsigned(178, 10), 241 => to_unsigned(660, 10), 242 => to_unsigned(24, 10), 243 => to_unsigned(628, 10), 244 => to_unsigned(985, 10), 245 => to_unsigned(961, 10), 246 => to_unsigned(71, 10), 247 => to_unsigned(80, 10), 248 => to_unsigned(192, 10), 249 => to_unsigned(756, 10), 250 => to_unsigned(136, 10), 251 => to_unsigned(850, 10), 252 => to_unsigned(548, 10), 253 => to_unsigned(534, 10), 254 => to_unsigned(230, 10), 255 => to_unsigned(502, 10), 256 => to_unsigned(82, 10), 257 => to_unsigned(317, 10), 258 => to_unsigned(564, 10), 259 => to_unsigned(630, 10), 260 => to_unsigned(346, 10), 261 => to_unsigned(565, 10), 262 => to_unsigned(906, 10), 263 => to_unsigned(522, 10), 264 => to_unsigned(948, 10), 265 => to_unsigned(315, 10), 266 => to_unsigned(111, 10), 267 => to_unsigned(812, 10), 268 => to_unsigned(816, 10), 269 => to_unsigned(339, 10), 270 => to_unsigned(762, 10), 271 => to_unsigned(426, 10), 272 => to_unsigned(528, 10), 273 => to_unsigned(231, 10), 274 => to_unsigned(381, 10), 275 => to_unsigned(558, 10), 276 => to_unsigned(548, 10), 277 => to_unsigned(494, 10), 278 => to_unsigned(460, 10), 279 => to_unsigned(219, 10), 280 => to_unsigned(867, 10), 281 => to_unsigned(16, 10), 282 => to_unsigned(391, 10), 283 => to_unsigned(137, 10), 284 => to_unsigned(746, 10), 285 => to_unsigned(825, 10), 286 => to_unsigned(709, 10), 287 => to_unsigned(262, 10), 288 => to_unsigned(547, 10), 289 => to_unsigned(624, 10), 290 => to_unsigned(656, 10), 291 => to_unsigned(583, 10), 292 => to_unsigned(862, 10), 293 => to_unsigned(621, 10), 294 => to_unsigned(320, 10), 295 => to_unsigned(567, 10), 296 => to_unsigned(455, 10), 297 => to_unsigned(771, 10), 298 => to_unsigned(47, 10), 299 => to_unsigned(899, 10), 300 => to_unsigned(152, 10), 301 => to_unsigned(513, 10), 302 => to_unsigned(133, 10), 303 => to_unsigned(676, 10), 304 => to_unsigned(662, 10), 305 => to_unsigned(217, 10), 306 => to_unsigned(645, 10), 307 => to_unsigned(821, 10), 308 => to_unsigned(910, 10), 309 => to_unsigned(127, 10), 310 => to_unsigned(207, 10), 311 => to_unsigned(165, 10), 312 => to_unsigned(562, 10), 313 => to_unsigned(322, 10), 314 => to_unsigned(989, 10), 315 => to_unsigned(819, 10), 316 => to_unsigned(186, 10), 317 => to_unsigned(322, 10), 318 => to_unsigned(71, 10), 319 => to_unsigned(895, 10), 320 => to_unsigned(583, 10), 321 => to_unsigned(912, 10), 322 => to_unsigned(20, 10), 323 => to_unsigned(999, 10), 324 => to_unsigned(594, 10), 325 => to_unsigned(685, 10), 326 => to_unsigned(361, 10), 327 => to_unsigned(1014, 10), 328 => to_unsigned(602, 10), 329 => to_unsigned(358, 10), 330 => to_unsigned(282, 10), 331 => to_unsigned(206, 10), 332 => to_unsigned(346, 10), 333 => to_unsigned(252, 10), 334 => to_unsigned(484, 10), 335 => to_unsigned(769, 10), 336 => to_unsigned(588, 10), 337 => to_unsigned(266, 10), 338 => to_unsigned(657, 10), 339 => to_unsigned(13, 10), 340 => to_unsigned(911, 10), 341 => to_unsigned(177, 10), 342 => to_unsigned(718, 10), 343 => to_unsigned(803, 10), 344 => to_unsigned(130, 10), 345 => to_unsigned(468, 10), 346 => to_unsigned(781, 10), 347 => to_unsigned(743, 10), 348 => to_unsigned(648, 10), 349 => to_unsigned(15, 10), 350 => to_unsigned(532, 10), 351 => to_unsigned(1023, 10), 352 => to_unsigned(148, 10), 353 => to_unsigned(914, 10), 354 => to_unsigned(519, 10), 355 => to_unsigned(990, 10), 356 => to_unsigned(603, 10), 357 => to_unsigned(248, 10), 358 => to_unsigned(203, 10), 359 => to_unsigned(514, 10), 360 => to_unsigned(640, 10), 361 => to_unsigned(303, 10), 362 => to_unsigned(960, 10), 363 => to_unsigned(861, 10), 364 => to_unsigned(298, 10), 365 => to_unsigned(1014, 10), 366 => to_unsigned(1010, 10), 367 => to_unsigned(483, 10), 368 => to_unsigned(682, 10), 369 => to_unsigned(540, 10), 370 => to_unsigned(1018, 10), 371 => to_unsigned(82, 10), 372 => to_unsigned(677, 10), 373 => to_unsigned(9, 10), 374 => to_unsigned(393, 10), 375 => to_unsigned(672, 10), 376 => to_unsigned(237, 10), 377 => to_unsigned(927, 10), 378 => to_unsigned(55, 10), 379 => to_unsigned(248, 10), 380 => to_unsigned(966, 10), 381 => to_unsigned(79, 10), 382 => to_unsigned(981, 10), 383 => to_unsigned(229, 10), 384 => to_unsigned(348, 10), 385 => to_unsigned(555, 10), 386 => to_unsigned(954, 10), 387 => to_unsigned(708, 10), 388 => to_unsigned(838, 10), 389 => to_unsigned(958, 10), 390 => to_unsigned(246, 10), 391 => to_unsigned(351, 10), 392 => to_unsigned(966, 10), 393 => to_unsigned(575, 10), 394 => to_unsigned(618, 10), 395 => to_unsigned(100, 10), 396 => to_unsigned(111, 10), 397 => to_unsigned(1000, 10), 398 => to_unsigned(112, 10), 399 => to_unsigned(242, 10), 400 => to_unsigned(923, 10), 401 => to_unsigned(360, 10), 402 => to_unsigned(315, 10), 403 => to_unsigned(943, 10), 404 => to_unsigned(855, 10), 405 => to_unsigned(603, 10), 406 => to_unsigned(410, 10), 407 => to_unsigned(413, 10), 408 => to_unsigned(257, 10), 409 => to_unsigned(717, 10), 410 => to_unsigned(678, 10), 411 => to_unsigned(719, 10), 412 => to_unsigned(250, 10), 413 => to_unsigned(860, 10), 414 => to_unsigned(487, 10), 415 => to_unsigned(221, 10), 416 => to_unsigned(419, 10), 417 => to_unsigned(460, 10), 418 => to_unsigned(664, 10), 419 => to_unsigned(289, 10), 420 => to_unsigned(879, 10), 421 => to_unsigned(234, 10), 422 => to_unsigned(898, 10), 423 => to_unsigned(616, 10), 424 => to_unsigned(318, 10), 425 => to_unsigned(877, 10), 426 => to_unsigned(63, 10), 427 => to_unsigned(693, 10), 428 => to_unsigned(432, 10), 429 => to_unsigned(940, 10), 430 => to_unsigned(165, 10), 431 => to_unsigned(16, 10), 432 => to_unsigned(295, 10), 433 => to_unsigned(336, 10), 434 => to_unsigned(686, 10), 435 => to_unsigned(826, 10), 436 => to_unsigned(292, 10), 437 => to_unsigned(769, 10), 438 => to_unsigned(93, 10), 439 => to_unsigned(85, 10), 440 => to_unsigned(461, 10), 441 => to_unsigned(321, 10), 442 => to_unsigned(160, 10), 443 => to_unsigned(800, 10), 444 => to_unsigned(266, 10), 445 => to_unsigned(158, 10), 446 => to_unsigned(447, 10), 447 => to_unsigned(547, 10), 448 => to_unsigned(334, 10), 449 => to_unsigned(211, 10), 450 => to_unsigned(386, 10), 451 => to_unsigned(547, 10), 452 => to_unsigned(822, 10), 453 => to_unsigned(560, 10), 454 => to_unsigned(703, 10), 455 => to_unsigned(937, 10), 456 => to_unsigned(293, 10), 457 => to_unsigned(414, 10), 458 => to_unsigned(161, 10), 459 => to_unsigned(525, 10), 460 => to_unsigned(533, 10), 461 => to_unsigned(629, 10), 462 => to_unsigned(414, 10), 463 => to_unsigned(524, 10), 464 => to_unsigned(435, 10), 465 => to_unsigned(218, 10), 466 => to_unsigned(79, 10), 467 => to_unsigned(29, 10), 468 => to_unsigned(71, 10), 469 => to_unsigned(557, 10), 470 => to_unsigned(239, 10), 471 => to_unsigned(719, 10), 472 => to_unsigned(394, 10), 473 => to_unsigned(872, 10), 474 => to_unsigned(247, 10), 475 => to_unsigned(639, 10), 476 => to_unsigned(152, 10), 477 => to_unsigned(81, 10), 478 => to_unsigned(987, 10), 479 => to_unsigned(171, 10), 480 => to_unsigned(323, 10), 481 => to_unsigned(268, 10), 482 => to_unsigned(436, 10), 483 => to_unsigned(170, 10), 484 => to_unsigned(889, 10), 485 => to_unsigned(977, 10), 486 => to_unsigned(803, 10), 487 => to_unsigned(931, 10), 488 => to_unsigned(407, 10), 489 => to_unsigned(114, 10), 490 => to_unsigned(1020, 10), 491 => to_unsigned(51, 10), 492 => to_unsigned(888, 10), 493 => to_unsigned(829, 10), 494 => to_unsigned(92, 10), 495 => to_unsigned(836, 10), 496 => to_unsigned(946, 10), 497 => to_unsigned(879, 10), 498 => to_unsigned(422, 10), 499 => to_unsigned(197, 10), 500 => to_unsigned(463, 10), 501 => to_unsigned(398, 10), 502 => to_unsigned(870, 10), 503 => to_unsigned(55, 10), 504 => to_unsigned(85, 10), 505 => to_unsigned(460, 10), 506 => to_unsigned(573, 10), 507 => to_unsigned(683, 10), 508 => to_unsigned(976, 10), 509 => to_unsigned(360, 10), 510 => to_unsigned(83, 10), 511 => to_unsigned(890, 10), 512 => to_unsigned(435, 10), 513 => to_unsigned(792, 10), 514 => to_unsigned(977, 10), 515 => to_unsigned(819, 10), 516 => to_unsigned(699, 10), 517 => to_unsigned(683, 10), 518 => to_unsigned(201, 10), 519 => to_unsigned(645, 10), 520 => to_unsigned(1010, 10), 521 => to_unsigned(483, 10), 522 => to_unsigned(793, 10), 523 => to_unsigned(457, 10), 524 => to_unsigned(708, 10), 525 => to_unsigned(593, 10), 526 => to_unsigned(93, 10), 527 => to_unsigned(202, 10), 528 => to_unsigned(981, 10), 529 => to_unsigned(497, 10), 530 => to_unsigned(29, 10), 531 => to_unsigned(296, 10), 532 => to_unsigned(185, 10), 533 => to_unsigned(665, 10), 534 => to_unsigned(297, 10), 535 => to_unsigned(580, 10), 536 => to_unsigned(65, 10), 537 => to_unsigned(698, 10), 538 => to_unsigned(678, 10), 539 => to_unsigned(492, 10), 540 => to_unsigned(130, 10), 541 => to_unsigned(480, 10), 542 => to_unsigned(434, 10), 543 => to_unsigned(641, 10), 544 => to_unsigned(886, 10), 545 => to_unsigned(430, 10), 546 => to_unsigned(1014, 10), 547 => to_unsigned(881, 10), 548 => to_unsigned(625, 10), 549 => to_unsigned(398, 10), 550 => to_unsigned(401, 10), 551 => to_unsigned(834, 10), 552 => to_unsigned(131, 10), 553 => to_unsigned(655, 10), 554 => to_unsigned(967, 10), 555 => to_unsigned(469, 10), 556 => to_unsigned(683, 10), 557 => to_unsigned(71, 10), 558 => to_unsigned(52, 10), 559 => to_unsigned(401, 10), 560 => to_unsigned(539, 10), 561 => to_unsigned(680, 10), 562 => to_unsigned(788, 10), 563 => to_unsigned(191, 10), 564 => to_unsigned(245, 10), 565 => to_unsigned(400, 10), 566 => to_unsigned(625, 10), 567 => to_unsigned(491, 10), 568 => to_unsigned(285, 10), 569 => to_unsigned(617, 10), 570 => to_unsigned(476, 10), 571 => to_unsigned(711, 10), 572 => to_unsigned(69, 10), 573 => to_unsigned(519, 10), 574 => to_unsigned(634, 10), 575 => to_unsigned(946, 10), 576 => to_unsigned(872, 10), 577 => to_unsigned(165, 10), 578 => to_unsigned(985, 10), 579 => to_unsigned(704, 10), 580 => to_unsigned(218, 10), 581 => to_unsigned(112, 10), 582 => to_unsigned(685, 10), 583 => to_unsigned(523, 10), 584 => to_unsigned(592, 10), 585 => to_unsigned(532, 10), 586 => to_unsigned(660, 10), 587 => to_unsigned(284, 10), 588 => to_unsigned(439, 10), 589 => to_unsigned(1009, 10), 590 => to_unsigned(402, 10), 591 => to_unsigned(329, 10), 592 => to_unsigned(482, 10), 593 => to_unsigned(323, 10), 594 => to_unsigned(641, 10), 595 => to_unsigned(581, 10), 596 => to_unsigned(355, 10), 597 => to_unsigned(403, 10), 598 => to_unsigned(860, 10), 599 => to_unsigned(531, 10), 600 => to_unsigned(556, 10), 601 => to_unsigned(50, 10), 602 => to_unsigned(259, 10), 603 => to_unsigned(275, 10), 604 => to_unsigned(437, 10), 605 => to_unsigned(501, 10), 606 => to_unsigned(522, 10), 607 => to_unsigned(881, 10), 608 => to_unsigned(612, 10), 609 => to_unsigned(483, 10), 610 => to_unsigned(829, 10), 611 => to_unsigned(594, 10), 612 => to_unsigned(273, 10), 613 => to_unsigned(874, 10), 614 => to_unsigned(445, 10), 615 => to_unsigned(950, 10), 616 => to_unsigned(693, 10), 617 => to_unsigned(860, 10), 618 => to_unsigned(612, 10), 619 => to_unsigned(655, 10), 620 => to_unsigned(933, 10), 621 => to_unsigned(818, 10), 622 => to_unsigned(758, 10), 623 => to_unsigned(934, 10), 624 => to_unsigned(395, 10), 625 => to_unsigned(719, 10), 626 => to_unsigned(234, 10), 627 => to_unsigned(822, 10), 628 => to_unsigned(821, 10), 629 => to_unsigned(712, 10), 630 => to_unsigned(957, 10), 631 => to_unsigned(875, 10), 632 => to_unsigned(601, 10), 633 => to_unsigned(463, 10), 634 => to_unsigned(591, 10), 635 => to_unsigned(320, 10), 636 => to_unsigned(175, 10), 637 => to_unsigned(949, 10), 638 => to_unsigned(890, 10), 639 => to_unsigned(744, 10), 640 => to_unsigned(212, 10), 641 => to_unsigned(493, 10), 642 => to_unsigned(463, 10), 643 => to_unsigned(937, 10), 644 => to_unsigned(809, 10), 645 => to_unsigned(537, 10), 646 => to_unsigned(460, 10), 647 => to_unsigned(464, 10), 648 => to_unsigned(466, 10), 649 => to_unsigned(301, 10), 650 => to_unsigned(91, 10), 651 => to_unsigned(25, 10), 652 => to_unsigned(110, 10), 653 => to_unsigned(655, 10), 654 => to_unsigned(564, 10), 655 => to_unsigned(292, 10), 656 => to_unsigned(844, 10), 657 => to_unsigned(334, 10), 658 => to_unsigned(503, 10), 659 => to_unsigned(841, 10), 660 => to_unsigned(924, 10), 661 => to_unsigned(808, 10), 662 => to_unsigned(297, 10), 663 => to_unsigned(989, 10), 664 => to_unsigned(557, 10), 665 => to_unsigned(522, 10), 666 => to_unsigned(798, 10), 667 => to_unsigned(520, 10), 668 => to_unsigned(742, 10), 669 => to_unsigned(132, 10), 670 => to_unsigned(1011, 10), 671 => to_unsigned(462, 10), 672 => to_unsigned(104, 10), 673 => to_unsigned(408, 10), 674 => to_unsigned(871, 10), 675 => to_unsigned(712, 10), 676 => to_unsigned(341, 10), 677 => to_unsigned(145, 10), 678 => to_unsigned(106, 10), 679 => to_unsigned(135, 10), 680 => to_unsigned(905, 10), 681 => to_unsigned(872, 10), 682 => to_unsigned(981, 10), 683 => to_unsigned(897, 10), 684 => to_unsigned(415, 10), 685 => to_unsigned(409, 10), 686 => to_unsigned(824, 10), 687 => to_unsigned(681, 10), 688 => to_unsigned(694, 10), 689 => to_unsigned(220, 10), 690 => to_unsigned(645, 10), 691 => to_unsigned(225, 10), 692 => to_unsigned(647, 10), 693 => to_unsigned(624, 10), 694 => to_unsigned(939, 10), 695 => to_unsigned(1004, 10), 696 => to_unsigned(553, 10), 697 => to_unsigned(204, 10), 698 => to_unsigned(770, 10), 699 => to_unsigned(918, 10), 700 => to_unsigned(98, 10), 701 => to_unsigned(882, 10), 702 => to_unsigned(646, 10), 703 => to_unsigned(1018, 10), 704 => to_unsigned(600, 10), 705 => to_unsigned(812, 10), 706 => to_unsigned(532, 10), 707 => to_unsigned(602, 10), 708 => to_unsigned(51, 10), 709 => to_unsigned(891, 10), 710 => to_unsigned(753, 10), 711 => to_unsigned(630, 10), 712 => to_unsigned(171, 10), 713 => to_unsigned(451, 10), 714 => to_unsigned(783, 10), 715 => to_unsigned(301, 10), 716 => to_unsigned(738, 10), 717 => to_unsigned(732, 10), 718 => to_unsigned(692, 10), 719 => to_unsigned(610, 10), 720 => to_unsigned(857, 10), 721 => to_unsigned(384, 10), 722 => to_unsigned(563, 10), 723 => to_unsigned(507, 10), 724 => to_unsigned(890, 10), 725 => to_unsigned(646, 10), 726 => to_unsigned(430, 10), 727 => to_unsigned(946, 10), 728 => to_unsigned(370, 10), 729 => to_unsigned(664, 10), 730 => to_unsigned(386, 10), 731 => to_unsigned(169, 10), 732 => to_unsigned(326, 10), 733 => to_unsigned(310, 10), 734 => to_unsigned(607, 10), 735 => to_unsigned(669, 10), 736 => to_unsigned(415, 10), 737 => to_unsigned(488, 10), 738 => to_unsigned(590, 10), 739 => to_unsigned(684, 10), 740 => to_unsigned(695, 10), 741 => to_unsigned(454, 10), 742 => to_unsigned(119, 10), 743 => to_unsigned(394, 10), 744 => to_unsigned(644, 10), 745 => to_unsigned(445, 10), 746 => to_unsigned(431, 10), 747 => to_unsigned(577, 10), 748 => to_unsigned(807, 10), 749 => to_unsigned(26, 10), 750 => to_unsigned(643, 10), 751 => to_unsigned(229, 10), 752 => to_unsigned(186, 10), 753 => to_unsigned(608, 10), 754 => to_unsigned(913, 10), 755 => to_unsigned(887, 10), 756 => to_unsigned(90, 10), 757 => to_unsigned(778, 10), 758 => to_unsigned(409, 10), 759 => to_unsigned(543, 10), 760 => to_unsigned(169, 10), 761 => to_unsigned(960, 10), 762 => to_unsigned(805, 10), 763 => to_unsigned(758, 10), 764 => to_unsigned(741, 10), 765 => to_unsigned(288, 10), 766 => to_unsigned(396, 10), 767 => to_unsigned(108, 10), 768 => to_unsigned(364, 10), 769 => to_unsigned(552, 10), 770 => to_unsigned(32, 10), 771 => to_unsigned(567, 10), 772 => to_unsigned(685, 10), 773 => to_unsigned(245, 10), 774 => to_unsigned(792, 10), 775 => to_unsigned(489, 10), 776 => to_unsigned(418, 10), 777 => to_unsigned(807, 10), 778 => to_unsigned(926, 10), 779 => to_unsigned(822, 10), 780 => to_unsigned(307, 10), 781 => to_unsigned(687, 10), 782 => to_unsigned(749, 10), 783 => to_unsigned(35, 10), 784 => to_unsigned(577, 10), 785 => to_unsigned(108, 10), 786 => to_unsigned(379, 10), 787 => to_unsigned(642, 10), 788 => to_unsigned(506, 10), 789 => to_unsigned(979, 10), 790 => to_unsigned(729, 10), 791 => to_unsigned(761, 10), 792 => to_unsigned(9, 10), 793 => to_unsigned(904, 10), 794 => to_unsigned(956, 10), 795 => to_unsigned(482, 10), 796 => to_unsigned(637, 10), 797 => to_unsigned(815, 10), 798 => to_unsigned(630, 10), 799 => to_unsigned(513, 10), 800 => to_unsigned(132, 10), 801 => to_unsigned(325, 10), 802 => to_unsigned(152, 10), 803 => to_unsigned(933, 10), 804 => to_unsigned(901, 10), 805 => to_unsigned(51, 10), 806 => to_unsigned(839, 10), 807 => to_unsigned(490, 10), 808 => to_unsigned(760, 10), 809 => to_unsigned(540, 10), 810 => to_unsigned(629, 10), 811 => to_unsigned(579, 10), 812 => to_unsigned(766, 10), 813 => to_unsigned(397, 10), 814 => to_unsigned(677, 10), 815 => to_unsigned(192, 10), 816 => to_unsigned(139, 10), 817 => to_unsigned(629, 10), 818 => to_unsigned(340, 10), 819 => to_unsigned(316, 10), 820 => to_unsigned(571, 10), 821 => to_unsigned(353, 10), 822 => to_unsigned(157, 10), 823 => to_unsigned(854, 10), 824 => to_unsigned(474, 10), 825 => to_unsigned(327, 10), 826 => to_unsigned(481, 10), 827 => to_unsigned(166, 10), 828 => to_unsigned(612, 10), 829 => to_unsigned(17, 10), 830 => to_unsigned(777, 10), 831 => to_unsigned(621, 10), 832 => to_unsigned(793, 10), 833 => to_unsigned(677, 10), 834 => to_unsigned(892, 10), 835 => to_unsigned(81, 10), 836 => to_unsigned(539, 10), 837 => to_unsigned(474, 10), 838 => to_unsigned(90, 10), 839 => to_unsigned(462, 10), 840 => to_unsigned(182, 10), 841 => to_unsigned(990, 10), 842 => to_unsigned(551, 10), 843 => to_unsigned(691, 10), 844 => to_unsigned(241, 10), 845 => to_unsigned(870, 10), 846 => to_unsigned(999, 10), 847 => to_unsigned(252, 10), 848 => to_unsigned(709, 10), 849 => to_unsigned(888, 10), 850 => to_unsigned(681, 10), 851 => to_unsigned(893, 10), 852 => to_unsigned(259, 10), 853 => to_unsigned(572, 10), 854 => to_unsigned(78, 10), 855 => to_unsigned(794, 10), 856 => to_unsigned(342, 10), 857 => to_unsigned(120, 10), 858 => to_unsigned(1013, 10), 859 => to_unsigned(690, 10), 860 => to_unsigned(339, 10), 861 => to_unsigned(46, 10), 862 => to_unsigned(970, 10), 863 => to_unsigned(749, 10), 864 => to_unsigned(854, 10), 865 => to_unsigned(626, 10), 866 => to_unsigned(332, 10), 867 => to_unsigned(339, 10), 868 => to_unsigned(797, 10), 869 => to_unsigned(353, 10), 870 => to_unsigned(504, 10), 871 => to_unsigned(752, 10), 872 => to_unsigned(323, 10), 873 => to_unsigned(218, 10), 874 => to_unsigned(988, 10), 875 => to_unsigned(559, 10), 876 => to_unsigned(739, 10), 877 => to_unsigned(931, 10), 878 => to_unsigned(179, 10), 879 => to_unsigned(201, 10), 880 => to_unsigned(604, 10), 881 => to_unsigned(85, 10), 882 => to_unsigned(440, 10), 883 => to_unsigned(14, 10), 884 => to_unsigned(335, 10), 885 => to_unsigned(248, 10), 886 => to_unsigned(158, 10), 887 => to_unsigned(499, 10), 888 => to_unsigned(765, 10), 889 => to_unsigned(177, 10), 890 => to_unsigned(136, 10), 891 => to_unsigned(496, 10), 892 => to_unsigned(827, 10), 893 => to_unsigned(148, 10), 894 => to_unsigned(730, 10), 895 => to_unsigned(565, 10), 896 => to_unsigned(123, 10), 897 => to_unsigned(14, 10), 898 => to_unsigned(156, 10), 899 => to_unsigned(936, 10), 900 => to_unsigned(988, 10), 901 => to_unsigned(211, 10), 902 => to_unsigned(244, 10), 903 => to_unsigned(931, 10), 904 => to_unsigned(515, 10), 905 => to_unsigned(627, 10), 906 => to_unsigned(333, 10), 907 => to_unsigned(336, 10), 908 => to_unsigned(549, 10), 909 => to_unsigned(75, 10), 910 => to_unsigned(974, 10), 911 => to_unsigned(74, 10), 912 => to_unsigned(182, 10), 913 => to_unsigned(89, 10), 914 => to_unsigned(163, 10), 915 => to_unsigned(473, 10), 916 => to_unsigned(174, 10), 917 => to_unsigned(161, 10), 918 => to_unsigned(201, 10), 919 => to_unsigned(858, 10), 920 => to_unsigned(586, 10), 921 => to_unsigned(346, 10), 922 => to_unsigned(262, 10), 923 => to_unsigned(361, 10), 924 => to_unsigned(639, 10), 925 => to_unsigned(804, 10), 926 => to_unsigned(797, 10), 927 => to_unsigned(403, 10), 928 => to_unsigned(579, 10), 929 => to_unsigned(820, 10), 930 => to_unsigned(674, 10), 931 => to_unsigned(104, 10), 932 => to_unsigned(370, 10), 933 => to_unsigned(232, 10), 934 => to_unsigned(1023, 10), 935 => to_unsigned(706, 10), 936 => to_unsigned(1011, 10), 937 => to_unsigned(455, 10), 938 => to_unsigned(733, 10), 939 => to_unsigned(242, 10), 940 => to_unsigned(913, 10), 941 => to_unsigned(944, 10), 942 => to_unsigned(183, 10), 943 => to_unsigned(169, 10), 944 => to_unsigned(54, 10), 945 => to_unsigned(861, 10), 946 => to_unsigned(790, 10), 947 => to_unsigned(417, 10), 948 => to_unsigned(461, 10), 949 => to_unsigned(401, 10), 950 => to_unsigned(263, 10), 951 => to_unsigned(814, 10), 952 => to_unsigned(676, 10), 953 => to_unsigned(708, 10), 954 => to_unsigned(539, 10), 955 => to_unsigned(788, 10), 956 => to_unsigned(490, 10), 957 => to_unsigned(646, 10), 958 => to_unsigned(113, 10), 959 => to_unsigned(75, 10), 960 => to_unsigned(942, 10), 961 => to_unsigned(407, 10), 962 => to_unsigned(457, 10), 963 => to_unsigned(760, 10), 964 => to_unsigned(117, 10), 965 => to_unsigned(478, 10), 966 => to_unsigned(825, 10), 967 => to_unsigned(551, 10), 968 => to_unsigned(15, 10), 969 => to_unsigned(268, 10), 970 => to_unsigned(538, 10), 971 => to_unsigned(760, 10), 972 => to_unsigned(133, 10), 973 => to_unsigned(894, 10), 974 => to_unsigned(357, 10), 975 => to_unsigned(581, 10), 976 => to_unsigned(568, 10), 977 => to_unsigned(338, 10), 978 => to_unsigned(397, 10), 979 => to_unsigned(309, 10), 980 => to_unsigned(126, 10), 981 => to_unsigned(192, 10), 982 => to_unsigned(1013, 10), 983 => to_unsigned(786, 10), 984 => to_unsigned(315, 10), 985 => to_unsigned(894, 10), 986 => to_unsigned(540, 10), 987 => to_unsigned(102, 10), 988 => to_unsigned(133, 10), 989 => to_unsigned(979, 10), 990 => to_unsigned(81, 10), 991 => to_unsigned(685, 10), 992 => to_unsigned(430, 10), 993 => to_unsigned(60, 10), 994 => to_unsigned(998, 10), 995 => to_unsigned(921, 10), 996 => to_unsigned(797, 10), 997 => to_unsigned(654, 10), 998 => to_unsigned(762, 10), 999 => to_unsigned(707, 10), 1000 => to_unsigned(482, 10), 1001 => to_unsigned(305, 10), 1002 => to_unsigned(963, 10), 1003 => to_unsigned(423, 10), 1004 => to_unsigned(971, 10), 1005 => to_unsigned(40, 10), 1006 => to_unsigned(681, 10), 1007 => to_unsigned(725, 10), 1008 => to_unsigned(28, 10), 1009 => to_unsigned(344, 10), 1010 => to_unsigned(582, 10), 1011 => to_unsigned(522, 10), 1012 => to_unsigned(849, 10), 1013 => to_unsigned(65, 10), 1014 => to_unsigned(274, 10), 1015 => to_unsigned(335, 10), 1016 => to_unsigned(867, 10), 1017 => to_unsigned(508, 10), 1018 => to_unsigned(460, 10), 1019 => to_unsigned(741, 10), 1020 => to_unsigned(444, 10), 1021 => to_unsigned(643, 10), 1022 => to_unsigned(437, 10), 1023 => to_unsigned(261, 10), 1024 => to_unsigned(958, 10), 1025 => to_unsigned(186, 10), 1026 => to_unsigned(977, 10), 1027 => to_unsigned(75, 10), 1028 => to_unsigned(62, 10), 1029 => to_unsigned(636, 10), 1030 => to_unsigned(179, 10), 1031 => to_unsigned(941, 10), 1032 => to_unsigned(916, 10), 1033 => to_unsigned(199, 10), 1034 => to_unsigned(510, 10), 1035 => to_unsigned(571, 10), 1036 => to_unsigned(90, 10), 1037 => to_unsigned(545, 10), 1038 => to_unsigned(355, 10), 1039 => to_unsigned(731, 10), 1040 => to_unsigned(858, 10), 1041 => to_unsigned(38, 10), 1042 => to_unsigned(357, 10), 1043 => to_unsigned(538, 10), 1044 => to_unsigned(474, 10), 1045 => to_unsigned(558, 10), 1046 => to_unsigned(982, 10), 1047 => to_unsigned(0, 10), 1048 => to_unsigned(852, 10), 1049 => to_unsigned(757, 10), 1050 => to_unsigned(68, 10), 1051 => to_unsigned(591, 10), 1052 => to_unsigned(764, 10), 1053 => to_unsigned(838, 10), 1054 => to_unsigned(859, 10), 1055 => to_unsigned(639, 10), 1056 => to_unsigned(917, 10), 1057 => to_unsigned(347, 10), 1058 => to_unsigned(174, 10), 1059 => to_unsigned(910, 10), 1060 => to_unsigned(599, 10), 1061 => to_unsigned(397, 10), 1062 => to_unsigned(380, 10), 1063 => to_unsigned(895, 10), 1064 => to_unsigned(929, 10), 1065 => to_unsigned(638, 10), 1066 => to_unsigned(650, 10), 1067 => to_unsigned(948, 10), 1068 => to_unsigned(92, 10), 1069 => to_unsigned(51, 10), 1070 => to_unsigned(1007, 10), 1071 => to_unsigned(376, 10), 1072 => to_unsigned(45, 10), 1073 => to_unsigned(346, 10), 1074 => to_unsigned(800, 10), 1075 => to_unsigned(1021, 10), 1076 => to_unsigned(661, 10), 1077 => to_unsigned(651, 10), 1078 => to_unsigned(339, 10), 1079 => to_unsigned(107, 10), 1080 => to_unsigned(889, 10), 1081 => to_unsigned(20, 10), 1082 => to_unsigned(167, 10), 1083 => to_unsigned(201, 10), 1084 => to_unsigned(490, 10), 1085 => to_unsigned(406, 10), 1086 => to_unsigned(868, 10), 1087 => to_unsigned(220, 10), 1088 => to_unsigned(629, 10), 1089 => to_unsigned(656, 10), 1090 => to_unsigned(227, 10), 1091 => to_unsigned(240, 10), 1092 => to_unsigned(256, 10), 1093 => to_unsigned(217, 10), 1094 => to_unsigned(996, 10), 1095 => to_unsigned(175, 10), 1096 => to_unsigned(568, 10), 1097 => to_unsigned(334, 10), 1098 => to_unsigned(213, 10), 1099 => to_unsigned(636, 10), 1100 => to_unsigned(57, 10), 1101 => to_unsigned(735, 10), 1102 => to_unsigned(330, 10), 1103 => to_unsigned(737, 10), 1104 => to_unsigned(441, 10), 1105 => to_unsigned(36, 10), 1106 => to_unsigned(927, 10), 1107 => to_unsigned(40, 10), 1108 => to_unsigned(375, 10), 1109 => to_unsigned(134, 10), 1110 => to_unsigned(790, 10), 1111 => to_unsigned(803, 10), 1112 => to_unsigned(657, 10), 1113 => to_unsigned(710, 10), 1114 => to_unsigned(259, 10), 1115 => to_unsigned(169, 10), 1116 => to_unsigned(907, 10), 1117 => to_unsigned(523, 10), 1118 => to_unsigned(401, 10), 1119 => to_unsigned(250, 10), 1120 => to_unsigned(823, 10), 1121 => to_unsigned(249, 10), 1122 => to_unsigned(744, 10), 1123 => to_unsigned(834, 10), 1124 => to_unsigned(666, 10), 1125 => to_unsigned(391, 10), 1126 => to_unsigned(722, 10), 1127 => to_unsigned(1009, 10), 1128 => to_unsigned(945, 10), 1129 => to_unsigned(67, 10), 1130 => to_unsigned(263, 10), 1131 => to_unsigned(764, 10), 1132 => to_unsigned(1007, 10), 1133 => to_unsigned(567, 10), 1134 => to_unsigned(683, 10), 1135 => to_unsigned(958, 10), 1136 => to_unsigned(654, 10), 1137 => to_unsigned(585, 10), 1138 => to_unsigned(493, 10), 1139 => to_unsigned(531, 10), 1140 => to_unsigned(753, 10), 1141 => to_unsigned(219, 10), 1142 => to_unsigned(648, 10), 1143 => to_unsigned(460, 10), 1144 => to_unsigned(498, 10), 1145 => to_unsigned(661, 10), 1146 => to_unsigned(638, 10), 1147 => to_unsigned(465, 10), 1148 => to_unsigned(315, 10), 1149 => to_unsigned(769, 10), 1150 => to_unsigned(89, 10), 1151 => to_unsigned(763, 10), 1152 => to_unsigned(100, 10), 1153 => to_unsigned(855, 10), 1154 => to_unsigned(59, 10), 1155 => to_unsigned(836, 10), 1156 => to_unsigned(570, 10), 1157 => to_unsigned(31, 10), 1158 => to_unsigned(484, 10), 1159 => to_unsigned(664, 10), 1160 => to_unsigned(424, 10), 1161 => to_unsigned(658, 10), 1162 => to_unsigned(343, 10), 1163 => to_unsigned(32, 10), 1164 => to_unsigned(504, 10), 1165 => to_unsigned(257, 10), 1166 => to_unsigned(231, 10), 1167 => to_unsigned(477, 10), 1168 => to_unsigned(433, 10), 1169 => to_unsigned(539, 10), 1170 => to_unsigned(975, 10), 1171 => to_unsigned(573, 10), 1172 => to_unsigned(580, 10), 1173 => to_unsigned(162, 10), 1174 => to_unsigned(708, 10), 1175 => to_unsigned(708, 10), 1176 => to_unsigned(960, 10), 1177 => to_unsigned(749, 10), 1178 => to_unsigned(508, 10), 1179 => to_unsigned(413, 10), 1180 => to_unsigned(790, 10), 1181 => to_unsigned(694, 10), 1182 => to_unsigned(31, 10), 1183 => to_unsigned(16, 10), 1184 => to_unsigned(772, 10), 1185 => to_unsigned(644, 10), 1186 => to_unsigned(439, 10), 1187 => to_unsigned(607, 10), 1188 => to_unsigned(350, 10), 1189 => to_unsigned(109, 10), 1190 => to_unsigned(823, 10), 1191 => to_unsigned(455, 10), 1192 => to_unsigned(962, 10), 1193 => to_unsigned(395, 10), 1194 => to_unsigned(866, 10), 1195 => to_unsigned(990, 10), 1196 => to_unsigned(758, 10), 1197 => to_unsigned(167, 10), 1198 => to_unsigned(177, 10), 1199 => to_unsigned(638, 10), 1200 => to_unsigned(354, 10), 1201 => to_unsigned(933, 10), 1202 => to_unsigned(14, 10), 1203 => to_unsigned(317, 10), 1204 => to_unsigned(765, 10), 1205 => to_unsigned(902, 10), 1206 => to_unsigned(248, 10), 1207 => to_unsigned(321, 10), 1208 => to_unsigned(1008, 10), 1209 => to_unsigned(355, 10), 1210 => to_unsigned(717, 10), 1211 => to_unsigned(771, 10), 1212 => to_unsigned(35, 10), 1213 => to_unsigned(474, 10), 1214 => to_unsigned(1006, 10), 1215 => to_unsigned(150, 10), 1216 => to_unsigned(319, 10), 1217 => to_unsigned(651, 10), 1218 => to_unsigned(798, 10), 1219 => to_unsigned(615, 10), 1220 => to_unsigned(706, 10), 1221 => to_unsigned(893, 10), 1222 => to_unsigned(282, 10), 1223 => to_unsigned(320, 10), 1224 => to_unsigned(460, 10), 1225 => to_unsigned(264, 10), 1226 => to_unsigned(119, 10), 1227 => to_unsigned(193, 10), 1228 => to_unsigned(379, 10), 1229 => to_unsigned(639, 10), 1230 => to_unsigned(431, 10), 1231 => to_unsigned(284, 10), 1232 => to_unsigned(181, 10), 1233 => to_unsigned(949, 10), 1234 => to_unsigned(631, 10), 1235 => to_unsigned(383, 10), 1236 => to_unsigned(664, 10), 1237 => to_unsigned(643, 10), 1238 => to_unsigned(799, 10), 1239 => to_unsigned(665, 10), 1240 => to_unsigned(562, 10), 1241 => to_unsigned(213, 10), 1242 => to_unsigned(441, 10), 1243 => to_unsigned(738, 10), 1244 => to_unsigned(590, 10), 1245 => to_unsigned(215, 10), 1246 => to_unsigned(693, 10), 1247 => to_unsigned(309, 10), 1248 => to_unsigned(45, 10), 1249 => to_unsigned(116, 10), 1250 => to_unsigned(704, 10), 1251 => to_unsigned(433, 10), 1252 => to_unsigned(388, 10), 1253 => to_unsigned(623, 10), 1254 => to_unsigned(678, 10), 1255 => to_unsigned(496, 10), 1256 => to_unsigned(639, 10), 1257 => to_unsigned(855, 10), 1258 => to_unsigned(748, 10), 1259 => to_unsigned(116, 10), 1260 => to_unsigned(731, 10), 1261 => to_unsigned(238, 10), 1262 => to_unsigned(848, 10), 1263 => to_unsigned(1, 10), 1264 => to_unsigned(355, 10), 1265 => to_unsigned(451, 10), 1266 => to_unsigned(852, 10), 1267 => to_unsigned(354, 10), 1268 => to_unsigned(7, 10), 1269 => to_unsigned(487, 10), 1270 => to_unsigned(620, 10), 1271 => to_unsigned(246, 10), 1272 => to_unsigned(208, 10), 1273 => to_unsigned(994, 10), 1274 => to_unsigned(526, 10), 1275 => to_unsigned(194, 10), 1276 => to_unsigned(532, 10), 1277 => to_unsigned(917, 10), 1278 => to_unsigned(37, 10), 1279 => to_unsigned(839, 10), 1280 => to_unsigned(153, 10), 1281 => to_unsigned(320, 10), 1282 => to_unsigned(450, 10), 1283 => to_unsigned(435, 10), 1284 => to_unsigned(84, 10), 1285 => to_unsigned(984, 10), 1286 => to_unsigned(294, 10), 1287 => to_unsigned(848, 10), 1288 => to_unsigned(850, 10), 1289 => to_unsigned(281, 10), 1290 => to_unsigned(880, 10), 1291 => to_unsigned(124, 10), 1292 => to_unsigned(107, 10), 1293 => to_unsigned(635, 10), 1294 => to_unsigned(549, 10), 1295 => to_unsigned(926, 10), 1296 => to_unsigned(36, 10), 1297 => to_unsigned(711, 10), 1298 => to_unsigned(69, 10), 1299 => to_unsigned(3, 10), 1300 => to_unsigned(972, 10), 1301 => to_unsigned(25, 10), 1302 => to_unsigned(597, 10), 1303 => to_unsigned(305, 10), 1304 => to_unsigned(185, 10), 1305 => to_unsigned(386, 10), 1306 => to_unsigned(75, 10), 1307 => to_unsigned(93, 10), 1308 => to_unsigned(567, 10), 1309 => to_unsigned(193, 10), 1310 => to_unsigned(820, 10), 1311 => to_unsigned(91, 10), 1312 => to_unsigned(694, 10), 1313 => to_unsigned(460, 10), 1314 => to_unsigned(95, 10), 1315 => to_unsigned(847, 10), 1316 => to_unsigned(926, 10), 1317 => to_unsigned(535, 10), 1318 => to_unsigned(188, 10), 1319 => to_unsigned(508, 10), 1320 => to_unsigned(867, 10), 1321 => to_unsigned(261, 10), 1322 => to_unsigned(856, 10), 1323 => to_unsigned(553, 10), 1324 => to_unsigned(336, 10), 1325 => to_unsigned(718, 10), 1326 => to_unsigned(3, 10), 1327 => to_unsigned(763, 10), 1328 => to_unsigned(487, 10), 1329 => to_unsigned(38, 10), 1330 => to_unsigned(493, 10), 1331 => to_unsigned(837, 10), 1332 => to_unsigned(221, 10), 1333 => to_unsigned(722, 10), 1334 => to_unsigned(219, 10), 1335 => to_unsigned(636, 10), 1336 => to_unsigned(868, 10), 1337 => to_unsigned(318, 10), 1338 => to_unsigned(131, 10), 1339 => to_unsigned(732, 10), 1340 => to_unsigned(271, 10), 1341 => to_unsigned(127, 10), 1342 => to_unsigned(124, 10), 1343 => to_unsigned(3, 10), 1344 => to_unsigned(461, 10), 1345 => to_unsigned(919, 10), 1346 => to_unsigned(630, 10), 1347 => to_unsigned(679, 10), 1348 => to_unsigned(421, 10), 1349 => to_unsigned(896, 10), 1350 => to_unsigned(609, 10), 1351 => to_unsigned(490, 10), 1352 => to_unsigned(35, 10), 1353 => to_unsigned(832, 10), 1354 => to_unsigned(558, 10), 1355 => to_unsigned(882, 10), 1356 => to_unsigned(385, 10), 1357 => to_unsigned(381, 10), 1358 => to_unsigned(174, 10), 1359 => to_unsigned(1000, 10), 1360 => to_unsigned(564, 10), 1361 => to_unsigned(572, 10), 1362 => to_unsigned(416, 10), 1363 => to_unsigned(551, 10), 1364 => to_unsigned(894, 10), 1365 => to_unsigned(717, 10), 1366 => to_unsigned(257, 10), 1367 => to_unsigned(131, 10), 1368 => to_unsigned(272, 10), 1369 => to_unsigned(181, 10), 1370 => to_unsigned(91, 10), 1371 => to_unsigned(942, 10), 1372 => to_unsigned(515, 10), 1373 => to_unsigned(788, 10), 1374 => to_unsigned(984, 10), 1375 => to_unsigned(30, 10), 1376 => to_unsigned(737, 10), 1377 => to_unsigned(111, 10), 1378 => to_unsigned(177, 10), 1379 => to_unsigned(787, 10), 1380 => to_unsigned(749, 10), 1381 => to_unsigned(902, 10), 1382 => to_unsigned(483, 10), 1383 => to_unsigned(45, 10), 1384 => to_unsigned(998, 10), 1385 => to_unsigned(578, 10), 1386 => to_unsigned(701, 10), 1387 => to_unsigned(126, 10), 1388 => to_unsigned(126, 10), 1389 => to_unsigned(711, 10), 1390 => to_unsigned(498, 10), 1391 => to_unsigned(33, 10), 1392 => to_unsigned(784, 10), 1393 => to_unsigned(108, 10), 1394 => to_unsigned(808, 10), 1395 => to_unsigned(156, 10), 1396 => to_unsigned(576, 10), 1397 => to_unsigned(220, 10), 1398 => to_unsigned(717, 10), 1399 => to_unsigned(998, 10), 1400 => to_unsigned(933, 10), 1401 => to_unsigned(1012, 10), 1402 => to_unsigned(280, 10), 1403 => to_unsigned(379, 10), 1404 => to_unsigned(556, 10), 1405 => to_unsigned(14, 10), 1406 => to_unsigned(413, 10), 1407 => to_unsigned(329, 10), 1408 => to_unsigned(531, 10), 1409 => to_unsigned(605, 10), 1410 => to_unsigned(32, 10), 1411 => to_unsigned(74, 10), 1412 => to_unsigned(884, 10), 1413 => to_unsigned(965, 10), 1414 => to_unsigned(58, 10), 1415 => to_unsigned(207, 10), 1416 => to_unsigned(626, 10), 1417 => to_unsigned(826, 10), 1418 => to_unsigned(182, 10), 1419 => to_unsigned(843, 10), 1420 => to_unsigned(961, 10), 1421 => to_unsigned(779, 10), 1422 => to_unsigned(57, 10), 1423 => to_unsigned(7, 10), 1424 => to_unsigned(522, 10), 1425 => to_unsigned(973, 10), 1426 => to_unsigned(52, 10), 1427 => to_unsigned(793, 10), 1428 => to_unsigned(399, 10), 1429 => to_unsigned(527, 10), 1430 => to_unsigned(893, 10), 1431 => to_unsigned(825, 10), 1432 => to_unsigned(846, 10), 1433 => to_unsigned(61, 10), 1434 => to_unsigned(443, 10), 1435 => to_unsigned(686, 10), 1436 => to_unsigned(918, 10), 1437 => to_unsigned(390, 10), 1438 => to_unsigned(209, 10), 1439 => to_unsigned(155, 10), 1440 => to_unsigned(570, 10), 1441 => to_unsigned(831, 10), 1442 => to_unsigned(167, 10), 1443 => to_unsigned(155, 10), 1444 => to_unsigned(365, 10), 1445 => to_unsigned(49, 10), 1446 => to_unsigned(16, 10), 1447 => to_unsigned(398, 10), 1448 => to_unsigned(339, 10), 1449 => to_unsigned(614, 10), 1450 => to_unsigned(919, 10), 1451 => to_unsigned(163, 10), 1452 => to_unsigned(925, 10), 1453 => to_unsigned(557, 10), 1454 => to_unsigned(25, 10), 1455 => to_unsigned(433, 10), 1456 => to_unsigned(557, 10), 1457 => to_unsigned(244, 10), 1458 => to_unsigned(414, 10), 1459 => to_unsigned(764, 10), 1460 => to_unsigned(392, 10), 1461 => to_unsigned(260, 10), 1462 => to_unsigned(199, 10), 1463 => to_unsigned(139, 10), 1464 => to_unsigned(479, 10), 1465 => to_unsigned(430, 10), 1466 => to_unsigned(816, 10), 1467 => to_unsigned(1003, 10), 1468 => to_unsigned(958, 10), 1469 => to_unsigned(38, 10), 1470 => to_unsigned(156, 10), 1471 => to_unsigned(251, 10), 1472 => to_unsigned(623, 10), 1473 => to_unsigned(1018, 10), 1474 => to_unsigned(369, 10), 1475 => to_unsigned(408, 10), 1476 => to_unsigned(185, 10), 1477 => to_unsigned(1008, 10), 1478 => to_unsigned(604, 10), 1479 => to_unsigned(62, 10), 1480 => to_unsigned(758, 10), 1481 => to_unsigned(129, 10), 1482 => to_unsigned(545, 10), 1483 => to_unsigned(208, 10), 1484 => to_unsigned(25, 10), 1485 => to_unsigned(332, 10), 1486 => to_unsigned(249, 10), 1487 => to_unsigned(510, 10), 1488 => to_unsigned(955, 10), 1489 => to_unsigned(460, 10), 1490 => to_unsigned(356, 10), 1491 => to_unsigned(21, 10), 1492 => to_unsigned(651, 10), 1493 => to_unsigned(644, 10), 1494 => to_unsigned(932, 10), 1495 => to_unsigned(995, 10), 1496 => to_unsigned(967, 10), 1497 => to_unsigned(433, 10), 1498 => to_unsigned(518, 10), 1499 => to_unsigned(405, 10), 1500 => to_unsigned(148, 10), 1501 => to_unsigned(833, 10), 1502 => to_unsigned(562, 10), 1503 => to_unsigned(1002, 10), 1504 => to_unsigned(873, 10), 1505 => to_unsigned(799, 10), 1506 => to_unsigned(932, 10), 1507 => to_unsigned(298, 10), 1508 => to_unsigned(813, 10), 1509 => to_unsigned(372, 10), 1510 => to_unsigned(10, 10), 1511 => to_unsigned(95, 10), 1512 => to_unsigned(342, 10), 1513 => to_unsigned(38, 10), 1514 => to_unsigned(864, 10), 1515 => to_unsigned(177, 10), 1516 => to_unsigned(196, 10), 1517 => to_unsigned(997, 10), 1518 => to_unsigned(936, 10), 1519 => to_unsigned(47, 10), 1520 => to_unsigned(477, 10), 1521 => to_unsigned(54, 10), 1522 => to_unsigned(753, 10), 1523 => to_unsigned(178, 10), 1524 => to_unsigned(368, 10), 1525 => to_unsigned(973, 10), 1526 => to_unsigned(728, 10), 1527 => to_unsigned(705, 10), 1528 => to_unsigned(304, 10), 1529 => to_unsigned(393, 10), 1530 => to_unsigned(943, 10), 1531 => to_unsigned(904, 10), 1532 => to_unsigned(149, 10), 1533 => to_unsigned(891, 10), 1534 => to_unsigned(286, 10), 1535 => to_unsigned(28, 10), 1536 => to_unsigned(893, 10), 1537 => to_unsigned(328, 10), 1538 => to_unsigned(636, 10), 1539 => to_unsigned(637, 10), 1540 => to_unsigned(103, 10), 1541 => to_unsigned(549, 10), 1542 => to_unsigned(250, 10), 1543 => to_unsigned(190, 10), 1544 => to_unsigned(149, 10), 1545 => to_unsigned(964, 10), 1546 => to_unsigned(453, 10), 1547 => to_unsigned(212, 10), 1548 => to_unsigned(483, 10), 1549 => to_unsigned(262, 10), 1550 => to_unsigned(248, 10), 1551 => to_unsigned(982, 10), 1552 => to_unsigned(652, 10), 1553 => to_unsigned(863, 10), 1554 => to_unsigned(989, 10), 1555 => to_unsigned(974, 10), 1556 => to_unsigned(730, 10), 1557 => to_unsigned(51, 10), 1558 => to_unsigned(88, 10), 1559 => to_unsigned(349, 10), 1560 => to_unsigned(188, 10), 1561 => to_unsigned(473, 10), 1562 => to_unsigned(252, 10), 1563 => to_unsigned(589, 10), 1564 => to_unsigned(899, 10), 1565 => to_unsigned(64, 10), 1566 => to_unsigned(887, 10), 1567 => to_unsigned(642, 10), 1568 => to_unsigned(823, 10), 1569 => to_unsigned(680, 10), 1570 => to_unsigned(469, 10), 1571 => to_unsigned(135, 10), 1572 => to_unsigned(678, 10), 1573 => to_unsigned(25, 10), 1574 => to_unsigned(198, 10), 1575 => to_unsigned(351, 10), 1576 => to_unsigned(928, 10), 1577 => to_unsigned(685, 10), 1578 => to_unsigned(13, 10), 1579 => to_unsigned(490, 10), 1580 => to_unsigned(853, 10), 1581 => to_unsigned(223, 10), 1582 => to_unsigned(247, 10), 1583 => to_unsigned(701, 10), 1584 => to_unsigned(921, 10), 1585 => to_unsigned(236, 10), 1586 => to_unsigned(77, 10), 1587 => to_unsigned(437, 10), 1588 => to_unsigned(813, 10), 1589 => to_unsigned(835, 10), 1590 => to_unsigned(813, 10), 1591 => to_unsigned(753, 10), 1592 => to_unsigned(229, 10), 1593 => to_unsigned(497, 10), 1594 => to_unsigned(620, 10), 1595 => to_unsigned(333, 10), 1596 => to_unsigned(807, 10), 1597 => to_unsigned(90, 10), 1598 => to_unsigned(420, 10), 1599 => to_unsigned(333, 10), 1600 => to_unsigned(145, 10), 1601 => to_unsigned(30, 10), 1602 => to_unsigned(499, 10), 1603 => to_unsigned(484, 10), 1604 => to_unsigned(999, 10), 1605 => to_unsigned(371, 10), 1606 => to_unsigned(802, 10), 1607 => to_unsigned(716, 10), 1608 => to_unsigned(132, 10), 1609 => to_unsigned(214, 10), 1610 => to_unsigned(81, 10), 1611 => to_unsigned(439, 10), 1612 => to_unsigned(360, 10), 1613 => to_unsigned(186, 10), 1614 => to_unsigned(99, 10), 1615 => to_unsigned(200, 10), 1616 => to_unsigned(345, 10), 1617 => to_unsigned(716, 10), 1618 => to_unsigned(283, 10), 1619 => to_unsigned(923, 10), 1620 => to_unsigned(365, 10), 1621 => to_unsigned(22, 10), 1622 => to_unsigned(394, 10), 1623 => to_unsigned(855, 10), 1624 => to_unsigned(495, 10), 1625 => to_unsigned(411, 10), 1626 => to_unsigned(729, 10), 1627 => to_unsigned(931, 10), 1628 => to_unsigned(82, 10), 1629 => to_unsigned(640, 10), 1630 => to_unsigned(220, 10), 1631 => to_unsigned(323, 10), 1632 => to_unsigned(437, 10), 1633 => to_unsigned(297, 10), 1634 => to_unsigned(251, 10), 1635 => to_unsigned(126, 10), 1636 => to_unsigned(155, 10), 1637 => to_unsigned(815, 10), 1638 => to_unsigned(260, 10), 1639 => to_unsigned(146, 10), 1640 => to_unsigned(134, 10), 1641 => to_unsigned(717, 10), 1642 => to_unsigned(466, 10), 1643 => to_unsigned(683, 10), 1644 => to_unsigned(264, 10), 1645 => to_unsigned(345, 10), 1646 => to_unsigned(17, 10), 1647 => to_unsigned(51, 10), 1648 => to_unsigned(720, 10), 1649 => to_unsigned(852, 10), 1650 => to_unsigned(337, 10), 1651 => to_unsigned(973, 10), 1652 => to_unsigned(256, 10), 1653 => to_unsigned(466, 10), 1654 => to_unsigned(421, 10), 1655 => to_unsigned(414, 10), 1656 => to_unsigned(852, 10), 1657 => to_unsigned(105, 10), 1658 => to_unsigned(436, 10), 1659 => to_unsigned(903, 10), 1660 => to_unsigned(71, 10), 1661 => to_unsigned(700, 10), 1662 => to_unsigned(775, 10), 1663 => to_unsigned(206, 10), 1664 => to_unsigned(902, 10), 1665 => to_unsigned(808, 10), 1666 => to_unsigned(463, 10), 1667 => to_unsigned(390, 10), 1668 => to_unsigned(837, 10), 1669 => to_unsigned(902, 10), 1670 => to_unsigned(727, 10), 1671 => to_unsigned(278, 10), 1672 => to_unsigned(306, 10), 1673 => to_unsigned(732, 10), 1674 => to_unsigned(75, 10), 1675 => to_unsigned(936, 10), 1676 => to_unsigned(903, 10), 1677 => to_unsigned(547, 10), 1678 => to_unsigned(658, 10), 1679 => to_unsigned(944, 10), 1680 => to_unsigned(766, 10), 1681 => to_unsigned(783, 10), 1682 => to_unsigned(139, 10), 1683 => to_unsigned(466, 10), 1684 => to_unsigned(196, 10), 1685 => to_unsigned(888, 10), 1686 => to_unsigned(731, 10), 1687 => to_unsigned(628, 10), 1688 => to_unsigned(65, 10), 1689 => to_unsigned(967, 10), 1690 => to_unsigned(19, 10), 1691 => to_unsigned(459, 10), 1692 => to_unsigned(710, 10), 1693 => to_unsigned(480, 10), 1694 => to_unsigned(581, 10), 1695 => to_unsigned(813, 10), 1696 => to_unsigned(679, 10), 1697 => to_unsigned(116, 10), 1698 => to_unsigned(851, 10), 1699 => to_unsigned(766, 10), 1700 => to_unsigned(68, 10), 1701 => to_unsigned(405, 10), 1702 => to_unsigned(668, 10), 1703 => to_unsigned(177, 10), 1704 => to_unsigned(920, 10), 1705 => to_unsigned(870, 10), 1706 => to_unsigned(139, 10), 1707 => to_unsigned(885, 10), 1708 => to_unsigned(467, 10), 1709 => to_unsigned(737, 10), 1710 => to_unsigned(44, 10), 1711 => to_unsigned(231, 10), 1712 => to_unsigned(463, 10), 1713 => to_unsigned(654, 10), 1714 => to_unsigned(403, 10), 1715 => to_unsigned(296, 10), 1716 => to_unsigned(996, 10), 1717 => to_unsigned(845, 10), 1718 => to_unsigned(700, 10), 1719 => to_unsigned(1000, 10), 1720 => to_unsigned(250, 10), 1721 => to_unsigned(361, 10), 1722 => to_unsigned(50, 10), 1723 => to_unsigned(308, 10), 1724 => to_unsigned(893, 10), 1725 => to_unsigned(858, 10), 1726 => to_unsigned(440, 10), 1727 => to_unsigned(351, 10), 1728 => to_unsigned(946, 10), 1729 => to_unsigned(679, 10), 1730 => to_unsigned(167, 10), 1731 => to_unsigned(955, 10), 1732 => to_unsigned(427, 10), 1733 => to_unsigned(165, 10), 1734 => to_unsigned(775, 10), 1735 => to_unsigned(440, 10), 1736 => to_unsigned(76, 10), 1737 => to_unsigned(426, 10), 1738 => to_unsigned(609, 10), 1739 => to_unsigned(80, 10), 1740 => to_unsigned(530, 10), 1741 => to_unsigned(482, 10), 1742 => to_unsigned(433, 10), 1743 => to_unsigned(838, 10), 1744 => to_unsigned(601, 10), 1745 => to_unsigned(767, 10), 1746 => to_unsigned(459, 10), 1747 => to_unsigned(597, 10), 1748 => to_unsigned(739, 10), 1749 => to_unsigned(185, 10), 1750 => to_unsigned(211, 10), 1751 => to_unsigned(109, 10), 1752 => to_unsigned(411, 10), 1753 => to_unsigned(198, 10), 1754 => to_unsigned(835, 10), 1755 => to_unsigned(512, 10), 1756 => to_unsigned(629, 10), 1757 => to_unsigned(267, 10), 1758 => to_unsigned(708, 10), 1759 => to_unsigned(703, 10), 1760 => to_unsigned(666, 10), 1761 => to_unsigned(613, 10), 1762 => to_unsigned(588, 10), 1763 => to_unsigned(502, 10), 1764 => to_unsigned(895, 10), 1765 => to_unsigned(962, 10), 1766 => to_unsigned(753, 10), 1767 => to_unsigned(950, 10), 1768 => to_unsigned(942, 10), 1769 => to_unsigned(311, 10), 1770 => to_unsigned(246, 10), 1771 => to_unsigned(439, 10), 1772 => to_unsigned(127, 10), 1773 => to_unsigned(438, 10), 1774 => to_unsigned(617, 10), 1775 => to_unsigned(727, 10), 1776 => to_unsigned(270, 10), 1777 => to_unsigned(613, 10), 1778 => to_unsigned(112, 10), 1779 => to_unsigned(926, 10), 1780 => to_unsigned(518, 10), 1781 => to_unsigned(397, 10), 1782 => to_unsigned(787, 10), 1783 => to_unsigned(937, 10), 1784 => to_unsigned(619, 10), 1785 => to_unsigned(703, 10), 1786 => to_unsigned(149, 10), 1787 => to_unsigned(453, 10), 1788 => to_unsigned(35, 10), 1789 => to_unsigned(399, 10), 1790 => to_unsigned(746, 10), 1791 => to_unsigned(870, 10), 1792 => to_unsigned(166, 10), 1793 => to_unsigned(547, 10), 1794 => to_unsigned(6, 10), 1795 => to_unsigned(188, 10), 1796 => to_unsigned(149, 10), 1797 => to_unsigned(250, 10), 1798 => to_unsigned(45, 10), 1799 => to_unsigned(717, 10), 1800 => to_unsigned(983, 10), 1801 => to_unsigned(351, 10), 1802 => to_unsigned(561, 10), 1803 => to_unsigned(541, 10), 1804 => to_unsigned(616, 10), 1805 => to_unsigned(737, 10), 1806 => to_unsigned(829, 10), 1807 => to_unsigned(543, 10), 1808 => to_unsigned(232, 10), 1809 => to_unsigned(474, 10), 1810 => to_unsigned(801, 10), 1811 => to_unsigned(213, 10), 1812 => to_unsigned(400, 10), 1813 => to_unsigned(520, 10), 1814 => to_unsigned(368, 10), 1815 => to_unsigned(511, 10), 1816 => to_unsigned(204, 10), 1817 => to_unsigned(807, 10), 1818 => to_unsigned(434, 10), 1819 => to_unsigned(908, 10), 1820 => to_unsigned(200, 10), 1821 => to_unsigned(667, 10), 1822 => to_unsigned(224, 10), 1823 => to_unsigned(170, 10), 1824 => to_unsigned(836, 10), 1825 => to_unsigned(428, 10), 1826 => to_unsigned(97, 10), 1827 => to_unsigned(490, 10), 1828 => to_unsigned(68, 10), 1829 => to_unsigned(831, 10), 1830 => to_unsigned(554, 10), 1831 => to_unsigned(497, 10), 1832 => to_unsigned(918, 10), 1833 => to_unsigned(336, 10), 1834 => to_unsigned(56, 10), 1835 => to_unsigned(592, 10), 1836 => to_unsigned(987, 10), 1837 => to_unsigned(844, 10), 1838 => to_unsigned(18, 10), 1839 => to_unsigned(650, 10), 1840 => to_unsigned(415, 10), 1841 => to_unsigned(1017, 10), 1842 => to_unsigned(316, 10), 1843 => to_unsigned(483, 10), 1844 => to_unsigned(519, 10), 1845 => to_unsigned(934, 10), 1846 => to_unsigned(90, 10), 1847 => to_unsigned(449, 10), 1848 => to_unsigned(465, 10), 1849 => to_unsigned(777, 10), 1850 => to_unsigned(810, 10), 1851 => to_unsigned(707, 10), 1852 => to_unsigned(472, 10), 1853 => to_unsigned(103, 10), 1854 => to_unsigned(647, 10), 1855 => to_unsigned(387, 10), 1856 => to_unsigned(273, 10), 1857 => to_unsigned(785, 10), 1858 => to_unsigned(864, 10), 1859 => to_unsigned(644, 10), 1860 => to_unsigned(227, 10), 1861 => to_unsigned(11, 10), 1862 => to_unsigned(463, 10), 1863 => to_unsigned(856, 10), 1864 => to_unsigned(866, 10), 1865 => to_unsigned(864, 10), 1866 => to_unsigned(264, 10), 1867 => to_unsigned(968, 10), 1868 => to_unsigned(991, 10), 1869 => to_unsigned(878, 10), 1870 => to_unsigned(615, 10), 1871 => to_unsigned(220, 10), 1872 => to_unsigned(500, 10), 1873 => to_unsigned(321, 10), 1874 => to_unsigned(98, 10), 1875 => to_unsigned(638, 10), 1876 => to_unsigned(454, 10), 1877 => to_unsigned(419, 10), 1878 => to_unsigned(224, 10), 1879 => to_unsigned(713, 10), 1880 => to_unsigned(82, 10), 1881 => to_unsigned(115, 10), 1882 => to_unsigned(222, 10), 1883 => to_unsigned(853, 10), 1884 => to_unsigned(836, 10), 1885 => to_unsigned(718, 10), 1886 => to_unsigned(562, 10), 1887 => to_unsigned(150, 10), 1888 => to_unsigned(330, 10), 1889 => to_unsigned(790, 10), 1890 => to_unsigned(270, 10), 1891 => to_unsigned(102, 10), 1892 => to_unsigned(876, 10), 1893 => to_unsigned(342, 10), 1894 => to_unsigned(419, 10), 1895 => to_unsigned(334, 10), 1896 => to_unsigned(366, 10), 1897 => to_unsigned(101, 10), 1898 => to_unsigned(1005, 10), 1899 => to_unsigned(709, 10), 1900 => to_unsigned(496, 10), 1901 => to_unsigned(856, 10), 1902 => to_unsigned(141, 10), 1903 => to_unsigned(1016, 10), 1904 => to_unsigned(259, 10), 1905 => to_unsigned(425, 10), 1906 => to_unsigned(690, 10), 1907 => to_unsigned(58, 10), 1908 => to_unsigned(554, 10), 1909 => to_unsigned(9, 10), 1910 => to_unsigned(510, 10), 1911 => to_unsigned(946, 10), 1912 => to_unsigned(416, 10), 1913 => to_unsigned(936, 10), 1914 => to_unsigned(705, 10), 1915 => to_unsigned(383, 10), 1916 => to_unsigned(354, 10), 1917 => to_unsigned(453, 10), 1918 => to_unsigned(311, 10), 1919 => to_unsigned(813, 10), 1920 => to_unsigned(35, 10), 1921 => to_unsigned(149, 10), 1922 => to_unsigned(948, 10), 1923 => to_unsigned(597, 10), 1924 => to_unsigned(155, 10), 1925 => to_unsigned(269, 10), 1926 => to_unsigned(564, 10), 1927 => to_unsigned(635, 10), 1928 => to_unsigned(380, 10), 1929 => to_unsigned(712, 10), 1930 => to_unsigned(861, 10), 1931 => to_unsigned(574, 10), 1932 => to_unsigned(661, 10), 1933 => to_unsigned(954, 10), 1934 => to_unsigned(563, 10), 1935 => to_unsigned(233, 10), 1936 => to_unsigned(871, 10), 1937 => to_unsigned(1, 10), 1938 => to_unsigned(41, 10), 1939 => to_unsigned(246, 10), 1940 => to_unsigned(888, 10), 1941 => to_unsigned(330, 10), 1942 => to_unsigned(454, 10), 1943 => to_unsigned(579, 10), 1944 => to_unsigned(527, 10), 1945 => to_unsigned(1001, 10), 1946 => to_unsigned(368, 10), 1947 => to_unsigned(450, 10), 1948 => to_unsigned(308, 10), 1949 => to_unsigned(729, 10), 1950 => to_unsigned(64, 10), 1951 => to_unsigned(42, 10), 1952 => to_unsigned(691, 10), 1953 => to_unsigned(132, 10), 1954 => to_unsigned(683, 10), 1955 => to_unsigned(672, 10), 1956 => to_unsigned(528, 10), 1957 => to_unsigned(1022, 10), 1958 => to_unsigned(14, 10), 1959 => to_unsigned(601, 10), 1960 => to_unsigned(214, 10), 1961 => to_unsigned(366, 10), 1962 => to_unsigned(381, 10), 1963 => to_unsigned(916, 10), 1964 => to_unsigned(381, 10), 1965 => to_unsigned(697, 10), 1966 => to_unsigned(667, 10), 1967 => to_unsigned(259, 10), 1968 => to_unsigned(182, 10), 1969 => to_unsigned(565, 10), 1970 => to_unsigned(273, 10), 1971 => to_unsigned(465, 10), 1972 => to_unsigned(694, 10), 1973 => to_unsigned(517, 10), 1974 => to_unsigned(395, 10), 1975 => to_unsigned(863, 10), 1976 => to_unsigned(63, 10), 1977 => to_unsigned(5, 10), 1978 => to_unsigned(755, 10), 1979 => to_unsigned(230, 10), 1980 => to_unsigned(36, 10), 1981 => to_unsigned(305, 10), 1982 => to_unsigned(596, 10), 1983 => to_unsigned(908, 10), 1984 => to_unsigned(460, 10), 1985 => to_unsigned(924, 10), 1986 => to_unsigned(323, 10), 1987 => to_unsigned(591, 10), 1988 => to_unsigned(318, 10), 1989 => to_unsigned(61, 10), 1990 => to_unsigned(936, 10), 1991 => to_unsigned(198, 10), 1992 => to_unsigned(315, 10), 1993 => to_unsigned(344, 10), 1994 => to_unsigned(315, 10), 1995 => to_unsigned(826, 10), 1996 => to_unsigned(346, 10), 1997 => to_unsigned(610, 10), 1998 => to_unsigned(913, 10), 1999 => to_unsigned(838, 10), 2000 => to_unsigned(599, 10), 2001 => to_unsigned(227, 10), 2002 => to_unsigned(782, 10), 2003 => to_unsigned(119, 10), 2004 => to_unsigned(454, 10), 2005 => to_unsigned(292, 10), 2006 => to_unsigned(783, 10), 2007 => to_unsigned(110, 10), 2008 => to_unsigned(794, 10), 2009 => to_unsigned(638, 10), 2010 => to_unsigned(792, 10), 2011 => to_unsigned(898, 10), 2012 => to_unsigned(959, 10), 2013 => to_unsigned(934, 10), 2014 => to_unsigned(794, 10), 2015 => to_unsigned(458, 10), 2016 => to_unsigned(766, 10), 2017 => to_unsigned(431, 10), 2018 => to_unsigned(934, 10), 2019 => to_unsigned(1008, 10), 2020 => to_unsigned(732, 10), 2021 => to_unsigned(84, 10), 2022 => to_unsigned(632, 10), 2023 => to_unsigned(424, 10), 2024 => to_unsigned(752, 10), 2025 => to_unsigned(248, 10), 2026 => to_unsigned(923, 10), 2027 => to_unsigned(925, 10), 2028 => to_unsigned(659, 10), 2029 => to_unsigned(617, 10), 2030 => to_unsigned(280, 10), 2031 => to_unsigned(342, 10), 2032 => to_unsigned(267, 10), 2033 => to_unsigned(843, 10), 2034 => to_unsigned(42, 10), 2035 => to_unsigned(255, 10), 2036 => to_unsigned(349, 10), 2037 => to_unsigned(960, 10), 2038 => to_unsigned(604, 10), 2039 => to_unsigned(76, 10), 2040 => to_unsigned(299, 10), 2041 => to_unsigned(219, 10), 2042 => to_unsigned(605, 10), 2043 => to_unsigned(755, 10), 2044 => to_unsigned(712, 10), 2045 => to_unsigned(895, 10), 2046 => to_unsigned(413, 10), 2047 => to_unsigned(999, 10))
        ),
        2 => (
            0 => (0 => to_unsigned(904, 10), 1 => to_unsigned(350, 10), 2 => to_unsigned(231, 10), 3 => to_unsigned(865, 10), 4 => to_unsigned(651, 10), 5 => to_unsigned(324, 10), 6 => to_unsigned(147, 10), 7 => to_unsigned(879, 10), 8 => to_unsigned(630, 10), 9 => to_unsigned(373, 10), 10 => to_unsigned(955, 10), 11 => to_unsigned(170, 10), 12 => to_unsigned(708, 10), 13 => to_unsigned(886, 10), 14 => to_unsigned(754, 10), 15 => to_unsigned(843, 10), 16 => to_unsigned(343, 10), 17 => to_unsigned(151, 10), 18 => to_unsigned(579, 10), 19 => to_unsigned(820, 10), 20 => to_unsigned(210, 10), 21 => to_unsigned(370, 10), 22 => to_unsigned(51, 10), 23 => to_unsigned(975, 10), 24 => to_unsigned(199, 10), 25 => to_unsigned(324, 10), 26 => to_unsigned(465, 10), 27 => to_unsigned(927, 10), 28 => to_unsigned(985, 10), 29 => to_unsigned(41, 10), 30 => to_unsigned(857, 10), 31 => to_unsigned(806, 10), 32 => to_unsigned(587, 10), 33 => to_unsigned(443, 10), 34 => to_unsigned(879, 10), 35 => to_unsigned(467, 10), 36 => to_unsigned(751, 10), 37 => to_unsigned(593, 10), 38 => to_unsigned(662, 10), 39 => to_unsigned(392, 10), 40 => to_unsigned(961, 10), 41 => to_unsigned(622, 10), 42 => to_unsigned(9, 10), 43 => to_unsigned(53, 10), 44 => to_unsigned(835, 10), 45 => to_unsigned(165, 10), 46 => to_unsigned(857, 10), 47 => to_unsigned(732, 10), 48 => to_unsigned(601, 10), 49 => to_unsigned(622, 10), 50 => to_unsigned(319, 10), 51 => to_unsigned(365, 10), 52 => to_unsigned(767, 10), 53 => to_unsigned(858, 10), 54 => to_unsigned(213, 10), 55 => to_unsigned(671, 10), 56 => to_unsigned(274, 10), 57 => to_unsigned(357, 10), 58 => to_unsigned(489, 10), 59 => to_unsigned(869, 10), 60 => to_unsigned(807, 10), 61 => to_unsigned(970, 10), 62 => to_unsigned(662, 10), 63 => to_unsigned(325, 10), 64 => to_unsigned(836, 10), 65 => to_unsigned(97, 10), 66 => to_unsigned(505, 10), 67 => to_unsigned(744, 10), 68 => to_unsigned(490, 10), 69 => to_unsigned(349, 10), 70 => to_unsigned(300, 10), 71 => to_unsigned(182, 10), 72 => to_unsigned(148, 10), 73 => to_unsigned(965, 10), 74 => to_unsigned(122, 10), 75 => to_unsigned(111, 10), 76 => to_unsigned(655, 10), 77 => to_unsigned(880, 10), 78 => to_unsigned(804, 10), 79 => to_unsigned(29, 10), 80 => to_unsigned(245, 10), 81 => to_unsigned(718, 10), 82 => to_unsigned(239, 10), 83 => to_unsigned(689, 10), 84 => to_unsigned(169, 10), 85 => to_unsigned(116, 10), 86 => to_unsigned(608, 10), 87 => to_unsigned(752, 10), 88 => to_unsigned(730, 10), 89 => to_unsigned(870, 10), 90 => to_unsigned(630, 10), 91 => to_unsigned(379, 10), 92 => to_unsigned(704, 10), 93 => to_unsigned(665, 10), 94 => to_unsigned(26, 10), 95 => to_unsigned(15, 10), 96 => to_unsigned(646, 10), 97 => to_unsigned(292, 10), 98 => to_unsigned(237, 10), 99 => to_unsigned(15, 10), 100 => to_unsigned(263, 10), 101 => to_unsigned(804, 10), 102 => to_unsigned(199, 10), 103 => to_unsigned(93, 10), 104 => to_unsigned(760, 10), 105 => to_unsigned(609, 10), 106 => to_unsigned(582, 10), 107 => to_unsigned(534, 10), 108 => to_unsigned(25, 10), 109 => to_unsigned(99, 10), 110 => to_unsigned(550, 10), 111 => to_unsigned(585, 10), 112 => to_unsigned(457, 10), 113 => to_unsigned(320, 10), 114 => to_unsigned(544, 10), 115 => to_unsigned(109, 10), 116 => to_unsigned(172, 10), 117 => to_unsigned(677, 10), 118 => to_unsigned(92, 10), 119 => to_unsigned(330, 10), 120 => to_unsigned(22, 10), 121 => to_unsigned(200, 10), 122 => to_unsigned(837, 10), 123 => to_unsigned(465, 10), 124 => to_unsigned(787, 10), 125 => to_unsigned(56, 10), 126 => to_unsigned(411, 10), 127 => to_unsigned(562, 10), 128 => to_unsigned(124, 10), 129 => to_unsigned(980, 10), 130 => to_unsigned(334, 10), 131 => to_unsigned(726, 10), 132 => to_unsigned(982, 10), 133 => to_unsigned(909, 10), 134 => to_unsigned(134, 10), 135 => to_unsigned(638, 10), 136 => to_unsigned(223, 10), 137 => to_unsigned(415, 10), 138 => to_unsigned(264, 10), 139 => to_unsigned(202, 10), 140 => to_unsigned(400, 10), 141 => to_unsigned(197, 10), 142 => to_unsigned(976, 10), 143 => to_unsigned(378, 10), 144 => to_unsigned(456, 10), 145 => to_unsigned(842, 10), 146 => to_unsigned(833, 10), 147 => to_unsigned(646, 10), 148 => to_unsigned(652, 10), 149 => to_unsigned(576, 10), 150 => to_unsigned(324, 10), 151 => to_unsigned(447, 10), 152 => to_unsigned(185, 10), 153 => to_unsigned(957, 10), 154 => to_unsigned(319, 10), 155 => to_unsigned(165, 10), 156 => to_unsigned(1017, 10), 157 => to_unsigned(258, 10), 158 => to_unsigned(506, 10), 159 => to_unsigned(427, 10), 160 => to_unsigned(479, 10), 161 => to_unsigned(389, 10), 162 => to_unsigned(57, 10), 163 => to_unsigned(402, 10), 164 => to_unsigned(647, 10), 165 => to_unsigned(233, 10), 166 => to_unsigned(98, 10), 167 => to_unsigned(307, 10), 168 => to_unsigned(205, 10), 169 => to_unsigned(189, 10), 170 => to_unsigned(54, 10), 171 => to_unsigned(19, 10), 172 => to_unsigned(739, 10), 173 => to_unsigned(787, 10), 174 => to_unsigned(466, 10), 175 => to_unsigned(761, 10), 176 => to_unsigned(879, 10), 177 => to_unsigned(1002, 10), 178 => to_unsigned(756, 10), 179 => to_unsigned(991, 10), 180 => to_unsigned(634, 10), 181 => to_unsigned(527, 10), 182 => to_unsigned(981, 10), 183 => to_unsigned(817, 10), 184 => to_unsigned(659, 10), 185 => to_unsigned(507, 10), 186 => to_unsigned(702, 10), 187 => to_unsigned(532, 10), 188 => to_unsigned(126, 10), 189 => to_unsigned(803, 10), 190 => to_unsigned(689, 10), 191 => to_unsigned(906, 10), 192 => to_unsigned(877, 10), 193 => to_unsigned(679, 10), 194 => to_unsigned(12, 10), 195 => to_unsigned(397, 10), 196 => to_unsigned(916, 10), 197 => to_unsigned(245, 10), 198 => to_unsigned(190, 10), 199 => to_unsigned(571, 10), 200 => to_unsigned(178, 10), 201 => to_unsigned(446, 10), 202 => to_unsigned(837, 10), 203 => to_unsigned(852, 10), 204 => to_unsigned(827, 10), 205 => to_unsigned(861, 10), 206 => to_unsigned(941, 10), 207 => to_unsigned(454, 10), 208 => to_unsigned(186, 10), 209 => to_unsigned(857, 10), 210 => to_unsigned(420, 10), 211 => to_unsigned(685, 10), 212 => to_unsigned(451, 10), 213 => to_unsigned(277, 10), 214 => to_unsigned(838, 10), 215 => to_unsigned(838, 10), 216 => to_unsigned(860, 10), 217 => to_unsigned(553, 10), 218 => to_unsigned(934, 10), 219 => to_unsigned(904, 10), 220 => to_unsigned(724, 10), 221 => to_unsigned(784, 10), 222 => to_unsigned(499, 10), 223 => to_unsigned(640, 10), 224 => to_unsigned(749, 10), 225 => to_unsigned(295, 10), 226 => to_unsigned(619, 10), 227 => to_unsigned(453, 10), 228 => to_unsigned(726, 10), 229 => to_unsigned(462, 10), 230 => to_unsigned(678, 10), 231 => to_unsigned(396, 10), 232 => to_unsigned(237, 10), 233 => to_unsigned(621, 10), 234 => to_unsigned(719, 10), 235 => to_unsigned(316, 10), 236 => to_unsigned(943, 10), 237 => to_unsigned(86, 10), 238 => to_unsigned(259, 10), 239 => to_unsigned(566, 10), 240 => to_unsigned(63, 10), 241 => to_unsigned(914, 10), 242 => to_unsigned(553, 10), 243 => to_unsigned(523, 10), 244 => to_unsigned(500, 10), 245 => to_unsigned(10, 10), 246 => to_unsigned(145, 10), 247 => to_unsigned(974, 10), 248 => to_unsigned(697, 10), 249 => to_unsigned(869, 10), 250 => to_unsigned(211, 10), 251 => to_unsigned(988, 10), 252 => to_unsigned(88, 10), 253 => to_unsigned(826, 10), 254 => to_unsigned(213, 10), 255 => to_unsigned(1001, 10), 256 => to_unsigned(770, 10), 257 => to_unsigned(812, 10), 258 => to_unsigned(391, 10), 259 => to_unsigned(746, 10), 260 => to_unsigned(760, 10), 261 => to_unsigned(1018, 10), 262 => to_unsigned(325, 10), 263 => to_unsigned(761, 10), 264 => to_unsigned(871, 10), 265 => to_unsigned(840, 10), 266 => to_unsigned(183, 10), 267 => to_unsigned(685, 10), 268 => to_unsigned(354, 10), 269 => to_unsigned(652, 10), 270 => to_unsigned(798, 10), 271 => to_unsigned(322, 10), 272 => to_unsigned(242, 10), 273 => to_unsigned(210, 10), 274 => to_unsigned(273, 10), 275 => to_unsigned(507, 10), 276 => to_unsigned(952, 10), 277 => to_unsigned(199, 10), 278 => to_unsigned(931, 10), 279 => to_unsigned(396, 10), 280 => to_unsigned(554, 10), 281 => to_unsigned(1017, 10), 282 => to_unsigned(190, 10), 283 => to_unsigned(404, 10), 284 => to_unsigned(641, 10), 285 => to_unsigned(519, 10), 286 => to_unsigned(766, 10), 287 => to_unsigned(438, 10), 288 => to_unsigned(719, 10), 289 => to_unsigned(925, 10), 290 => to_unsigned(253, 10), 291 => to_unsigned(452, 10), 292 => to_unsigned(140, 10), 293 => to_unsigned(839, 10), 294 => to_unsigned(71, 10), 295 => to_unsigned(819, 10), 296 => to_unsigned(498, 10), 297 => to_unsigned(618, 10), 298 => to_unsigned(908, 10), 299 => to_unsigned(708, 10), 300 => to_unsigned(778, 10), 301 => to_unsigned(1020, 10), 302 => to_unsigned(447, 10), 303 => to_unsigned(126, 10), 304 => to_unsigned(251, 10), 305 => to_unsigned(119, 10), 306 => to_unsigned(315, 10), 307 => to_unsigned(735, 10), 308 => to_unsigned(525, 10), 309 => to_unsigned(88, 10), 310 => to_unsigned(471, 10), 311 => to_unsigned(123, 10), 312 => to_unsigned(300, 10), 313 => to_unsigned(522, 10), 314 => to_unsigned(213, 10), 315 => to_unsigned(746, 10), 316 => to_unsigned(1000, 10), 317 => to_unsigned(889, 10), 318 => to_unsigned(242, 10), 319 => to_unsigned(902, 10), 320 => to_unsigned(980, 10), 321 => to_unsigned(556, 10), 322 => to_unsigned(260, 10), 323 => to_unsigned(351, 10), 324 => to_unsigned(863, 10), 325 => to_unsigned(871, 10), 326 => to_unsigned(988, 10), 327 => to_unsigned(16, 10), 328 => to_unsigned(577, 10), 329 => to_unsigned(747, 10), 330 => to_unsigned(992, 10), 331 => to_unsigned(194, 10), 332 => to_unsigned(119, 10), 333 => to_unsigned(157, 10), 334 => to_unsigned(330, 10), 335 => to_unsigned(152, 10), 336 => to_unsigned(776, 10), 337 => to_unsigned(815, 10), 338 => to_unsigned(94, 10), 339 => to_unsigned(793, 10), 340 => to_unsigned(521, 10), 341 => to_unsigned(328, 10), 342 => to_unsigned(764, 10), 343 => to_unsigned(759, 10), 344 => to_unsigned(195, 10), 345 => to_unsigned(170, 10), 346 => to_unsigned(485, 10), 347 => to_unsigned(269, 10), 348 => to_unsigned(31, 10), 349 => to_unsigned(46, 10), 350 => to_unsigned(661, 10), 351 => to_unsigned(384, 10), 352 => to_unsigned(637, 10), 353 => to_unsigned(963, 10), 354 => to_unsigned(763, 10), 355 => to_unsigned(826, 10), 356 => to_unsigned(838, 10), 357 => to_unsigned(460, 10), 358 => to_unsigned(856, 10), 359 => to_unsigned(382, 10), 360 => to_unsigned(309, 10), 361 => to_unsigned(15, 10), 362 => to_unsigned(900, 10), 363 => to_unsigned(440, 10), 364 => to_unsigned(393, 10), 365 => to_unsigned(541, 10), 366 => to_unsigned(29, 10), 367 => to_unsigned(538, 10), 368 => to_unsigned(4, 10), 369 => to_unsigned(155, 10), 370 => to_unsigned(541, 10), 371 => to_unsigned(400, 10), 372 => to_unsigned(112, 10), 373 => to_unsigned(270, 10), 374 => to_unsigned(900, 10), 375 => to_unsigned(585, 10), 376 => to_unsigned(462, 10), 377 => to_unsigned(267, 10), 378 => to_unsigned(23, 10), 379 => to_unsigned(754, 10), 380 => to_unsigned(246, 10), 381 => to_unsigned(88, 10), 382 => to_unsigned(149, 10), 383 => to_unsigned(617, 10), 384 => to_unsigned(193, 10), 385 => to_unsigned(32, 10), 386 => to_unsigned(716, 10), 387 => to_unsigned(512, 10), 388 => to_unsigned(479, 10), 389 => to_unsigned(36, 10), 390 => to_unsigned(667, 10), 391 => to_unsigned(516, 10), 392 => to_unsigned(572, 10), 393 => to_unsigned(950, 10), 394 => to_unsigned(111, 10), 395 => to_unsigned(294, 10), 396 => to_unsigned(434, 10), 397 => to_unsigned(418, 10), 398 => to_unsigned(323, 10), 399 => to_unsigned(595, 10), 400 => to_unsigned(358, 10), 401 => to_unsigned(996, 10), 402 => to_unsigned(565, 10), 403 => to_unsigned(445, 10), 404 => to_unsigned(881, 10), 405 => to_unsigned(379, 10), 406 => to_unsigned(467, 10), 407 => to_unsigned(772, 10), 408 => to_unsigned(857, 10), 409 => to_unsigned(341, 10), 410 => to_unsigned(995, 10), 411 => to_unsigned(932, 10), 412 => to_unsigned(477, 10), 413 => to_unsigned(274, 10), 414 => to_unsigned(257, 10), 415 => to_unsigned(955, 10), 416 => to_unsigned(154, 10), 417 => to_unsigned(628, 10), 418 => to_unsigned(285, 10), 419 => to_unsigned(664, 10), 420 => to_unsigned(54, 10), 421 => to_unsigned(450, 10), 422 => to_unsigned(49, 10), 423 => to_unsigned(219, 10), 424 => to_unsigned(690, 10), 425 => to_unsigned(888, 10), 426 => to_unsigned(877, 10), 427 => to_unsigned(93, 10), 428 => to_unsigned(122, 10), 429 => to_unsigned(331, 10), 430 => to_unsigned(566, 10), 431 => to_unsigned(512, 10), 432 => to_unsigned(712, 10), 433 => to_unsigned(219, 10), 434 => to_unsigned(264, 10), 435 => to_unsigned(678, 10), 436 => to_unsigned(746, 10), 437 => to_unsigned(692, 10), 438 => to_unsigned(336, 10), 439 => to_unsigned(653, 10), 440 => to_unsigned(696, 10), 441 => to_unsigned(675, 10), 442 => to_unsigned(155, 10), 443 => to_unsigned(23, 10), 444 => to_unsigned(943, 10), 445 => to_unsigned(885, 10), 446 => to_unsigned(911, 10), 447 => to_unsigned(178, 10), 448 => to_unsigned(888, 10), 449 => to_unsigned(317, 10), 450 => to_unsigned(648, 10), 451 => to_unsigned(721, 10), 452 => to_unsigned(464, 10), 453 => to_unsigned(920, 10), 454 => to_unsigned(244, 10), 455 => to_unsigned(567, 10), 456 => to_unsigned(270, 10), 457 => to_unsigned(336, 10), 458 => to_unsigned(840, 10), 459 => to_unsigned(761, 10), 460 => to_unsigned(571, 10), 461 => to_unsigned(87, 10), 462 => to_unsigned(917, 10), 463 => to_unsigned(202, 10), 464 => to_unsigned(929, 10), 465 => to_unsigned(824, 10), 466 => to_unsigned(992, 10), 467 => to_unsigned(549, 10), 468 => to_unsigned(742, 10), 469 => to_unsigned(110, 10), 470 => to_unsigned(975, 10), 471 => to_unsigned(433, 10), 472 => to_unsigned(617, 10), 473 => to_unsigned(204, 10), 474 => to_unsigned(178, 10), 475 => to_unsigned(593, 10), 476 => to_unsigned(459, 10), 477 => to_unsigned(804, 10), 478 => to_unsigned(824, 10), 479 => to_unsigned(154, 10), 480 => to_unsigned(730, 10), 481 => to_unsigned(635, 10), 482 => to_unsigned(613, 10), 483 => to_unsigned(937, 10), 484 => to_unsigned(534, 10), 485 => to_unsigned(454, 10), 486 => to_unsigned(660, 10), 487 => to_unsigned(826, 10), 488 => to_unsigned(395, 10), 489 => to_unsigned(808, 10), 490 => to_unsigned(193, 10), 491 => to_unsigned(62, 10), 492 => to_unsigned(281, 10), 493 => to_unsigned(456, 10), 494 => to_unsigned(1001, 10), 495 => to_unsigned(196, 10), 496 => to_unsigned(635, 10), 497 => to_unsigned(127, 10), 498 => to_unsigned(619, 10), 499 => to_unsigned(570, 10), 500 => to_unsigned(389, 10), 501 => to_unsigned(834, 10), 502 => to_unsigned(692, 10), 503 => to_unsigned(727, 10), 504 => to_unsigned(204, 10), 505 => to_unsigned(442, 10), 506 => to_unsigned(340, 10), 507 => to_unsigned(696, 10), 508 => to_unsigned(125, 10), 509 => to_unsigned(61, 10), 510 => to_unsigned(894, 10), 511 => to_unsigned(296, 10), 512 => to_unsigned(237, 10), 513 => to_unsigned(190, 10), 514 => to_unsigned(971, 10), 515 => to_unsigned(919, 10), 516 => to_unsigned(896, 10), 517 => to_unsigned(873, 10), 518 => to_unsigned(755, 10), 519 => to_unsigned(346, 10), 520 => to_unsigned(729, 10), 521 => to_unsigned(164, 10), 522 => to_unsigned(430, 10), 523 => to_unsigned(313, 10), 524 => to_unsigned(1023, 10), 525 => to_unsigned(541, 10), 526 => to_unsigned(233, 10), 527 => to_unsigned(533, 10), 528 => to_unsigned(650, 10), 529 => to_unsigned(503, 10), 530 => to_unsigned(884, 10), 531 => to_unsigned(976, 10), 532 => to_unsigned(752, 10), 533 => to_unsigned(473, 10), 534 => to_unsigned(769, 10), 535 => to_unsigned(114, 10), 536 => to_unsigned(365, 10), 537 => to_unsigned(307, 10), 538 => to_unsigned(170, 10), 539 => to_unsigned(649, 10), 540 => to_unsigned(1010, 10), 541 => to_unsigned(70, 10), 542 => to_unsigned(181, 10), 543 => to_unsigned(70, 10), 544 => to_unsigned(267, 10), 545 => to_unsigned(577, 10), 546 => to_unsigned(199, 10), 547 => to_unsigned(340, 10), 548 => to_unsigned(105, 10), 549 => to_unsigned(739, 10), 550 => to_unsigned(807, 10), 551 => to_unsigned(494, 10), 552 => to_unsigned(642, 10), 553 => to_unsigned(547, 10), 554 => to_unsigned(129, 10), 555 => to_unsigned(651, 10), 556 => to_unsigned(912, 10), 557 => to_unsigned(249, 10), 558 => to_unsigned(990, 10), 559 => to_unsigned(943, 10), 560 => to_unsigned(400, 10), 561 => to_unsigned(978, 10), 562 => to_unsigned(747, 10), 563 => to_unsigned(1017, 10), 564 => to_unsigned(485, 10), 565 => to_unsigned(331, 10), 566 => to_unsigned(315, 10), 567 => to_unsigned(729, 10), 568 => to_unsigned(536, 10), 569 => to_unsigned(446, 10), 570 => to_unsigned(233, 10), 571 => to_unsigned(107, 10), 572 => to_unsigned(281, 10), 573 => to_unsigned(218, 10), 574 => to_unsigned(1012, 10), 575 => to_unsigned(145, 10), 576 => to_unsigned(41, 10), 577 => to_unsigned(342, 10), 578 => to_unsigned(910, 10), 579 => to_unsigned(324, 10), 580 => to_unsigned(531, 10), 581 => to_unsigned(715, 10), 582 => to_unsigned(607, 10), 583 => to_unsigned(371, 10), 584 => to_unsigned(756, 10), 585 => to_unsigned(133, 10), 586 => to_unsigned(357, 10), 587 => to_unsigned(757, 10), 588 => to_unsigned(816, 10), 589 => to_unsigned(451, 10), 590 => to_unsigned(609, 10), 591 => to_unsigned(497, 10), 592 => to_unsigned(622, 10), 593 => to_unsigned(760, 10), 594 => to_unsigned(497, 10), 595 => to_unsigned(30, 10), 596 => to_unsigned(386, 10), 597 => to_unsigned(870, 10), 598 => to_unsigned(311, 10), 599 => to_unsigned(438, 10), 600 => to_unsigned(55, 10), 601 => to_unsigned(24, 10), 602 => to_unsigned(503, 10), 603 => to_unsigned(14, 10), 604 => to_unsigned(769, 10), 605 => to_unsigned(950, 10), 606 => to_unsigned(180, 10), 607 => to_unsigned(660, 10), 608 => to_unsigned(661, 10), 609 => to_unsigned(327, 10), 610 => to_unsigned(406, 10), 611 => to_unsigned(89, 10), 612 => to_unsigned(900, 10), 613 => to_unsigned(507, 10), 614 => to_unsigned(336, 10), 615 => to_unsigned(501, 10), 616 => to_unsigned(39, 10), 617 => to_unsigned(534, 10), 618 => to_unsigned(300, 10), 619 => to_unsigned(616, 10), 620 => to_unsigned(616, 10), 621 => to_unsigned(680, 10), 622 => to_unsigned(577, 10), 623 => to_unsigned(968, 10), 624 => to_unsigned(115, 10), 625 => to_unsigned(42, 10), 626 => to_unsigned(245, 10), 627 => to_unsigned(648, 10), 628 => to_unsigned(439, 10), 629 => to_unsigned(455, 10), 630 => to_unsigned(319, 10), 631 => to_unsigned(540, 10), 632 => to_unsigned(616, 10), 633 => to_unsigned(358, 10), 634 => to_unsigned(516, 10), 635 => to_unsigned(340, 10), 636 => to_unsigned(611, 10), 637 => to_unsigned(438, 10), 638 => to_unsigned(491, 10), 639 => to_unsigned(628, 10), 640 => to_unsigned(250, 10), 641 => to_unsigned(839, 10), 642 => to_unsigned(937, 10), 643 => to_unsigned(205, 10), 644 => to_unsigned(957, 10), 645 => to_unsigned(568, 10), 646 => to_unsigned(659, 10), 647 => to_unsigned(32, 10), 648 => to_unsigned(73, 10), 649 => to_unsigned(94, 10), 650 => to_unsigned(631, 10), 651 => to_unsigned(933, 10), 652 => to_unsigned(108, 10), 653 => to_unsigned(383, 10), 654 => to_unsigned(845, 10), 655 => to_unsigned(238, 10), 656 => to_unsigned(350, 10), 657 => to_unsigned(833, 10), 658 => to_unsigned(588, 10), 659 => to_unsigned(1014, 10), 660 => to_unsigned(132, 10), 661 => to_unsigned(89, 10), 662 => to_unsigned(362, 10), 663 => to_unsigned(27, 10), 664 => to_unsigned(9, 10), 665 => to_unsigned(72, 10), 666 => to_unsigned(445, 10), 667 => to_unsigned(355, 10), 668 => to_unsigned(408, 10), 669 => to_unsigned(481, 10), 670 => to_unsigned(521, 10), 671 => to_unsigned(383, 10), 672 => to_unsigned(113, 10), 673 => to_unsigned(580, 10), 674 => to_unsigned(785, 10), 675 => to_unsigned(1010, 10), 676 => to_unsigned(490, 10), 677 => to_unsigned(66, 10), 678 => to_unsigned(917, 10), 679 => to_unsigned(118, 10), 680 => to_unsigned(267, 10), 681 => to_unsigned(610, 10), 682 => to_unsigned(796, 10), 683 => to_unsigned(125, 10), 684 => to_unsigned(989, 10), 685 => to_unsigned(483, 10), 686 => to_unsigned(660, 10), 687 => to_unsigned(67, 10), 688 => to_unsigned(191, 10), 689 => to_unsigned(926, 10), 690 => to_unsigned(496, 10), 691 => to_unsigned(156, 10), 692 => to_unsigned(741, 10), 693 => to_unsigned(474, 10), 694 => to_unsigned(724, 10), 695 => to_unsigned(35, 10), 696 => to_unsigned(690, 10), 697 => to_unsigned(558, 10), 698 => to_unsigned(83, 10), 699 => to_unsigned(413, 10), 700 => to_unsigned(738, 10), 701 => to_unsigned(606, 10), 702 => to_unsigned(48, 10), 703 => to_unsigned(284, 10), 704 => to_unsigned(975, 10), 705 => to_unsigned(164, 10), 706 => to_unsigned(625, 10), 707 => to_unsigned(778, 10), 708 => to_unsigned(965, 10), 709 => to_unsigned(659, 10), 710 => to_unsigned(130, 10), 711 => to_unsigned(381, 10), 712 => to_unsigned(241, 10), 713 => to_unsigned(710, 10), 714 => to_unsigned(960, 10), 715 => to_unsigned(57, 10), 716 => to_unsigned(158, 10), 717 => to_unsigned(900, 10), 718 => to_unsigned(512, 10), 719 => to_unsigned(854, 10), 720 => to_unsigned(983, 10), 721 => to_unsigned(10, 10), 722 => to_unsigned(902, 10), 723 => to_unsigned(958, 10), 724 => to_unsigned(992, 10), 725 => to_unsigned(323, 10), 726 => to_unsigned(548, 10), 727 => to_unsigned(737, 10), 728 => to_unsigned(638, 10), 729 => to_unsigned(224, 10), 730 => to_unsigned(6, 10), 731 => to_unsigned(709, 10), 732 => to_unsigned(101, 10), 733 => to_unsigned(831, 10), 734 => to_unsigned(79, 10), 735 => to_unsigned(483, 10), 736 => to_unsigned(857, 10), 737 => to_unsigned(19, 10), 738 => to_unsigned(385, 10), 739 => to_unsigned(1003, 10), 740 => to_unsigned(536, 10), 741 => to_unsigned(630, 10), 742 => to_unsigned(213, 10), 743 => to_unsigned(226, 10), 744 => to_unsigned(654, 10), 745 => to_unsigned(628, 10), 746 => to_unsigned(386, 10), 747 => to_unsigned(583, 10), 748 => to_unsigned(101, 10), 749 => to_unsigned(279, 10), 750 => to_unsigned(694, 10), 751 => to_unsigned(422, 10), 752 => to_unsigned(287, 10), 753 => to_unsigned(705, 10), 754 => to_unsigned(1023, 10), 755 => to_unsigned(103, 10), 756 => to_unsigned(443, 10), 757 => to_unsigned(762, 10), 758 => to_unsigned(17, 10), 759 => to_unsigned(52, 10), 760 => to_unsigned(461, 10), 761 => to_unsigned(798, 10), 762 => to_unsigned(867, 10), 763 => to_unsigned(313, 10), 764 => to_unsigned(854, 10), 765 => to_unsigned(211, 10), 766 => to_unsigned(251, 10), 767 => to_unsigned(412, 10), 768 => to_unsigned(326, 10), 769 => to_unsigned(193, 10), 770 => to_unsigned(505, 10), 771 => to_unsigned(5, 10), 772 => to_unsigned(523, 10), 773 => to_unsigned(53, 10), 774 => to_unsigned(920, 10), 775 => to_unsigned(346, 10), 776 => to_unsigned(760, 10), 777 => to_unsigned(815, 10), 778 => to_unsigned(321, 10), 779 => to_unsigned(869, 10), 780 => to_unsigned(682, 10), 781 => to_unsigned(447, 10), 782 => to_unsigned(160, 10), 783 => to_unsigned(523, 10), 784 => to_unsigned(914, 10), 785 => to_unsigned(639, 10), 786 => to_unsigned(536, 10), 787 => to_unsigned(132, 10), 788 => to_unsigned(903, 10), 789 => to_unsigned(544, 10), 790 => to_unsigned(399, 10), 791 => to_unsigned(1, 10), 792 => to_unsigned(369, 10), 793 => to_unsigned(88, 10), 794 => to_unsigned(933, 10), 795 => to_unsigned(886, 10), 796 => to_unsigned(593, 10), 797 => to_unsigned(372, 10), 798 => to_unsigned(31, 10), 799 => to_unsigned(927, 10), 800 => to_unsigned(456, 10), 801 => to_unsigned(961, 10), 802 => to_unsigned(372, 10), 803 => to_unsigned(753, 10), 804 => to_unsigned(52, 10), 805 => to_unsigned(256, 10), 806 => to_unsigned(669, 10), 807 => to_unsigned(824, 10), 808 => to_unsigned(897, 10), 809 => to_unsigned(153, 10), 810 => to_unsigned(745, 10), 811 => to_unsigned(834, 10), 812 => to_unsigned(44, 10), 813 => to_unsigned(786, 10), 814 => to_unsigned(724, 10), 815 => to_unsigned(231, 10), 816 => to_unsigned(993, 10), 817 => to_unsigned(509, 10), 818 => to_unsigned(819, 10), 819 => to_unsigned(845, 10), 820 => to_unsigned(287, 10), 821 => to_unsigned(885, 10), 822 => to_unsigned(132, 10), 823 => to_unsigned(680, 10), 824 => to_unsigned(995, 10), 825 => to_unsigned(376, 10), 826 => to_unsigned(119, 10), 827 => to_unsigned(883, 10), 828 => to_unsigned(610, 10), 829 => to_unsigned(382, 10), 830 => to_unsigned(407, 10), 831 => to_unsigned(606, 10), 832 => to_unsigned(312, 10), 833 => to_unsigned(441, 10), 834 => to_unsigned(829, 10), 835 => to_unsigned(3, 10), 836 => to_unsigned(333, 10), 837 => to_unsigned(686, 10), 838 => to_unsigned(283, 10), 839 => to_unsigned(494, 10), 840 => to_unsigned(96, 10), 841 => to_unsigned(257, 10), 842 => to_unsigned(3, 10), 843 => to_unsigned(98, 10), 844 => to_unsigned(740, 10), 845 => to_unsigned(267, 10), 846 => to_unsigned(699, 10), 847 => to_unsigned(103, 10), 848 => to_unsigned(470, 10), 849 => to_unsigned(401, 10), 850 => to_unsigned(156, 10), 851 => to_unsigned(679, 10), 852 => to_unsigned(66, 10), 853 => to_unsigned(820, 10), 854 => to_unsigned(857, 10), 855 => to_unsigned(656, 10), 856 => to_unsigned(684, 10), 857 => to_unsigned(623, 10), 858 => to_unsigned(752, 10), 859 => to_unsigned(118, 10), 860 => to_unsigned(343, 10), 861 => to_unsigned(245, 10), 862 => to_unsigned(746, 10), 863 => to_unsigned(132, 10), 864 => to_unsigned(844, 10), 865 => to_unsigned(455, 10), 866 => to_unsigned(1002, 10), 867 => to_unsigned(535, 10), 868 => to_unsigned(88, 10), 869 => to_unsigned(447, 10), 870 => to_unsigned(209, 10), 871 => to_unsigned(756, 10), 872 => to_unsigned(939, 10), 873 => to_unsigned(732, 10), 874 => to_unsigned(453, 10), 875 => to_unsigned(362, 10), 876 => to_unsigned(342, 10), 877 => to_unsigned(912, 10), 878 => to_unsigned(815, 10), 879 => to_unsigned(1018, 10), 880 => to_unsigned(617, 10), 881 => to_unsigned(642, 10), 882 => to_unsigned(709, 10), 883 => to_unsigned(683, 10), 884 => to_unsigned(406, 10), 885 => to_unsigned(753, 10), 886 => to_unsigned(275, 10), 887 => to_unsigned(724, 10), 888 => to_unsigned(550, 10), 889 => to_unsigned(338, 10), 890 => to_unsigned(649, 10), 891 => to_unsigned(87, 10), 892 => to_unsigned(835, 10), 893 => to_unsigned(430, 10), 894 => to_unsigned(134, 10), 895 => to_unsigned(140, 10), 896 => to_unsigned(235, 10), 897 => to_unsigned(137, 10), 898 => to_unsigned(26, 10), 899 => to_unsigned(1005, 10), 900 => to_unsigned(457, 10), 901 => to_unsigned(651, 10), 902 => to_unsigned(453, 10), 903 => to_unsigned(256, 10), 904 => to_unsigned(967, 10), 905 => to_unsigned(438, 10), 906 => to_unsigned(829, 10), 907 => to_unsigned(469, 10), 908 => to_unsigned(713, 10), 909 => to_unsigned(412, 10), 910 => to_unsigned(80, 10), 911 => to_unsigned(46, 10), 912 => to_unsigned(308, 10), 913 => to_unsigned(980, 10), 914 => to_unsigned(635, 10), 915 => to_unsigned(808, 10), 916 => to_unsigned(885, 10), 917 => to_unsigned(606, 10), 918 => to_unsigned(526, 10), 919 => to_unsigned(552, 10), 920 => to_unsigned(980, 10), 921 => to_unsigned(385, 10), 922 => to_unsigned(684, 10), 923 => to_unsigned(540, 10), 924 => to_unsigned(505, 10), 925 => to_unsigned(395, 10), 926 => to_unsigned(997, 10), 927 => to_unsigned(701, 10), 928 => to_unsigned(507, 10), 929 => to_unsigned(706, 10), 930 => to_unsigned(289, 10), 931 => to_unsigned(635, 10), 932 => to_unsigned(536, 10), 933 => to_unsigned(260, 10), 934 => to_unsigned(932, 10), 935 => to_unsigned(178, 10), 936 => to_unsigned(828, 10), 937 => to_unsigned(92, 10), 938 => to_unsigned(645, 10), 939 => to_unsigned(989, 10), 940 => to_unsigned(434, 10), 941 => to_unsigned(599, 10), 942 => to_unsigned(293, 10), 943 => to_unsigned(519, 10), 944 => to_unsigned(718, 10), 945 => to_unsigned(96, 10), 946 => to_unsigned(866, 10), 947 => to_unsigned(621, 10), 948 => to_unsigned(707, 10), 949 => to_unsigned(360, 10), 950 => to_unsigned(966, 10), 951 => to_unsigned(100, 10), 952 => to_unsigned(748, 10), 953 => to_unsigned(929, 10), 954 => to_unsigned(446, 10), 955 => to_unsigned(572, 10), 956 => to_unsigned(244, 10), 957 => to_unsigned(389, 10), 958 => to_unsigned(644, 10), 959 => to_unsigned(363, 10), 960 => to_unsigned(172, 10), 961 => to_unsigned(916, 10), 962 => to_unsigned(34, 10), 963 => to_unsigned(313, 10), 964 => to_unsigned(1019, 10), 965 => to_unsigned(126, 10), 966 => to_unsigned(352, 10), 967 => to_unsigned(626, 10), 968 => to_unsigned(151, 10), 969 => to_unsigned(340, 10), 970 => to_unsigned(780, 10), 971 => to_unsigned(501, 10), 972 => to_unsigned(88, 10), 973 => to_unsigned(142, 10), 974 => to_unsigned(462, 10), 975 => to_unsigned(378, 10), 976 => to_unsigned(534, 10), 977 => to_unsigned(134, 10), 978 => to_unsigned(1017, 10), 979 => to_unsigned(868, 10), 980 => to_unsigned(188, 10), 981 => to_unsigned(509, 10), 982 => to_unsigned(241, 10), 983 => to_unsigned(758, 10), 984 => to_unsigned(372, 10), 985 => to_unsigned(812, 10), 986 => to_unsigned(852, 10), 987 => to_unsigned(619, 10), 988 => to_unsigned(648, 10), 989 => to_unsigned(379, 10), 990 => to_unsigned(315, 10), 991 => to_unsigned(575, 10), 992 => to_unsigned(468, 10), 993 => to_unsigned(200, 10), 994 => to_unsigned(322, 10), 995 => to_unsigned(803, 10), 996 => to_unsigned(441, 10), 997 => to_unsigned(461, 10), 998 => to_unsigned(233, 10), 999 => to_unsigned(332, 10), 1000 => to_unsigned(1005, 10), 1001 => to_unsigned(370, 10), 1002 => to_unsigned(825, 10), 1003 => to_unsigned(562, 10), 1004 => to_unsigned(278, 10), 1005 => to_unsigned(132, 10), 1006 => to_unsigned(42, 10), 1007 => to_unsigned(954, 10), 1008 => to_unsigned(42, 10), 1009 => to_unsigned(488, 10), 1010 => to_unsigned(493, 10), 1011 => to_unsigned(875, 10), 1012 => to_unsigned(544, 10), 1013 => to_unsigned(374, 10), 1014 => to_unsigned(965, 10), 1015 => to_unsigned(619, 10), 1016 => to_unsigned(136, 10), 1017 => to_unsigned(704, 10), 1018 => to_unsigned(303, 10), 1019 => to_unsigned(348, 10), 1020 => to_unsigned(695, 10), 1021 => to_unsigned(856, 10), 1022 => to_unsigned(916, 10), 1023 => to_unsigned(267, 10), 1024 => to_unsigned(385, 10), 1025 => to_unsigned(601, 10), 1026 => to_unsigned(311, 10), 1027 => to_unsigned(879, 10), 1028 => to_unsigned(37, 10), 1029 => to_unsigned(928, 10), 1030 => to_unsigned(305, 10), 1031 => to_unsigned(75, 10), 1032 => to_unsigned(325, 10), 1033 => to_unsigned(400, 10), 1034 => to_unsigned(808, 10), 1035 => to_unsigned(908, 10), 1036 => to_unsigned(496, 10), 1037 => to_unsigned(983, 10), 1038 => to_unsigned(235, 10), 1039 => to_unsigned(601, 10), 1040 => to_unsigned(680, 10), 1041 => to_unsigned(234, 10), 1042 => to_unsigned(833, 10), 1043 => to_unsigned(217, 10), 1044 => to_unsigned(918, 10), 1045 => to_unsigned(321, 10), 1046 => to_unsigned(183, 10), 1047 => to_unsigned(333, 10), 1048 => to_unsigned(149, 10), 1049 => to_unsigned(358, 10), 1050 => to_unsigned(124, 10), 1051 => to_unsigned(163, 10), 1052 => to_unsigned(314, 10), 1053 => to_unsigned(608, 10), 1054 => to_unsigned(143, 10), 1055 => to_unsigned(630, 10), 1056 => to_unsigned(711, 10), 1057 => to_unsigned(695, 10), 1058 => to_unsigned(393, 10), 1059 => to_unsigned(969, 10), 1060 => to_unsigned(793, 10), 1061 => to_unsigned(255, 10), 1062 => to_unsigned(754, 10), 1063 => to_unsigned(731, 10), 1064 => to_unsigned(693, 10), 1065 => to_unsigned(984, 10), 1066 => to_unsigned(738, 10), 1067 => to_unsigned(429, 10), 1068 => to_unsigned(920, 10), 1069 => to_unsigned(847, 10), 1070 => to_unsigned(514, 10), 1071 => to_unsigned(300, 10), 1072 => to_unsigned(511, 10), 1073 => to_unsigned(382, 10), 1074 => to_unsigned(772, 10), 1075 => to_unsigned(391, 10), 1076 => to_unsigned(25, 10), 1077 => to_unsigned(974, 10), 1078 => to_unsigned(925, 10), 1079 => to_unsigned(341, 10), 1080 => to_unsigned(332, 10), 1081 => to_unsigned(658, 10), 1082 => to_unsigned(502, 10), 1083 => to_unsigned(752, 10), 1084 => to_unsigned(494, 10), 1085 => to_unsigned(523, 10), 1086 => to_unsigned(869, 10), 1087 => to_unsigned(11, 10), 1088 => to_unsigned(513, 10), 1089 => to_unsigned(207, 10), 1090 => to_unsigned(756, 10), 1091 => to_unsigned(912, 10), 1092 => to_unsigned(411, 10), 1093 => to_unsigned(717, 10), 1094 => to_unsigned(679, 10), 1095 => to_unsigned(543, 10), 1096 => to_unsigned(356, 10), 1097 => to_unsigned(713, 10), 1098 => to_unsigned(679, 10), 1099 => to_unsigned(209, 10), 1100 => to_unsigned(814, 10), 1101 => to_unsigned(584, 10), 1102 => to_unsigned(548, 10), 1103 => to_unsigned(290, 10), 1104 => to_unsigned(171, 10), 1105 => to_unsigned(775, 10), 1106 => to_unsigned(122, 10), 1107 => to_unsigned(675, 10), 1108 => to_unsigned(890, 10), 1109 => to_unsigned(409, 10), 1110 => to_unsigned(395, 10), 1111 => to_unsigned(34, 10), 1112 => to_unsigned(535, 10), 1113 => to_unsigned(103, 10), 1114 => to_unsigned(444, 10), 1115 => to_unsigned(401, 10), 1116 => to_unsigned(689, 10), 1117 => to_unsigned(692, 10), 1118 => to_unsigned(981, 10), 1119 => to_unsigned(474, 10), 1120 => to_unsigned(110, 10), 1121 => to_unsigned(762, 10), 1122 => to_unsigned(203, 10), 1123 => to_unsigned(889, 10), 1124 => to_unsigned(34, 10), 1125 => to_unsigned(246, 10), 1126 => to_unsigned(130, 10), 1127 => to_unsigned(73, 10), 1128 => to_unsigned(367, 10), 1129 => to_unsigned(420, 10), 1130 => to_unsigned(637, 10), 1131 => to_unsigned(385, 10), 1132 => to_unsigned(186, 10), 1133 => to_unsigned(319, 10), 1134 => to_unsigned(311, 10), 1135 => to_unsigned(573, 10), 1136 => to_unsigned(457, 10), 1137 => to_unsigned(811, 10), 1138 => to_unsigned(843, 10), 1139 => to_unsigned(788, 10), 1140 => to_unsigned(773, 10), 1141 => to_unsigned(36, 10), 1142 => to_unsigned(619, 10), 1143 => to_unsigned(56, 10), 1144 => to_unsigned(979, 10), 1145 => to_unsigned(950, 10), 1146 => to_unsigned(711, 10), 1147 => to_unsigned(946, 10), 1148 => to_unsigned(826, 10), 1149 => to_unsigned(931, 10), 1150 => to_unsigned(6, 10), 1151 => to_unsigned(545, 10), 1152 => to_unsigned(216, 10), 1153 => to_unsigned(259, 10), 1154 => to_unsigned(729, 10), 1155 => to_unsigned(657, 10), 1156 => to_unsigned(744, 10), 1157 => to_unsigned(943, 10), 1158 => to_unsigned(588, 10), 1159 => to_unsigned(1004, 10), 1160 => to_unsigned(751, 10), 1161 => to_unsigned(305, 10), 1162 => to_unsigned(565, 10), 1163 => to_unsigned(523, 10), 1164 => to_unsigned(648, 10), 1165 => to_unsigned(1014, 10), 1166 => to_unsigned(733, 10), 1167 => to_unsigned(817, 10), 1168 => to_unsigned(536, 10), 1169 => to_unsigned(668, 10), 1170 => to_unsigned(288, 10), 1171 => to_unsigned(339, 10), 1172 => to_unsigned(302, 10), 1173 => to_unsigned(840, 10), 1174 => to_unsigned(888, 10), 1175 => to_unsigned(345, 10), 1176 => to_unsigned(144, 10), 1177 => to_unsigned(460, 10), 1178 => to_unsigned(246, 10), 1179 => to_unsigned(366, 10), 1180 => to_unsigned(163, 10), 1181 => to_unsigned(894, 10), 1182 => to_unsigned(235, 10), 1183 => to_unsigned(126, 10), 1184 => to_unsigned(615, 10), 1185 => to_unsigned(312, 10), 1186 => to_unsigned(547, 10), 1187 => to_unsigned(29, 10), 1188 => to_unsigned(846, 10), 1189 => to_unsigned(717, 10), 1190 => to_unsigned(109, 10), 1191 => to_unsigned(394, 10), 1192 => to_unsigned(912, 10), 1193 => to_unsigned(387, 10), 1194 => to_unsigned(767, 10), 1195 => to_unsigned(277, 10), 1196 => to_unsigned(542, 10), 1197 => to_unsigned(667, 10), 1198 => to_unsigned(615, 10), 1199 => to_unsigned(650, 10), 1200 => to_unsigned(311, 10), 1201 => to_unsigned(864, 10), 1202 => to_unsigned(265, 10), 1203 => to_unsigned(474, 10), 1204 => to_unsigned(605, 10), 1205 => to_unsigned(1007, 10), 1206 => to_unsigned(891, 10), 1207 => to_unsigned(435, 10), 1208 => to_unsigned(20, 10), 1209 => to_unsigned(924, 10), 1210 => to_unsigned(558, 10), 1211 => to_unsigned(887, 10), 1212 => to_unsigned(920, 10), 1213 => to_unsigned(800, 10), 1214 => to_unsigned(907, 10), 1215 => to_unsigned(63, 10), 1216 => to_unsigned(196, 10), 1217 => to_unsigned(523, 10), 1218 => to_unsigned(539, 10), 1219 => to_unsigned(168, 10), 1220 => to_unsigned(781, 10), 1221 => to_unsigned(766, 10), 1222 => to_unsigned(58, 10), 1223 => to_unsigned(128, 10), 1224 => to_unsigned(164, 10), 1225 => to_unsigned(804, 10), 1226 => to_unsigned(75, 10), 1227 => to_unsigned(661, 10), 1228 => to_unsigned(374, 10), 1229 => to_unsigned(460, 10), 1230 => to_unsigned(733, 10), 1231 => to_unsigned(182, 10), 1232 => to_unsigned(750, 10), 1233 => to_unsigned(1014, 10), 1234 => to_unsigned(984, 10), 1235 => to_unsigned(650, 10), 1236 => to_unsigned(663, 10), 1237 => to_unsigned(770, 10), 1238 => to_unsigned(607, 10), 1239 => to_unsigned(358, 10), 1240 => to_unsigned(476, 10), 1241 => to_unsigned(699, 10), 1242 => to_unsigned(804, 10), 1243 => to_unsigned(375, 10), 1244 => to_unsigned(44, 10), 1245 => to_unsigned(812, 10), 1246 => to_unsigned(342, 10), 1247 => to_unsigned(964, 10), 1248 => to_unsigned(328, 10), 1249 => to_unsigned(902, 10), 1250 => to_unsigned(590, 10), 1251 => to_unsigned(148, 10), 1252 => to_unsigned(440, 10), 1253 => to_unsigned(834, 10), 1254 => to_unsigned(595, 10), 1255 => to_unsigned(371, 10), 1256 => to_unsigned(45, 10), 1257 => to_unsigned(580, 10), 1258 => to_unsigned(255, 10), 1259 => to_unsigned(838, 10), 1260 => to_unsigned(696, 10), 1261 => to_unsigned(104, 10), 1262 => to_unsigned(852, 10), 1263 => to_unsigned(568, 10), 1264 => to_unsigned(673, 10), 1265 => to_unsigned(409, 10), 1266 => to_unsigned(640, 10), 1267 => to_unsigned(905, 10), 1268 => to_unsigned(90, 10), 1269 => to_unsigned(981, 10), 1270 => to_unsigned(717, 10), 1271 => to_unsigned(976, 10), 1272 => to_unsigned(409, 10), 1273 => to_unsigned(906, 10), 1274 => to_unsigned(891, 10), 1275 => to_unsigned(955, 10), 1276 => to_unsigned(831, 10), 1277 => to_unsigned(261, 10), 1278 => to_unsigned(138, 10), 1279 => to_unsigned(924, 10), 1280 => to_unsigned(914, 10), 1281 => to_unsigned(107, 10), 1282 => to_unsigned(702, 10), 1283 => to_unsigned(661, 10), 1284 => to_unsigned(826, 10), 1285 => to_unsigned(687, 10), 1286 => to_unsigned(356, 10), 1287 => to_unsigned(591, 10), 1288 => to_unsigned(450, 10), 1289 => to_unsigned(889, 10), 1290 => to_unsigned(457, 10), 1291 => to_unsigned(57, 10), 1292 => to_unsigned(915, 10), 1293 => to_unsigned(104, 10), 1294 => to_unsigned(697, 10), 1295 => to_unsigned(487, 10), 1296 => to_unsigned(306, 10), 1297 => to_unsigned(750, 10), 1298 => to_unsigned(669, 10), 1299 => to_unsigned(775, 10), 1300 => to_unsigned(523, 10), 1301 => to_unsigned(599, 10), 1302 => to_unsigned(374, 10), 1303 => to_unsigned(72, 10), 1304 => to_unsigned(663, 10), 1305 => to_unsigned(836, 10), 1306 => to_unsigned(384, 10), 1307 => to_unsigned(282, 10), 1308 => to_unsigned(501, 10), 1309 => to_unsigned(340, 10), 1310 => to_unsigned(704, 10), 1311 => to_unsigned(337, 10), 1312 => to_unsigned(223, 10), 1313 => to_unsigned(948, 10), 1314 => to_unsigned(709, 10), 1315 => to_unsigned(775, 10), 1316 => to_unsigned(997, 10), 1317 => to_unsigned(503, 10), 1318 => to_unsigned(293, 10), 1319 => to_unsigned(20, 10), 1320 => to_unsigned(620, 10), 1321 => to_unsigned(361, 10), 1322 => to_unsigned(84, 10), 1323 => to_unsigned(158, 10), 1324 => to_unsigned(399, 10), 1325 => to_unsigned(934, 10), 1326 => to_unsigned(156, 10), 1327 => to_unsigned(305, 10), 1328 => to_unsigned(597, 10), 1329 => to_unsigned(494, 10), 1330 => to_unsigned(985, 10), 1331 => to_unsigned(911, 10), 1332 => to_unsigned(432, 10), 1333 => to_unsigned(99, 10), 1334 => to_unsigned(268, 10), 1335 => to_unsigned(632, 10), 1336 => to_unsigned(23, 10), 1337 => to_unsigned(872, 10), 1338 => to_unsigned(677, 10), 1339 => to_unsigned(368, 10), 1340 => to_unsigned(203, 10), 1341 => to_unsigned(465, 10), 1342 => to_unsigned(472, 10), 1343 => to_unsigned(396, 10), 1344 => to_unsigned(503, 10), 1345 => to_unsigned(426, 10), 1346 => to_unsigned(572, 10), 1347 => to_unsigned(411, 10), 1348 => to_unsigned(992, 10), 1349 => to_unsigned(902, 10), 1350 => to_unsigned(826, 10), 1351 => to_unsigned(630, 10), 1352 => to_unsigned(813, 10), 1353 => to_unsigned(620, 10), 1354 => to_unsigned(744, 10), 1355 => to_unsigned(1001, 10), 1356 => to_unsigned(406, 10), 1357 => to_unsigned(140, 10), 1358 => to_unsigned(341, 10), 1359 => to_unsigned(384, 10), 1360 => to_unsigned(874, 10), 1361 => to_unsigned(156, 10), 1362 => to_unsigned(555, 10), 1363 => to_unsigned(739, 10), 1364 => to_unsigned(1008, 10), 1365 => to_unsigned(449, 10), 1366 => to_unsigned(657, 10), 1367 => to_unsigned(375, 10), 1368 => to_unsigned(25, 10), 1369 => to_unsigned(399, 10), 1370 => to_unsigned(717, 10), 1371 => to_unsigned(119, 10), 1372 => to_unsigned(127, 10), 1373 => to_unsigned(277, 10), 1374 => to_unsigned(2, 10), 1375 => to_unsigned(486, 10), 1376 => to_unsigned(654, 10), 1377 => to_unsigned(20, 10), 1378 => to_unsigned(881, 10), 1379 => to_unsigned(535, 10), 1380 => to_unsigned(34, 10), 1381 => to_unsigned(614, 10), 1382 => to_unsigned(246, 10), 1383 => to_unsigned(328, 10), 1384 => to_unsigned(790, 10), 1385 => to_unsigned(7, 10), 1386 => to_unsigned(820, 10), 1387 => to_unsigned(235, 10), 1388 => to_unsigned(831, 10), 1389 => to_unsigned(1, 10), 1390 => to_unsigned(968, 10), 1391 => to_unsigned(412, 10), 1392 => to_unsigned(987, 10), 1393 => to_unsigned(226, 10), 1394 => to_unsigned(157, 10), 1395 => to_unsigned(954, 10), 1396 => to_unsigned(222, 10), 1397 => to_unsigned(905, 10), 1398 => to_unsigned(60, 10), 1399 => to_unsigned(848, 10), 1400 => to_unsigned(1014, 10), 1401 => to_unsigned(631, 10), 1402 => to_unsigned(232, 10), 1403 => to_unsigned(413, 10), 1404 => to_unsigned(176, 10), 1405 => to_unsigned(857, 10), 1406 => to_unsigned(993, 10), 1407 => to_unsigned(321, 10), 1408 => to_unsigned(929, 10), 1409 => to_unsigned(978, 10), 1410 => to_unsigned(284, 10), 1411 => to_unsigned(816, 10), 1412 => to_unsigned(747, 10), 1413 => to_unsigned(616, 10), 1414 => to_unsigned(565, 10), 1415 => to_unsigned(850, 10), 1416 => to_unsigned(326, 10), 1417 => to_unsigned(547, 10), 1418 => to_unsigned(873, 10), 1419 => to_unsigned(393, 10), 1420 => to_unsigned(280, 10), 1421 => to_unsigned(898, 10), 1422 => to_unsigned(27, 10), 1423 => to_unsigned(880, 10), 1424 => to_unsigned(190, 10), 1425 => to_unsigned(578, 10), 1426 => to_unsigned(79, 10), 1427 => to_unsigned(642, 10), 1428 => to_unsigned(587, 10), 1429 => to_unsigned(795, 10), 1430 => to_unsigned(995, 10), 1431 => to_unsigned(111, 10), 1432 => to_unsigned(878, 10), 1433 => to_unsigned(271, 10), 1434 => to_unsigned(36, 10), 1435 => to_unsigned(343, 10), 1436 => to_unsigned(909, 10), 1437 => to_unsigned(306, 10), 1438 => to_unsigned(329, 10), 1439 => to_unsigned(59, 10), 1440 => to_unsigned(636, 10), 1441 => to_unsigned(659, 10), 1442 => to_unsigned(598, 10), 1443 => to_unsigned(758, 10), 1444 => to_unsigned(101, 10), 1445 => to_unsigned(420, 10), 1446 => to_unsigned(828, 10), 1447 => to_unsigned(655, 10), 1448 => to_unsigned(937, 10), 1449 => to_unsigned(187, 10), 1450 => to_unsigned(94, 10), 1451 => to_unsigned(525, 10), 1452 => to_unsigned(1002, 10), 1453 => to_unsigned(580, 10), 1454 => to_unsigned(578, 10), 1455 => to_unsigned(278, 10), 1456 => to_unsigned(470, 10), 1457 => to_unsigned(971, 10), 1458 => to_unsigned(892, 10), 1459 => to_unsigned(598, 10), 1460 => to_unsigned(605, 10), 1461 => to_unsigned(420, 10), 1462 => to_unsigned(98, 10), 1463 => to_unsigned(480, 10), 1464 => to_unsigned(608, 10), 1465 => to_unsigned(920, 10), 1466 => to_unsigned(824, 10), 1467 => to_unsigned(922, 10), 1468 => to_unsigned(279, 10), 1469 => to_unsigned(104, 10), 1470 => to_unsigned(374, 10), 1471 => to_unsigned(756, 10), 1472 => to_unsigned(722, 10), 1473 => to_unsigned(835, 10), 1474 => to_unsigned(984, 10), 1475 => to_unsigned(338, 10), 1476 => to_unsigned(629, 10), 1477 => to_unsigned(25, 10), 1478 => to_unsigned(799, 10), 1479 => to_unsigned(440, 10), 1480 => to_unsigned(553, 10), 1481 => to_unsigned(268, 10), 1482 => to_unsigned(562, 10), 1483 => to_unsigned(799, 10), 1484 => to_unsigned(160, 10), 1485 => to_unsigned(47, 10), 1486 => to_unsigned(264, 10), 1487 => to_unsigned(903, 10), 1488 => to_unsigned(105, 10), 1489 => to_unsigned(373, 10), 1490 => to_unsigned(666, 10), 1491 => to_unsigned(590, 10), 1492 => to_unsigned(222, 10), 1493 => to_unsigned(40, 10), 1494 => to_unsigned(686, 10), 1495 => to_unsigned(650, 10), 1496 => to_unsigned(843, 10), 1497 => to_unsigned(126, 10), 1498 => to_unsigned(968, 10), 1499 => to_unsigned(943, 10), 1500 => to_unsigned(401, 10), 1501 => to_unsigned(545, 10), 1502 => to_unsigned(35, 10), 1503 => to_unsigned(638, 10), 1504 => to_unsigned(928, 10), 1505 => to_unsigned(755, 10), 1506 => to_unsigned(945, 10), 1507 => to_unsigned(906, 10), 1508 => to_unsigned(846, 10), 1509 => to_unsigned(644, 10), 1510 => to_unsigned(630, 10), 1511 => to_unsigned(960, 10), 1512 => to_unsigned(805, 10), 1513 => to_unsigned(290, 10), 1514 => to_unsigned(53, 10), 1515 => to_unsigned(596, 10), 1516 => to_unsigned(965, 10), 1517 => to_unsigned(638, 10), 1518 => to_unsigned(399, 10), 1519 => to_unsigned(525, 10), 1520 => to_unsigned(710, 10), 1521 => to_unsigned(620, 10), 1522 => to_unsigned(495, 10), 1523 => to_unsigned(302, 10), 1524 => to_unsigned(114, 10), 1525 => to_unsigned(764, 10), 1526 => to_unsigned(195, 10), 1527 => to_unsigned(488, 10), 1528 => to_unsigned(245, 10), 1529 => to_unsigned(172, 10), 1530 => to_unsigned(51, 10), 1531 => to_unsigned(781, 10), 1532 => to_unsigned(781, 10), 1533 => to_unsigned(391, 10), 1534 => to_unsigned(474, 10), 1535 => to_unsigned(690, 10), 1536 => to_unsigned(864, 10), 1537 => to_unsigned(870, 10), 1538 => to_unsigned(794, 10), 1539 => to_unsigned(332, 10), 1540 => to_unsigned(815, 10), 1541 => to_unsigned(111, 10), 1542 => to_unsigned(241, 10), 1543 => to_unsigned(701, 10), 1544 => to_unsigned(407, 10), 1545 => to_unsigned(2, 10), 1546 => to_unsigned(435, 10), 1547 => to_unsigned(979, 10), 1548 => to_unsigned(211, 10), 1549 => to_unsigned(731, 10), 1550 => to_unsigned(137, 10), 1551 => to_unsigned(420, 10), 1552 => to_unsigned(978, 10), 1553 => to_unsigned(288, 10), 1554 => to_unsigned(913, 10), 1555 => to_unsigned(389, 10), 1556 => to_unsigned(670, 10), 1557 => to_unsigned(158, 10), 1558 => to_unsigned(1017, 10), 1559 => to_unsigned(821, 10), 1560 => to_unsigned(769, 10), 1561 => to_unsigned(122, 10), 1562 => to_unsigned(444, 10), 1563 => to_unsigned(73, 10), 1564 => to_unsigned(482, 10), 1565 => to_unsigned(652, 10), 1566 => to_unsigned(697, 10), 1567 => to_unsigned(694, 10), 1568 => to_unsigned(638, 10), 1569 => to_unsigned(200, 10), 1570 => to_unsigned(38, 10), 1571 => to_unsigned(55, 10), 1572 => to_unsigned(574, 10), 1573 => to_unsigned(986, 10), 1574 => to_unsigned(316, 10), 1575 => to_unsigned(395, 10), 1576 => to_unsigned(1011, 10), 1577 => to_unsigned(817, 10), 1578 => to_unsigned(893, 10), 1579 => to_unsigned(452, 10), 1580 => to_unsigned(133, 10), 1581 => to_unsigned(301, 10), 1582 => to_unsigned(289, 10), 1583 => to_unsigned(756, 10), 1584 => to_unsigned(856, 10), 1585 => to_unsigned(972, 10), 1586 => to_unsigned(861, 10), 1587 => to_unsigned(192, 10), 1588 => to_unsigned(219, 10), 1589 => to_unsigned(69, 10), 1590 => to_unsigned(1000, 10), 1591 => to_unsigned(429, 10), 1592 => to_unsigned(850, 10), 1593 => to_unsigned(690, 10), 1594 => to_unsigned(34, 10), 1595 => to_unsigned(506, 10), 1596 => to_unsigned(63, 10), 1597 => to_unsigned(529, 10), 1598 => to_unsigned(909, 10), 1599 => to_unsigned(85, 10), 1600 => to_unsigned(485, 10), 1601 => to_unsigned(970, 10), 1602 => to_unsigned(579, 10), 1603 => to_unsigned(913, 10), 1604 => to_unsigned(122, 10), 1605 => to_unsigned(178, 10), 1606 => to_unsigned(227, 10), 1607 => to_unsigned(588, 10), 1608 => to_unsigned(367, 10), 1609 => to_unsigned(176, 10), 1610 => to_unsigned(450, 10), 1611 => to_unsigned(657, 10), 1612 => to_unsigned(540, 10), 1613 => to_unsigned(272, 10), 1614 => to_unsigned(4, 10), 1615 => to_unsigned(32, 10), 1616 => to_unsigned(689, 10), 1617 => to_unsigned(81, 10), 1618 => to_unsigned(967, 10), 1619 => to_unsigned(18, 10), 1620 => to_unsigned(312, 10), 1621 => to_unsigned(70, 10), 1622 => to_unsigned(962, 10), 1623 => to_unsigned(568, 10), 1624 => to_unsigned(466, 10), 1625 => to_unsigned(870, 10), 1626 => to_unsigned(824, 10), 1627 => to_unsigned(656, 10), 1628 => to_unsigned(742, 10), 1629 => to_unsigned(151, 10), 1630 => to_unsigned(793, 10), 1631 => to_unsigned(822, 10), 1632 => to_unsigned(556, 10), 1633 => to_unsigned(884, 10), 1634 => to_unsigned(87, 10), 1635 => to_unsigned(339, 10), 1636 => to_unsigned(684, 10), 1637 => to_unsigned(927, 10), 1638 => to_unsigned(94, 10), 1639 => to_unsigned(961, 10), 1640 => to_unsigned(97, 10), 1641 => to_unsigned(24, 10), 1642 => to_unsigned(982, 10), 1643 => to_unsigned(929, 10), 1644 => to_unsigned(723, 10), 1645 => to_unsigned(926, 10), 1646 => to_unsigned(1021, 10), 1647 => to_unsigned(602, 10), 1648 => to_unsigned(546, 10), 1649 => to_unsigned(980, 10), 1650 => to_unsigned(1008, 10), 1651 => to_unsigned(740, 10), 1652 => to_unsigned(81, 10), 1653 => to_unsigned(528, 10), 1654 => to_unsigned(303, 10), 1655 => to_unsigned(826, 10), 1656 => to_unsigned(731, 10), 1657 => to_unsigned(857, 10), 1658 => to_unsigned(674, 10), 1659 => to_unsigned(227, 10), 1660 => to_unsigned(507, 10), 1661 => to_unsigned(870, 10), 1662 => to_unsigned(390, 10), 1663 => to_unsigned(30, 10), 1664 => to_unsigned(824, 10), 1665 => to_unsigned(849, 10), 1666 => to_unsigned(845, 10), 1667 => to_unsigned(304, 10), 1668 => to_unsigned(948, 10), 1669 => to_unsigned(493, 10), 1670 => to_unsigned(379, 10), 1671 => to_unsigned(629, 10), 1672 => to_unsigned(130, 10), 1673 => to_unsigned(26, 10), 1674 => to_unsigned(636, 10), 1675 => to_unsigned(951, 10), 1676 => to_unsigned(152, 10), 1677 => to_unsigned(1007, 10), 1678 => to_unsigned(284, 10), 1679 => to_unsigned(968, 10), 1680 => to_unsigned(503, 10), 1681 => to_unsigned(228, 10), 1682 => to_unsigned(204, 10), 1683 => to_unsigned(37, 10), 1684 => to_unsigned(895, 10), 1685 => to_unsigned(1001, 10), 1686 => to_unsigned(965, 10), 1687 => to_unsigned(129, 10), 1688 => to_unsigned(233, 10), 1689 => to_unsigned(808, 10), 1690 => to_unsigned(338, 10), 1691 => to_unsigned(248, 10), 1692 => to_unsigned(170, 10), 1693 => to_unsigned(341, 10), 1694 => to_unsigned(64, 10), 1695 => to_unsigned(336, 10), 1696 => to_unsigned(681, 10), 1697 => to_unsigned(236, 10), 1698 => to_unsigned(39, 10), 1699 => to_unsigned(223, 10), 1700 => to_unsigned(613, 10), 1701 => to_unsigned(108, 10), 1702 => to_unsigned(472, 10), 1703 => to_unsigned(115, 10), 1704 => to_unsigned(539, 10), 1705 => to_unsigned(869, 10), 1706 => to_unsigned(589, 10), 1707 => to_unsigned(668, 10), 1708 => to_unsigned(58, 10), 1709 => to_unsigned(993, 10), 1710 => to_unsigned(961, 10), 1711 => to_unsigned(534, 10), 1712 => to_unsigned(77, 10), 1713 => to_unsigned(270, 10), 1714 => to_unsigned(996, 10), 1715 => to_unsigned(89, 10), 1716 => to_unsigned(416, 10), 1717 => to_unsigned(198, 10), 1718 => to_unsigned(273, 10), 1719 => to_unsigned(39, 10), 1720 => to_unsigned(4, 10), 1721 => to_unsigned(628, 10), 1722 => to_unsigned(154, 10), 1723 => to_unsigned(94, 10), 1724 => to_unsigned(136, 10), 1725 => to_unsigned(142, 10), 1726 => to_unsigned(184, 10), 1727 => to_unsigned(90, 10), 1728 => to_unsigned(785, 10), 1729 => to_unsigned(980, 10), 1730 => to_unsigned(28, 10), 1731 => to_unsigned(811, 10), 1732 => to_unsigned(259, 10), 1733 => to_unsigned(448, 10), 1734 => to_unsigned(12, 10), 1735 => to_unsigned(595, 10), 1736 => to_unsigned(62, 10), 1737 => to_unsigned(638, 10), 1738 => to_unsigned(567, 10), 1739 => to_unsigned(703, 10), 1740 => to_unsigned(442, 10), 1741 => to_unsigned(340, 10), 1742 => to_unsigned(521, 10), 1743 => to_unsigned(936, 10), 1744 => to_unsigned(817, 10), 1745 => to_unsigned(195, 10), 1746 => to_unsigned(607, 10), 1747 => to_unsigned(269, 10), 1748 => to_unsigned(108, 10), 1749 => to_unsigned(343, 10), 1750 => to_unsigned(274, 10), 1751 => to_unsigned(255, 10), 1752 => to_unsigned(572, 10), 1753 => to_unsigned(327, 10), 1754 => to_unsigned(684, 10), 1755 => to_unsigned(432, 10), 1756 => to_unsigned(811, 10), 1757 => to_unsigned(982, 10), 1758 => to_unsigned(489, 10), 1759 => to_unsigned(695, 10), 1760 => to_unsigned(683, 10), 1761 => to_unsigned(52, 10), 1762 => to_unsigned(181, 10), 1763 => to_unsigned(406, 10), 1764 => to_unsigned(322, 10), 1765 => to_unsigned(1006, 10), 1766 => to_unsigned(566, 10), 1767 => to_unsigned(965, 10), 1768 => to_unsigned(591, 10), 1769 => to_unsigned(1023, 10), 1770 => to_unsigned(903, 10), 1771 => to_unsigned(889, 10), 1772 => to_unsigned(225, 10), 1773 => to_unsigned(986, 10), 1774 => to_unsigned(918, 10), 1775 => to_unsigned(674, 10), 1776 => to_unsigned(220, 10), 1777 => to_unsigned(260, 10), 1778 => to_unsigned(1001, 10), 1779 => to_unsigned(999, 10), 1780 => to_unsigned(439, 10), 1781 => to_unsigned(73, 10), 1782 => to_unsigned(80, 10), 1783 => to_unsigned(956, 10), 1784 => to_unsigned(282, 10), 1785 => to_unsigned(805, 10), 1786 => to_unsigned(894, 10), 1787 => to_unsigned(45, 10), 1788 => to_unsigned(890, 10), 1789 => to_unsigned(486, 10), 1790 => to_unsigned(324, 10), 1791 => to_unsigned(395, 10), 1792 => to_unsigned(701, 10), 1793 => to_unsigned(402, 10), 1794 => to_unsigned(992, 10), 1795 => to_unsigned(215, 10), 1796 => to_unsigned(400, 10), 1797 => to_unsigned(127, 10), 1798 => to_unsigned(141, 10), 1799 => to_unsigned(259, 10), 1800 => to_unsigned(240, 10), 1801 => to_unsigned(396, 10), 1802 => to_unsigned(123, 10), 1803 => to_unsigned(945, 10), 1804 => to_unsigned(839, 10), 1805 => to_unsigned(860, 10), 1806 => to_unsigned(282, 10), 1807 => to_unsigned(620, 10), 1808 => to_unsigned(91, 10), 1809 => to_unsigned(392, 10), 1810 => to_unsigned(869, 10), 1811 => to_unsigned(157, 10), 1812 => to_unsigned(613, 10), 1813 => to_unsigned(229, 10), 1814 => to_unsigned(441, 10), 1815 => to_unsigned(699, 10), 1816 => to_unsigned(48, 10), 1817 => to_unsigned(143, 10), 1818 => to_unsigned(1017, 10), 1819 => to_unsigned(737, 10), 1820 => to_unsigned(518, 10), 1821 => to_unsigned(199, 10), 1822 => to_unsigned(455, 10), 1823 => to_unsigned(164, 10), 1824 => to_unsigned(148, 10), 1825 => to_unsigned(424, 10), 1826 => to_unsigned(176, 10), 1827 => to_unsigned(235, 10), 1828 => to_unsigned(84, 10), 1829 => to_unsigned(417, 10), 1830 => to_unsigned(675, 10), 1831 => to_unsigned(214, 10), 1832 => to_unsigned(570, 10), 1833 => to_unsigned(909, 10), 1834 => to_unsigned(942, 10), 1835 => to_unsigned(451, 10), 1836 => to_unsigned(370, 10), 1837 => to_unsigned(842, 10), 1838 => to_unsigned(32, 10), 1839 => to_unsigned(896, 10), 1840 => to_unsigned(264, 10), 1841 => to_unsigned(62, 10), 1842 => to_unsigned(419, 10), 1843 => to_unsigned(706, 10), 1844 => to_unsigned(10, 10), 1845 => to_unsigned(176, 10), 1846 => to_unsigned(287, 10), 1847 => to_unsigned(941, 10), 1848 => to_unsigned(979, 10), 1849 => to_unsigned(446, 10), 1850 => to_unsigned(501, 10), 1851 => to_unsigned(339, 10), 1852 => to_unsigned(867, 10), 1853 => to_unsigned(646, 10), 1854 => to_unsigned(440, 10), 1855 => to_unsigned(467, 10), 1856 => to_unsigned(315, 10), 1857 => to_unsigned(230, 10), 1858 => to_unsigned(502, 10), 1859 => to_unsigned(956, 10), 1860 => to_unsigned(849, 10), 1861 => to_unsigned(318, 10), 1862 => to_unsigned(282, 10), 1863 => to_unsigned(250, 10), 1864 => to_unsigned(770, 10), 1865 => to_unsigned(875, 10), 1866 => to_unsigned(344, 10), 1867 => to_unsigned(473, 10), 1868 => to_unsigned(808, 10), 1869 => to_unsigned(499, 10), 1870 => to_unsigned(113, 10), 1871 => to_unsigned(340, 10), 1872 => to_unsigned(970, 10), 1873 => to_unsigned(691, 10), 1874 => to_unsigned(914, 10), 1875 => to_unsigned(189, 10), 1876 => to_unsigned(741, 10), 1877 => to_unsigned(839, 10), 1878 => to_unsigned(236, 10), 1879 => to_unsigned(516, 10), 1880 => to_unsigned(161, 10), 1881 => to_unsigned(903, 10), 1882 => to_unsigned(553, 10), 1883 => to_unsigned(770, 10), 1884 => to_unsigned(446, 10), 1885 => to_unsigned(938, 10), 1886 => to_unsigned(760, 10), 1887 => to_unsigned(924, 10), 1888 => to_unsigned(537, 10), 1889 => to_unsigned(56, 10), 1890 => to_unsigned(25, 10), 1891 => to_unsigned(982, 10), 1892 => to_unsigned(433, 10), 1893 => to_unsigned(181, 10), 1894 => to_unsigned(221, 10), 1895 => to_unsigned(958, 10), 1896 => to_unsigned(218, 10), 1897 => to_unsigned(958, 10), 1898 => to_unsigned(829, 10), 1899 => to_unsigned(371, 10), 1900 => to_unsigned(829, 10), 1901 => to_unsigned(638, 10), 1902 => to_unsigned(120, 10), 1903 => to_unsigned(600, 10), 1904 => to_unsigned(123, 10), 1905 => to_unsigned(275, 10), 1906 => to_unsigned(736, 10), 1907 => to_unsigned(809, 10), 1908 => to_unsigned(880, 10), 1909 => to_unsigned(1008, 10), 1910 => to_unsigned(535, 10), 1911 => to_unsigned(53, 10), 1912 => to_unsigned(524, 10), 1913 => to_unsigned(736, 10), 1914 => to_unsigned(78, 10), 1915 => to_unsigned(937, 10), 1916 => to_unsigned(305, 10), 1917 => to_unsigned(540, 10), 1918 => to_unsigned(952, 10), 1919 => to_unsigned(551, 10), 1920 => to_unsigned(473, 10), 1921 => to_unsigned(73, 10), 1922 => to_unsigned(460, 10), 1923 => to_unsigned(753, 10), 1924 => to_unsigned(269, 10), 1925 => to_unsigned(1016, 10), 1926 => to_unsigned(805, 10), 1927 => to_unsigned(475, 10), 1928 => to_unsigned(840, 10), 1929 => to_unsigned(553, 10), 1930 => to_unsigned(574, 10), 1931 => to_unsigned(808, 10), 1932 => to_unsigned(545, 10), 1933 => to_unsigned(765, 10), 1934 => to_unsigned(0, 10), 1935 => to_unsigned(15, 10), 1936 => to_unsigned(294, 10), 1937 => to_unsigned(419, 10), 1938 => to_unsigned(275, 10), 1939 => to_unsigned(484, 10), 1940 => to_unsigned(806, 10), 1941 => to_unsigned(865, 10), 1942 => to_unsigned(103, 10), 1943 => to_unsigned(461, 10), 1944 => to_unsigned(548, 10), 1945 => to_unsigned(619, 10), 1946 => to_unsigned(320, 10), 1947 => to_unsigned(168, 10), 1948 => to_unsigned(394, 10), 1949 => to_unsigned(295, 10), 1950 => to_unsigned(232, 10), 1951 => to_unsigned(274, 10), 1952 => to_unsigned(366, 10), 1953 => to_unsigned(940, 10), 1954 => to_unsigned(422, 10), 1955 => to_unsigned(3, 10), 1956 => to_unsigned(739, 10), 1957 => to_unsigned(997, 10), 1958 => to_unsigned(253, 10), 1959 => to_unsigned(754, 10), 1960 => to_unsigned(767, 10), 1961 => to_unsigned(334, 10), 1962 => to_unsigned(978, 10), 1963 => to_unsigned(593, 10), 1964 => to_unsigned(245, 10), 1965 => to_unsigned(133, 10), 1966 => to_unsigned(73, 10), 1967 => to_unsigned(819, 10), 1968 => to_unsigned(591, 10), 1969 => to_unsigned(458, 10), 1970 => to_unsigned(934, 10), 1971 => to_unsigned(884, 10), 1972 => to_unsigned(158, 10), 1973 => to_unsigned(645, 10), 1974 => to_unsigned(203, 10), 1975 => to_unsigned(278, 10), 1976 => to_unsigned(489, 10), 1977 => to_unsigned(892, 10), 1978 => to_unsigned(599, 10), 1979 => to_unsigned(921, 10), 1980 => to_unsigned(789, 10), 1981 => to_unsigned(71, 10), 1982 => to_unsigned(945, 10), 1983 => to_unsigned(529, 10), 1984 => to_unsigned(862, 10), 1985 => to_unsigned(714, 10), 1986 => to_unsigned(897, 10), 1987 => to_unsigned(329, 10), 1988 => to_unsigned(367, 10), 1989 => to_unsigned(648, 10), 1990 => to_unsigned(901, 10), 1991 => to_unsigned(970, 10), 1992 => to_unsigned(996, 10), 1993 => to_unsigned(605, 10), 1994 => to_unsigned(430, 10), 1995 => to_unsigned(440, 10), 1996 => to_unsigned(699, 10), 1997 => to_unsigned(369, 10), 1998 => to_unsigned(288, 10), 1999 => to_unsigned(225, 10), 2000 => to_unsigned(511, 10), 2001 => to_unsigned(653, 10), 2002 => to_unsigned(277, 10), 2003 => to_unsigned(890, 10), 2004 => to_unsigned(538, 10), 2005 => to_unsigned(636, 10), 2006 => to_unsigned(904, 10), 2007 => to_unsigned(925, 10), 2008 => to_unsigned(748, 10), 2009 => to_unsigned(698, 10), 2010 => to_unsigned(962, 10), 2011 => to_unsigned(279, 10), 2012 => to_unsigned(258, 10), 2013 => to_unsigned(725, 10), 2014 => to_unsigned(827, 10), 2015 => to_unsigned(731, 10), 2016 => to_unsigned(537, 10), 2017 => to_unsigned(192, 10), 2018 => to_unsigned(403, 10), 2019 => to_unsigned(131, 10), 2020 => to_unsigned(628, 10), 2021 => to_unsigned(941, 10), 2022 => to_unsigned(483, 10), 2023 => to_unsigned(1015, 10), 2024 => to_unsigned(962, 10), 2025 => to_unsigned(707, 10), 2026 => to_unsigned(229, 10), 2027 => to_unsigned(449, 10), 2028 => to_unsigned(243, 10), 2029 => to_unsigned(585, 10), 2030 => to_unsigned(96, 10), 2031 => to_unsigned(230, 10), 2032 => to_unsigned(181, 10), 2033 => to_unsigned(602, 10), 2034 => to_unsigned(620, 10), 2035 => to_unsigned(515, 10), 2036 => to_unsigned(615, 10), 2037 => to_unsigned(319, 10), 2038 => to_unsigned(543, 10), 2039 => to_unsigned(166, 10), 2040 => to_unsigned(124, 10), 2041 => to_unsigned(510, 10), 2042 => to_unsigned(100, 10), 2043 => to_unsigned(284, 10), 2044 => to_unsigned(772, 10), 2045 => to_unsigned(178, 10), 2046 => to_unsigned(319, 10), 2047 => to_unsigned(393, 10)),
            1 => (0 => to_unsigned(168, 10), 1 => to_unsigned(784, 10), 2 => to_unsigned(974, 10), 3 => to_unsigned(744, 10), 4 => to_unsigned(474, 10), 5 => to_unsigned(735, 10), 6 => to_unsigned(851, 10), 7 => to_unsigned(430, 10), 8 => to_unsigned(596, 10), 9 => to_unsigned(971, 10), 10 => to_unsigned(689, 10), 11 => to_unsigned(906, 10), 12 => to_unsigned(880, 10), 13 => to_unsigned(405, 10), 14 => to_unsigned(711, 10), 15 => to_unsigned(501, 10), 16 => to_unsigned(940, 10), 17 => to_unsigned(886, 10), 18 => to_unsigned(768, 10), 19 => to_unsigned(882, 10), 20 => to_unsigned(462, 10), 21 => to_unsigned(45, 10), 22 => to_unsigned(203, 10), 23 => to_unsigned(560, 10), 24 => to_unsigned(584, 10), 25 => to_unsigned(823, 10), 26 => to_unsigned(239, 10), 27 => to_unsigned(1015, 10), 28 => to_unsigned(412, 10), 29 => to_unsigned(974, 10), 30 => to_unsigned(742, 10), 31 => to_unsigned(599, 10), 32 => to_unsigned(307, 10), 33 => to_unsigned(706, 10), 34 => to_unsigned(1007, 10), 35 => to_unsigned(438, 10), 36 => to_unsigned(933, 10), 37 => to_unsigned(699, 10), 38 => to_unsigned(827, 10), 39 => to_unsigned(743, 10), 40 => to_unsigned(614, 10), 41 => to_unsigned(184, 10), 42 => to_unsigned(315, 10), 43 => to_unsigned(396, 10), 44 => to_unsigned(816, 10), 45 => to_unsigned(807, 10), 46 => to_unsigned(774, 10), 47 => to_unsigned(780, 10), 48 => to_unsigned(422, 10), 49 => to_unsigned(524, 10), 50 => to_unsigned(131, 10), 51 => to_unsigned(336, 10), 52 => to_unsigned(728, 10), 53 => to_unsigned(288, 10), 54 => to_unsigned(296, 10), 55 => to_unsigned(643, 10), 56 => to_unsigned(143, 10), 57 => to_unsigned(740, 10), 58 => to_unsigned(911, 10), 59 => to_unsigned(199, 10), 60 => to_unsigned(327, 10), 61 => to_unsigned(313, 10), 62 => to_unsigned(247, 10), 63 => to_unsigned(282, 10), 64 => to_unsigned(262, 10), 65 => to_unsigned(554, 10), 66 => to_unsigned(372, 10), 67 => to_unsigned(510, 10), 68 => to_unsigned(858, 10), 69 => to_unsigned(943, 10), 70 => to_unsigned(50, 10), 71 => to_unsigned(788, 10), 72 => to_unsigned(702, 10), 73 => to_unsigned(604, 10), 74 => to_unsigned(210, 10), 75 => to_unsigned(383, 10), 76 => to_unsigned(799, 10), 77 => to_unsigned(140, 10), 78 => to_unsigned(220, 10), 79 => to_unsigned(710, 10), 80 => to_unsigned(158, 10), 81 => to_unsigned(232, 10), 82 => to_unsigned(373, 10), 83 => to_unsigned(820, 10), 84 => to_unsigned(585, 10), 85 => to_unsigned(938, 10), 86 => to_unsigned(525, 10), 87 => to_unsigned(366, 10), 88 => to_unsigned(97, 10), 89 => to_unsigned(241, 10), 90 => to_unsigned(642, 10), 91 => to_unsigned(190, 10), 92 => to_unsigned(684, 10), 93 => to_unsigned(112, 10), 94 => to_unsigned(532, 10), 95 => to_unsigned(218, 10), 96 => to_unsigned(925, 10), 97 => to_unsigned(355, 10), 98 => to_unsigned(727, 10), 99 => to_unsigned(717, 10), 100 => to_unsigned(445, 10), 101 => to_unsigned(639, 10), 102 => to_unsigned(191, 10), 103 => to_unsigned(67, 10), 104 => to_unsigned(986, 10), 105 => to_unsigned(870, 10), 106 => to_unsigned(803, 10), 107 => to_unsigned(735, 10), 108 => to_unsigned(1003, 10), 109 => to_unsigned(861, 10), 110 => to_unsigned(471, 10), 111 => to_unsigned(987, 10), 112 => to_unsigned(975, 10), 113 => to_unsigned(398, 10), 114 => to_unsigned(251, 10), 115 => to_unsigned(643, 10), 116 => to_unsigned(716, 10), 117 => to_unsigned(565, 10), 118 => to_unsigned(724, 10), 119 => to_unsigned(553, 10), 120 => to_unsigned(299, 10), 121 => to_unsigned(767, 10), 122 => to_unsigned(756, 10), 123 => to_unsigned(78, 10), 124 => to_unsigned(268, 10), 125 => to_unsigned(978, 10), 126 => to_unsigned(1011, 10), 127 => to_unsigned(74, 10), 128 => to_unsigned(822, 10), 129 => to_unsigned(903, 10), 130 => to_unsigned(718, 10), 131 => to_unsigned(839, 10), 132 => to_unsigned(342, 10), 133 => to_unsigned(859, 10), 134 => to_unsigned(107, 10), 135 => to_unsigned(774, 10), 136 => to_unsigned(491, 10), 137 => to_unsigned(241, 10), 138 => to_unsigned(470, 10), 139 => to_unsigned(110, 10), 140 => to_unsigned(281, 10), 141 => to_unsigned(629, 10), 142 => to_unsigned(112, 10), 143 => to_unsigned(890, 10), 144 => to_unsigned(566, 10), 145 => to_unsigned(714, 10), 146 => to_unsigned(629, 10), 147 => to_unsigned(610, 10), 148 => to_unsigned(461, 10), 149 => to_unsigned(191, 10), 150 => to_unsigned(1006, 10), 151 => to_unsigned(205, 10), 152 => to_unsigned(925, 10), 153 => to_unsigned(7, 10), 154 => to_unsigned(682, 10), 155 => to_unsigned(448, 10), 156 => to_unsigned(886, 10), 157 => to_unsigned(700, 10), 158 => to_unsigned(616, 10), 159 => to_unsigned(818, 10), 160 => to_unsigned(1023, 10), 161 => to_unsigned(734, 10), 162 => to_unsigned(187, 10), 163 => to_unsigned(301, 10), 164 => to_unsigned(885, 10), 165 => to_unsigned(1014, 10), 166 => to_unsigned(882, 10), 167 => to_unsigned(308, 10), 168 => to_unsigned(476, 10), 169 => to_unsigned(275, 10), 170 => to_unsigned(489, 10), 171 => to_unsigned(594, 10), 172 => to_unsigned(807, 10), 173 => to_unsigned(147, 10), 174 => to_unsigned(4, 10), 175 => to_unsigned(1016, 10), 176 => to_unsigned(287, 10), 177 => to_unsigned(660, 10), 178 => to_unsigned(872, 10), 179 => to_unsigned(170, 10), 180 => to_unsigned(72, 10), 181 => to_unsigned(266, 10), 182 => to_unsigned(170, 10), 183 => to_unsigned(812, 10), 184 => to_unsigned(632, 10), 185 => to_unsigned(895, 10), 186 => to_unsigned(149, 10), 187 => to_unsigned(247, 10), 188 => to_unsigned(392, 10), 189 => to_unsigned(567, 10), 190 => to_unsigned(35, 10), 191 => to_unsigned(367, 10), 192 => to_unsigned(351, 10), 193 => to_unsigned(451, 10), 194 => to_unsigned(9, 10), 195 => to_unsigned(557, 10), 196 => to_unsigned(46, 10), 197 => to_unsigned(764, 10), 198 => to_unsigned(816, 10), 199 => to_unsigned(277, 10), 200 => to_unsigned(986, 10), 201 => to_unsigned(585, 10), 202 => to_unsigned(551, 10), 203 => to_unsigned(943, 10), 204 => to_unsigned(884, 10), 205 => to_unsigned(901, 10), 206 => to_unsigned(590, 10), 207 => to_unsigned(272, 10), 208 => to_unsigned(147, 10), 209 => to_unsigned(49, 10), 210 => to_unsigned(322, 10), 211 => to_unsigned(16, 10), 212 => to_unsigned(565, 10), 213 => to_unsigned(1014, 10), 214 => to_unsigned(1002, 10), 215 => to_unsigned(362, 10), 216 => to_unsigned(386, 10), 217 => to_unsigned(905, 10), 218 => to_unsigned(807, 10), 219 => to_unsigned(583, 10), 220 => to_unsigned(304, 10), 221 => to_unsigned(736, 10), 222 => to_unsigned(343, 10), 223 => to_unsigned(688, 10), 224 => to_unsigned(807, 10), 225 => to_unsigned(880, 10), 226 => to_unsigned(507, 10), 227 => to_unsigned(123, 10), 228 => to_unsigned(937, 10), 229 => to_unsigned(524, 10), 230 => to_unsigned(588, 10), 231 => to_unsigned(751, 10), 232 => to_unsigned(611, 10), 233 => to_unsigned(460, 10), 234 => to_unsigned(616, 10), 235 => to_unsigned(383, 10), 236 => to_unsigned(893, 10), 237 => to_unsigned(584, 10), 238 => to_unsigned(801, 10), 239 => to_unsigned(797, 10), 240 => to_unsigned(48, 10), 241 => to_unsigned(288, 10), 242 => to_unsigned(121, 10), 243 => to_unsigned(202, 10), 244 => to_unsigned(752, 10), 245 => to_unsigned(344, 10), 246 => to_unsigned(693, 10), 247 => to_unsigned(477, 10), 248 => to_unsigned(192, 10), 249 => to_unsigned(196, 10), 250 => to_unsigned(599, 10), 251 => to_unsigned(16, 10), 252 => to_unsigned(208, 10), 253 => to_unsigned(197, 10), 254 => to_unsigned(428, 10), 255 => to_unsigned(194, 10), 256 => to_unsigned(617, 10), 257 => to_unsigned(824, 10), 258 => to_unsigned(783, 10), 259 => to_unsigned(691, 10), 260 => to_unsigned(884, 10), 261 => to_unsigned(475, 10), 262 => to_unsigned(644, 10), 263 => to_unsigned(889, 10), 264 => to_unsigned(868, 10), 265 => to_unsigned(302, 10), 266 => to_unsigned(733, 10), 267 => to_unsigned(338, 10), 268 => to_unsigned(419, 10), 269 => to_unsigned(93, 10), 270 => to_unsigned(375, 10), 271 => to_unsigned(869, 10), 272 => to_unsigned(473, 10), 273 => to_unsigned(16, 10), 274 => to_unsigned(487, 10), 275 => to_unsigned(714, 10), 276 => to_unsigned(535, 10), 277 => to_unsigned(451, 10), 278 => to_unsigned(644, 10), 279 => to_unsigned(557, 10), 280 => to_unsigned(135, 10), 281 => to_unsigned(311, 10), 282 => to_unsigned(218, 10), 283 => to_unsigned(896, 10), 284 => to_unsigned(723, 10), 285 => to_unsigned(156, 10), 286 => to_unsigned(95, 10), 287 => to_unsigned(754, 10), 288 => to_unsigned(954, 10), 289 => to_unsigned(70, 10), 290 => to_unsigned(871, 10), 291 => to_unsigned(485, 10), 292 => to_unsigned(0, 10), 293 => to_unsigned(95, 10), 294 => to_unsigned(149, 10), 295 => to_unsigned(688, 10), 296 => to_unsigned(207, 10), 297 => to_unsigned(575, 10), 298 => to_unsigned(107, 10), 299 => to_unsigned(270, 10), 300 => to_unsigned(149, 10), 301 => to_unsigned(508, 10), 302 => to_unsigned(573, 10), 303 => to_unsigned(110, 10), 304 => to_unsigned(599, 10), 305 => to_unsigned(855, 10), 306 => to_unsigned(369, 10), 307 => to_unsigned(447, 10), 308 => to_unsigned(651, 10), 309 => to_unsigned(39, 10), 310 => to_unsigned(132, 10), 311 => to_unsigned(928, 10), 312 => to_unsigned(876, 10), 313 => to_unsigned(187, 10), 314 => to_unsigned(114, 10), 315 => to_unsigned(494, 10), 316 => to_unsigned(449, 10), 317 => to_unsigned(575, 10), 318 => to_unsigned(921, 10), 319 => to_unsigned(810, 10), 320 => to_unsigned(83, 10), 321 => to_unsigned(847, 10), 322 => to_unsigned(393, 10), 323 => to_unsigned(232, 10), 324 => to_unsigned(78, 10), 325 => to_unsigned(458, 10), 326 => to_unsigned(276, 10), 327 => to_unsigned(457, 10), 328 => to_unsigned(645, 10), 329 => to_unsigned(467, 10), 330 => to_unsigned(520, 10), 331 => to_unsigned(527, 10), 332 => to_unsigned(698, 10), 333 => to_unsigned(79, 10), 334 => to_unsigned(980, 10), 335 => to_unsigned(138, 10), 336 => to_unsigned(294, 10), 337 => to_unsigned(106, 10), 338 => to_unsigned(1023, 10), 339 => to_unsigned(586, 10), 340 => to_unsigned(191, 10), 341 => to_unsigned(359, 10), 342 => to_unsigned(139, 10), 343 => to_unsigned(117, 10), 344 => to_unsigned(931, 10), 345 => to_unsigned(802, 10), 346 => to_unsigned(753, 10), 347 => to_unsigned(207, 10), 348 => to_unsigned(683, 10), 349 => to_unsigned(865, 10), 350 => to_unsigned(265, 10), 351 => to_unsigned(850, 10), 352 => to_unsigned(351, 10), 353 => to_unsigned(766, 10), 354 => to_unsigned(545, 10), 355 => to_unsigned(49, 10), 356 => to_unsigned(498, 10), 357 => to_unsigned(158, 10), 358 => to_unsigned(454, 10), 359 => to_unsigned(575, 10), 360 => to_unsigned(269, 10), 361 => to_unsigned(510, 10), 362 => to_unsigned(648, 10), 363 => to_unsigned(455, 10), 364 => to_unsigned(802, 10), 365 => to_unsigned(280, 10), 366 => to_unsigned(3, 10), 367 => to_unsigned(661, 10), 368 => to_unsigned(941, 10), 369 => to_unsigned(131, 10), 370 => to_unsigned(248, 10), 371 => to_unsigned(729, 10), 372 => to_unsigned(171, 10), 373 => to_unsigned(567, 10), 374 => to_unsigned(227, 10), 375 => to_unsigned(423, 10), 376 => to_unsigned(358, 10), 377 => to_unsigned(193, 10), 378 => to_unsigned(786, 10), 379 => to_unsigned(102, 10), 380 => to_unsigned(215, 10), 381 => to_unsigned(497, 10), 382 => to_unsigned(608, 10), 383 => to_unsigned(395, 10), 384 => to_unsigned(673, 10), 385 => to_unsigned(1008, 10), 386 => to_unsigned(477, 10), 387 => to_unsigned(859, 10), 388 => to_unsigned(372, 10), 389 => to_unsigned(419, 10), 390 => to_unsigned(979, 10), 391 => to_unsigned(611, 10), 392 => to_unsigned(845, 10), 393 => to_unsigned(158, 10), 394 => to_unsigned(183, 10), 395 => to_unsigned(715, 10), 396 => to_unsigned(269, 10), 397 => to_unsigned(372, 10), 398 => to_unsigned(597, 10), 399 => to_unsigned(809, 10), 400 => to_unsigned(515, 10), 401 => to_unsigned(798, 10), 402 => to_unsigned(410, 10), 403 => to_unsigned(434, 10), 404 => to_unsigned(675, 10), 405 => to_unsigned(563, 10), 406 => to_unsigned(710, 10), 407 => to_unsigned(321, 10), 408 => to_unsigned(892, 10), 409 => to_unsigned(800, 10), 410 => to_unsigned(594, 10), 411 => to_unsigned(764, 10), 412 => to_unsigned(161, 10), 413 => to_unsigned(337, 10), 414 => to_unsigned(897, 10), 415 => to_unsigned(585, 10), 416 => to_unsigned(311, 10), 417 => to_unsigned(1005, 10), 418 => to_unsigned(836, 10), 419 => to_unsigned(423, 10), 420 => to_unsigned(97, 10), 421 => to_unsigned(136, 10), 422 => to_unsigned(646, 10), 423 => to_unsigned(368, 10), 424 => to_unsigned(904, 10), 425 => to_unsigned(297, 10), 426 => to_unsigned(617, 10), 427 => to_unsigned(941, 10), 428 => to_unsigned(599, 10), 429 => to_unsigned(320, 10), 430 => to_unsigned(7, 10), 431 => to_unsigned(400, 10), 432 => to_unsigned(653, 10), 433 => to_unsigned(589, 10), 434 => to_unsigned(428, 10), 435 => to_unsigned(866, 10), 436 => to_unsigned(149, 10), 437 => to_unsigned(431, 10), 438 => to_unsigned(288, 10), 439 => to_unsigned(229, 10), 440 => to_unsigned(475, 10), 441 => to_unsigned(888, 10), 442 => to_unsigned(841, 10), 443 => to_unsigned(281, 10), 444 => to_unsigned(891, 10), 445 => to_unsigned(206, 10), 446 => to_unsigned(179, 10), 447 => to_unsigned(1022, 10), 448 => to_unsigned(195, 10), 449 => to_unsigned(333, 10), 450 => to_unsigned(628, 10), 451 => to_unsigned(914, 10), 452 => to_unsigned(140, 10), 453 => to_unsigned(489, 10), 454 => to_unsigned(33, 10), 455 => to_unsigned(551, 10), 456 => to_unsigned(703, 10), 457 => to_unsigned(570, 10), 458 => to_unsigned(273, 10), 459 => to_unsigned(629, 10), 460 => to_unsigned(925, 10), 461 => to_unsigned(762, 10), 462 => to_unsigned(65, 10), 463 => to_unsigned(968, 10), 464 => to_unsigned(606, 10), 465 => to_unsigned(425, 10), 466 => to_unsigned(85, 10), 467 => to_unsigned(289, 10), 468 => to_unsigned(857, 10), 469 => to_unsigned(358, 10), 470 => to_unsigned(822, 10), 471 => to_unsigned(626, 10), 472 => to_unsigned(921, 10), 473 => to_unsigned(640, 10), 474 => to_unsigned(516, 10), 475 => to_unsigned(561, 10), 476 => to_unsigned(51, 10), 477 => to_unsigned(743, 10), 478 => to_unsigned(970, 10), 479 => to_unsigned(665, 10), 480 => to_unsigned(929, 10), 481 => to_unsigned(260, 10), 482 => to_unsigned(666, 10), 483 => to_unsigned(306, 10), 484 => to_unsigned(431, 10), 485 => to_unsigned(349, 10), 486 => to_unsigned(682, 10), 487 => to_unsigned(460, 10), 488 => to_unsigned(440, 10), 489 => to_unsigned(515, 10), 490 => to_unsigned(167, 10), 491 => to_unsigned(926, 10), 492 => to_unsigned(86, 10), 493 => to_unsigned(266, 10), 494 => to_unsigned(929, 10), 495 => to_unsigned(272, 10), 496 => to_unsigned(321, 10), 497 => to_unsigned(294, 10), 498 => to_unsigned(365, 10), 499 => to_unsigned(783, 10), 500 => to_unsigned(125, 10), 501 => to_unsigned(546, 10), 502 => to_unsigned(216, 10), 503 => to_unsigned(976, 10), 504 => to_unsigned(712, 10), 505 => to_unsigned(962, 10), 506 => to_unsigned(554, 10), 507 => to_unsigned(334, 10), 508 => to_unsigned(746, 10), 509 => to_unsigned(519, 10), 510 => to_unsigned(184, 10), 511 => to_unsigned(938, 10), 512 => to_unsigned(253, 10), 513 => to_unsigned(853, 10), 514 => to_unsigned(709, 10), 515 => to_unsigned(513, 10), 516 => to_unsigned(741, 10), 517 => to_unsigned(74, 10), 518 => to_unsigned(544, 10), 519 => to_unsigned(584, 10), 520 => to_unsigned(262, 10), 521 => to_unsigned(873, 10), 522 => to_unsigned(9, 10), 523 => to_unsigned(50, 10), 524 => to_unsigned(303, 10), 525 => to_unsigned(157, 10), 526 => to_unsigned(204, 10), 527 => to_unsigned(786, 10), 528 => to_unsigned(155, 10), 529 => to_unsigned(1006, 10), 530 => to_unsigned(916, 10), 531 => to_unsigned(580, 10), 532 => to_unsigned(748, 10), 533 => to_unsigned(254, 10), 534 => to_unsigned(395, 10), 535 => to_unsigned(80, 10), 536 => to_unsigned(361, 10), 537 => to_unsigned(39, 10), 538 => to_unsigned(644, 10), 539 => to_unsigned(49, 10), 540 => to_unsigned(687, 10), 541 => to_unsigned(870, 10), 542 => to_unsigned(463, 10), 543 => to_unsigned(92, 10), 544 => to_unsigned(981, 10), 545 => to_unsigned(726, 10), 546 => to_unsigned(903, 10), 547 => to_unsigned(227, 10), 548 => to_unsigned(465, 10), 549 => to_unsigned(389, 10), 550 => to_unsigned(1020, 10), 551 => to_unsigned(187, 10), 552 => to_unsigned(953, 10), 553 => to_unsigned(528, 10), 554 => to_unsigned(536, 10), 555 => to_unsigned(929, 10), 556 => to_unsigned(722, 10), 557 => to_unsigned(140, 10), 558 => to_unsigned(592, 10), 559 => to_unsigned(959, 10), 560 => to_unsigned(777, 10), 561 => to_unsigned(546, 10), 562 => to_unsigned(823, 10), 563 => to_unsigned(864, 10), 564 => to_unsigned(217, 10), 565 => to_unsigned(153, 10), 566 => to_unsigned(570, 10), 567 => to_unsigned(159, 10), 568 => to_unsigned(676, 10), 569 => to_unsigned(95, 10), 570 => to_unsigned(972, 10), 571 => to_unsigned(12, 10), 572 => to_unsigned(338, 10), 573 => to_unsigned(242, 10), 574 => to_unsigned(935, 10), 575 => to_unsigned(842, 10), 576 => to_unsigned(582, 10), 577 => to_unsigned(188, 10), 578 => to_unsigned(409, 10), 579 => to_unsigned(122, 10), 580 => to_unsigned(775, 10), 581 => to_unsigned(776, 10), 582 => to_unsigned(511, 10), 583 => to_unsigned(176, 10), 584 => to_unsigned(805, 10), 585 => to_unsigned(173, 10), 586 => to_unsigned(385, 10), 587 => to_unsigned(506, 10), 588 => to_unsigned(122, 10), 589 => to_unsigned(835, 10), 590 => to_unsigned(711, 10), 591 => to_unsigned(535, 10), 592 => to_unsigned(611, 10), 593 => to_unsigned(599, 10), 594 => to_unsigned(130, 10), 595 => to_unsigned(721, 10), 596 => to_unsigned(15, 10), 597 => to_unsigned(638, 10), 598 => to_unsigned(361, 10), 599 => to_unsigned(142, 10), 600 => to_unsigned(331, 10), 601 => to_unsigned(235, 10), 602 => to_unsigned(484, 10), 603 => to_unsigned(785, 10), 604 => to_unsigned(437, 10), 605 => to_unsigned(742, 10), 606 => to_unsigned(800, 10), 607 => to_unsigned(311, 10), 608 => to_unsigned(573, 10), 609 => to_unsigned(805, 10), 610 => to_unsigned(260, 10), 611 => to_unsigned(271, 10), 612 => to_unsigned(838, 10), 613 => to_unsigned(326, 10), 614 => to_unsigned(628, 10), 615 => to_unsigned(569, 10), 616 => to_unsigned(342, 10), 617 => to_unsigned(785, 10), 618 => to_unsigned(592, 10), 619 => to_unsigned(67, 10), 620 => to_unsigned(576, 10), 621 => to_unsigned(478, 10), 622 => to_unsigned(415, 10), 623 => to_unsigned(875, 10), 624 => to_unsigned(799, 10), 625 => to_unsigned(787, 10), 626 => to_unsigned(845, 10), 627 => to_unsigned(500, 10), 628 => to_unsigned(126, 10), 629 => to_unsigned(173, 10), 630 => to_unsigned(350, 10), 631 => to_unsigned(451, 10), 632 => to_unsigned(310, 10), 633 => to_unsigned(986, 10), 634 => to_unsigned(837, 10), 635 => to_unsigned(54, 10), 636 => to_unsigned(822, 10), 637 => to_unsigned(832, 10), 638 => to_unsigned(123, 10), 639 => to_unsigned(76, 10), 640 => to_unsigned(45, 10), 641 => to_unsigned(688, 10), 642 => to_unsigned(261, 10), 643 => to_unsigned(1001, 10), 644 => to_unsigned(653, 10), 645 => to_unsigned(237, 10), 646 => to_unsigned(351, 10), 647 => to_unsigned(587, 10), 648 => to_unsigned(44, 10), 649 => to_unsigned(96, 10), 650 => to_unsigned(975, 10), 651 => to_unsigned(672, 10), 652 => to_unsigned(295, 10), 653 => to_unsigned(691, 10), 654 => to_unsigned(307, 10), 655 => to_unsigned(699, 10), 656 => to_unsigned(1012, 10), 657 => to_unsigned(476, 10), 658 => to_unsigned(626, 10), 659 => to_unsigned(879, 10), 660 => to_unsigned(800, 10), 661 => to_unsigned(582, 10), 662 => to_unsigned(522, 10), 663 => to_unsigned(731, 10), 664 => to_unsigned(468, 10), 665 => to_unsigned(988, 10), 666 => to_unsigned(104, 10), 667 => to_unsigned(106, 10), 668 => to_unsigned(204, 10), 669 => to_unsigned(429, 10), 670 => to_unsigned(72, 10), 671 => to_unsigned(386, 10), 672 => to_unsigned(732, 10), 673 => to_unsigned(45, 10), 674 => to_unsigned(552, 10), 675 => to_unsigned(300, 10), 676 => to_unsigned(493, 10), 677 => to_unsigned(492, 10), 678 => to_unsigned(145, 10), 679 => to_unsigned(202, 10), 680 => to_unsigned(518, 10), 681 => to_unsigned(386, 10), 682 => to_unsigned(344, 10), 683 => to_unsigned(286, 10), 684 => to_unsigned(412, 10), 685 => to_unsigned(446, 10), 686 => to_unsigned(872, 10), 687 => to_unsigned(219, 10), 688 => to_unsigned(470, 10), 689 => to_unsigned(652, 10), 690 => to_unsigned(452, 10), 691 => to_unsigned(787, 10), 692 => to_unsigned(601, 10), 693 => to_unsigned(434, 10), 694 => to_unsigned(535, 10), 695 => to_unsigned(97, 10), 696 => to_unsigned(42, 10), 697 => to_unsigned(619, 10), 698 => to_unsigned(429, 10), 699 => to_unsigned(14, 10), 700 => to_unsigned(603, 10), 701 => to_unsigned(852, 10), 702 => to_unsigned(400, 10), 703 => to_unsigned(933, 10), 704 => to_unsigned(411, 10), 705 => to_unsigned(727, 10), 706 => to_unsigned(881, 10), 707 => to_unsigned(152, 10), 708 => to_unsigned(629, 10), 709 => to_unsigned(519, 10), 710 => to_unsigned(403, 10), 711 => to_unsigned(113, 10), 712 => to_unsigned(607, 10), 713 => to_unsigned(306, 10), 714 => to_unsigned(835, 10), 715 => to_unsigned(302, 10), 716 => to_unsigned(1010, 10), 717 => to_unsigned(678, 10), 718 => to_unsigned(186, 10), 719 => to_unsigned(492, 10), 720 => to_unsigned(817, 10), 721 => to_unsigned(504, 10), 722 => to_unsigned(68, 10), 723 => to_unsigned(576, 10), 724 => to_unsigned(354, 10), 725 => to_unsigned(111, 10), 726 => to_unsigned(675, 10), 727 => to_unsigned(620, 10), 728 => to_unsigned(306, 10), 729 => to_unsigned(847, 10), 730 => to_unsigned(458, 10), 731 => to_unsigned(600, 10), 732 => to_unsigned(576, 10), 733 => to_unsigned(860, 10), 734 => to_unsigned(807, 10), 735 => to_unsigned(942, 10), 736 => to_unsigned(891, 10), 737 => to_unsigned(159, 10), 738 => to_unsigned(168, 10), 739 => to_unsigned(783, 10), 740 => to_unsigned(710, 10), 741 => to_unsigned(51, 10), 742 => to_unsigned(448, 10), 743 => to_unsigned(371, 10), 744 => to_unsigned(690, 10), 745 => to_unsigned(851, 10), 746 => to_unsigned(423, 10), 747 => to_unsigned(235, 10), 748 => to_unsigned(459, 10), 749 => to_unsigned(980, 10), 750 => to_unsigned(571, 10), 751 => to_unsigned(338, 10), 752 => to_unsigned(148, 10), 753 => to_unsigned(308, 10), 754 => to_unsigned(116, 10), 755 => to_unsigned(344, 10), 756 => to_unsigned(498, 10), 757 => to_unsigned(803, 10), 758 => to_unsigned(777, 10), 759 => to_unsigned(24, 10), 760 => to_unsigned(454, 10), 761 => to_unsigned(276, 10), 762 => to_unsigned(798, 10), 763 => to_unsigned(671, 10), 764 => to_unsigned(392, 10), 765 => to_unsigned(207, 10), 766 => to_unsigned(179, 10), 767 => to_unsigned(826, 10), 768 => to_unsigned(313, 10), 769 => to_unsigned(730, 10), 770 => to_unsigned(405, 10), 771 => to_unsigned(642, 10), 772 => to_unsigned(847, 10), 773 => to_unsigned(384, 10), 774 => to_unsigned(29, 10), 775 => to_unsigned(405, 10), 776 => to_unsigned(812, 10), 777 => to_unsigned(301, 10), 778 => to_unsigned(964, 10), 779 => to_unsigned(648, 10), 780 => to_unsigned(223, 10), 781 => to_unsigned(674, 10), 782 => to_unsigned(173, 10), 783 => to_unsigned(52, 10), 784 => to_unsigned(595, 10), 785 => to_unsigned(337, 10), 786 => to_unsigned(694, 10), 787 => to_unsigned(785, 10), 788 => to_unsigned(957, 10), 789 => to_unsigned(291, 10), 790 => to_unsigned(792, 10), 791 => to_unsigned(929, 10), 792 => to_unsigned(511, 10), 793 => to_unsigned(131, 10), 794 => to_unsigned(972, 10), 795 => to_unsigned(216, 10), 796 => to_unsigned(804, 10), 797 => to_unsigned(297, 10), 798 => to_unsigned(147, 10), 799 => to_unsigned(260, 10), 800 => to_unsigned(488, 10), 801 => to_unsigned(695, 10), 802 => to_unsigned(634, 10), 803 => to_unsigned(1002, 10), 804 => to_unsigned(642, 10), 805 => to_unsigned(454, 10), 806 => to_unsigned(596, 10), 807 => to_unsigned(490, 10), 808 => to_unsigned(646, 10), 809 => to_unsigned(127, 10), 810 => to_unsigned(664, 10), 811 => to_unsigned(623, 10), 812 => to_unsigned(588, 10), 813 => to_unsigned(971, 10), 814 => to_unsigned(465, 10), 815 => to_unsigned(31, 10), 816 => to_unsigned(100, 10), 817 => to_unsigned(212, 10), 818 => to_unsigned(648, 10), 819 => to_unsigned(646, 10), 820 => to_unsigned(581, 10), 821 => to_unsigned(386, 10), 822 => to_unsigned(492, 10), 823 => to_unsigned(144, 10), 824 => to_unsigned(113, 10), 825 => to_unsigned(12, 10), 826 => to_unsigned(551, 10), 827 => to_unsigned(390, 10), 828 => to_unsigned(981, 10), 829 => to_unsigned(170, 10), 830 => to_unsigned(87, 10), 831 => to_unsigned(31, 10), 832 => to_unsigned(631, 10), 833 => to_unsigned(146, 10), 834 => to_unsigned(696, 10), 835 => to_unsigned(97, 10), 836 => to_unsigned(122, 10), 837 => to_unsigned(160, 10), 838 => to_unsigned(677, 10), 839 => to_unsigned(828, 10), 840 => to_unsigned(509, 10), 841 => to_unsigned(871, 10), 842 => to_unsigned(889, 10), 843 => to_unsigned(409, 10), 844 => to_unsigned(863, 10), 845 => to_unsigned(229, 10), 846 => to_unsigned(601, 10), 847 => to_unsigned(991, 10), 848 => to_unsigned(172, 10), 849 => to_unsigned(779, 10), 850 => to_unsigned(246, 10), 851 => to_unsigned(628, 10), 852 => to_unsigned(640, 10), 853 => to_unsigned(354, 10), 854 => to_unsigned(474, 10), 855 => to_unsigned(982, 10), 856 => to_unsigned(269, 10), 857 => to_unsigned(508, 10), 858 => to_unsigned(728, 10), 859 => to_unsigned(514, 10), 860 => to_unsigned(898, 10), 861 => to_unsigned(115, 10), 862 => to_unsigned(636, 10), 863 => to_unsigned(156, 10), 864 => to_unsigned(557, 10), 865 => to_unsigned(334, 10), 866 => to_unsigned(319, 10), 867 => to_unsigned(719, 10), 868 => to_unsigned(155, 10), 869 => to_unsigned(66, 10), 870 => to_unsigned(440, 10), 871 => to_unsigned(81, 10), 872 => to_unsigned(560, 10), 873 => to_unsigned(136, 10), 874 => to_unsigned(475, 10), 875 => to_unsigned(319, 10), 876 => to_unsigned(632, 10), 877 => to_unsigned(990, 10), 878 => to_unsigned(773, 10), 879 => to_unsigned(573, 10), 880 => to_unsigned(667, 10), 881 => to_unsigned(504, 10), 882 => to_unsigned(1022, 10), 883 => to_unsigned(41, 10), 884 => to_unsigned(146, 10), 885 => to_unsigned(145, 10), 886 => to_unsigned(704, 10), 887 => to_unsigned(964, 10), 888 => to_unsigned(97, 10), 889 => to_unsigned(102, 10), 890 => to_unsigned(361, 10), 891 => to_unsigned(908, 10), 892 => to_unsigned(994, 10), 893 => to_unsigned(890, 10), 894 => to_unsigned(726, 10), 895 => to_unsigned(154, 10), 896 => to_unsigned(268, 10), 897 => to_unsigned(205, 10), 898 => to_unsigned(249, 10), 899 => to_unsigned(352, 10), 900 => to_unsigned(883, 10), 901 => to_unsigned(320, 10), 902 => to_unsigned(791, 10), 903 => to_unsigned(219, 10), 904 => to_unsigned(268, 10), 905 => to_unsigned(974, 10), 906 => to_unsigned(284, 10), 907 => to_unsigned(52, 10), 908 => to_unsigned(195, 10), 909 => to_unsigned(153, 10), 910 => to_unsigned(890, 10), 911 => to_unsigned(839, 10), 912 => to_unsigned(320, 10), 913 => to_unsigned(341, 10), 914 => to_unsigned(752, 10), 915 => to_unsigned(10, 10), 916 => to_unsigned(968, 10), 917 => to_unsigned(116, 10), 918 => to_unsigned(107, 10), 919 => to_unsigned(915, 10), 920 => to_unsigned(138, 10), 921 => to_unsigned(161, 10), 922 => to_unsigned(765, 10), 923 => to_unsigned(524, 10), 924 => to_unsigned(380, 10), 925 => to_unsigned(540, 10), 926 => to_unsigned(925, 10), 927 => to_unsigned(320, 10), 928 => to_unsigned(223, 10), 929 => to_unsigned(436, 10), 930 => to_unsigned(934, 10), 931 => to_unsigned(310, 10), 932 => to_unsigned(776, 10), 933 => to_unsigned(747, 10), 934 => to_unsigned(661, 10), 935 => to_unsigned(493, 10), 936 => to_unsigned(864, 10), 937 => to_unsigned(919, 10), 938 => to_unsigned(600, 10), 939 => to_unsigned(381, 10), 940 => to_unsigned(122, 10), 941 => to_unsigned(646, 10), 942 => to_unsigned(910, 10), 943 => to_unsigned(293, 10), 944 => to_unsigned(463, 10), 945 => to_unsigned(475, 10), 946 => to_unsigned(256, 10), 947 => to_unsigned(837, 10), 948 => to_unsigned(668, 10), 949 => to_unsigned(847, 10), 950 => to_unsigned(421, 10), 951 => to_unsigned(833, 10), 952 => to_unsigned(461, 10), 953 => to_unsigned(174, 10), 954 => to_unsigned(81, 10), 955 => to_unsigned(122, 10), 956 => to_unsigned(546, 10), 957 => to_unsigned(23, 10), 958 => to_unsigned(827, 10), 959 => to_unsigned(101, 10), 960 => to_unsigned(182, 10), 961 => to_unsigned(564, 10), 962 => to_unsigned(915, 10), 963 => to_unsigned(879, 10), 964 => to_unsigned(207, 10), 965 => to_unsigned(344, 10), 966 => to_unsigned(650, 10), 967 => to_unsigned(120, 10), 968 => to_unsigned(721, 10), 969 => to_unsigned(846, 10), 970 => to_unsigned(271, 10), 971 => to_unsigned(231, 10), 972 => to_unsigned(752, 10), 973 => to_unsigned(944, 10), 974 => to_unsigned(441, 10), 975 => to_unsigned(991, 10), 976 => to_unsigned(209, 10), 977 => to_unsigned(438, 10), 978 => to_unsigned(708, 10), 979 => to_unsigned(170, 10), 980 => to_unsigned(426, 10), 981 => to_unsigned(655, 10), 982 => to_unsigned(940, 10), 983 => to_unsigned(841, 10), 984 => to_unsigned(419, 10), 985 => to_unsigned(498, 10), 986 => to_unsigned(404, 10), 987 => to_unsigned(375, 10), 988 => to_unsigned(116, 10), 989 => to_unsigned(796, 10), 990 => to_unsigned(773, 10), 991 => to_unsigned(776, 10), 992 => to_unsigned(264, 10), 993 => to_unsigned(214, 10), 994 => to_unsigned(314, 10), 995 => to_unsigned(891, 10), 996 => to_unsigned(215, 10), 997 => to_unsigned(677, 10), 998 => to_unsigned(956, 10), 999 => to_unsigned(632, 10), 1000 => to_unsigned(817, 10), 1001 => to_unsigned(896, 10), 1002 => to_unsigned(217, 10), 1003 => to_unsigned(523, 10), 1004 => to_unsigned(166, 10), 1005 => to_unsigned(243, 10), 1006 => to_unsigned(702, 10), 1007 => to_unsigned(836, 10), 1008 => to_unsigned(677, 10), 1009 => to_unsigned(492, 10), 1010 => to_unsigned(103, 10), 1011 => to_unsigned(531, 10), 1012 => to_unsigned(242, 10), 1013 => to_unsigned(389, 10), 1014 => to_unsigned(181, 10), 1015 => to_unsigned(8, 10), 1016 => to_unsigned(541, 10), 1017 => to_unsigned(314, 10), 1018 => to_unsigned(501, 10), 1019 => to_unsigned(1009, 10), 1020 => to_unsigned(985, 10), 1021 => to_unsigned(191, 10), 1022 => to_unsigned(928, 10), 1023 => to_unsigned(286, 10), 1024 => to_unsigned(328, 10), 1025 => to_unsigned(768, 10), 1026 => to_unsigned(182, 10), 1027 => to_unsigned(916, 10), 1028 => to_unsigned(494, 10), 1029 => to_unsigned(1010, 10), 1030 => to_unsigned(538, 10), 1031 => to_unsigned(388, 10), 1032 => to_unsigned(840, 10), 1033 => to_unsigned(52, 10), 1034 => to_unsigned(267, 10), 1035 => to_unsigned(371, 10), 1036 => to_unsigned(228, 10), 1037 => to_unsigned(862, 10), 1038 => to_unsigned(360, 10), 1039 => to_unsigned(425, 10), 1040 => to_unsigned(477, 10), 1041 => to_unsigned(487, 10), 1042 => to_unsigned(730, 10), 1043 => to_unsigned(848, 10), 1044 => to_unsigned(629, 10), 1045 => to_unsigned(404, 10), 1046 => to_unsigned(591, 10), 1047 => to_unsigned(331, 10), 1048 => to_unsigned(732, 10), 1049 => to_unsigned(947, 10), 1050 => to_unsigned(971, 10), 1051 => to_unsigned(652, 10), 1052 => to_unsigned(55, 10), 1053 => to_unsigned(100, 10), 1054 => to_unsigned(830, 10), 1055 => to_unsigned(352, 10), 1056 => to_unsigned(779, 10), 1057 => to_unsigned(883, 10), 1058 => to_unsigned(834, 10), 1059 => to_unsigned(871, 10), 1060 => to_unsigned(201, 10), 1061 => to_unsigned(1009, 10), 1062 => to_unsigned(300, 10), 1063 => to_unsigned(10, 10), 1064 => to_unsigned(725, 10), 1065 => to_unsigned(885, 10), 1066 => to_unsigned(419, 10), 1067 => to_unsigned(372, 10), 1068 => to_unsigned(268, 10), 1069 => to_unsigned(653, 10), 1070 => to_unsigned(631, 10), 1071 => to_unsigned(127, 10), 1072 => to_unsigned(887, 10), 1073 => to_unsigned(763, 10), 1074 => to_unsigned(366, 10), 1075 => to_unsigned(303, 10), 1076 => to_unsigned(425, 10), 1077 => to_unsigned(115, 10), 1078 => to_unsigned(785, 10), 1079 => to_unsigned(675, 10), 1080 => to_unsigned(806, 10), 1081 => to_unsigned(187, 10), 1082 => to_unsigned(675, 10), 1083 => to_unsigned(1006, 10), 1084 => to_unsigned(610, 10), 1085 => to_unsigned(221, 10), 1086 => to_unsigned(39, 10), 1087 => to_unsigned(945, 10), 1088 => to_unsigned(440, 10), 1089 => to_unsigned(93, 10), 1090 => to_unsigned(85, 10), 1091 => to_unsigned(650, 10), 1092 => to_unsigned(75, 10), 1093 => to_unsigned(613, 10), 1094 => to_unsigned(116, 10), 1095 => to_unsigned(620, 10), 1096 => to_unsigned(583, 10), 1097 => to_unsigned(381, 10), 1098 => to_unsigned(789, 10), 1099 => to_unsigned(520, 10), 1100 => to_unsigned(595, 10), 1101 => to_unsigned(526, 10), 1102 => to_unsigned(938, 10), 1103 => to_unsigned(279, 10), 1104 => to_unsigned(501, 10), 1105 => to_unsigned(284, 10), 1106 => to_unsigned(538, 10), 1107 => to_unsigned(218, 10), 1108 => to_unsigned(715, 10), 1109 => to_unsigned(502, 10), 1110 => to_unsigned(996, 10), 1111 => to_unsigned(16, 10), 1112 => to_unsigned(571, 10), 1113 => to_unsigned(176, 10), 1114 => to_unsigned(174, 10), 1115 => to_unsigned(666, 10), 1116 => to_unsigned(128, 10), 1117 => to_unsigned(251, 10), 1118 => to_unsigned(688, 10), 1119 => to_unsigned(699, 10), 1120 => to_unsigned(172, 10), 1121 => to_unsigned(548, 10), 1122 => to_unsigned(290, 10), 1123 => to_unsigned(158, 10), 1124 => to_unsigned(887, 10), 1125 => to_unsigned(474, 10), 1126 => to_unsigned(166, 10), 1127 => to_unsigned(693, 10), 1128 => to_unsigned(279, 10), 1129 => to_unsigned(839, 10), 1130 => to_unsigned(840, 10), 1131 => to_unsigned(277, 10), 1132 => to_unsigned(821, 10), 1133 => to_unsigned(53, 10), 1134 => to_unsigned(587, 10), 1135 => to_unsigned(831, 10), 1136 => to_unsigned(80, 10), 1137 => to_unsigned(94, 10), 1138 => to_unsigned(670, 10), 1139 => to_unsigned(734, 10), 1140 => to_unsigned(954, 10), 1141 => to_unsigned(322, 10), 1142 => to_unsigned(904, 10), 1143 => to_unsigned(943, 10), 1144 => to_unsigned(347, 10), 1145 => to_unsigned(29, 10), 1146 => to_unsigned(718, 10), 1147 => to_unsigned(818, 10), 1148 => to_unsigned(693, 10), 1149 => to_unsigned(300, 10), 1150 => to_unsigned(730, 10), 1151 => to_unsigned(379, 10), 1152 => to_unsigned(248, 10), 1153 => to_unsigned(562, 10), 1154 => to_unsigned(741, 10), 1155 => to_unsigned(495, 10), 1156 => to_unsigned(700, 10), 1157 => to_unsigned(552, 10), 1158 => to_unsigned(636, 10), 1159 => to_unsigned(585, 10), 1160 => to_unsigned(807, 10), 1161 => to_unsigned(975, 10), 1162 => to_unsigned(508, 10), 1163 => to_unsigned(821, 10), 1164 => to_unsigned(25, 10), 1165 => to_unsigned(635, 10), 1166 => to_unsigned(182, 10), 1167 => to_unsigned(881, 10), 1168 => to_unsigned(746, 10), 1169 => to_unsigned(859, 10), 1170 => to_unsigned(959, 10), 1171 => to_unsigned(79, 10), 1172 => to_unsigned(285, 10), 1173 => to_unsigned(740, 10), 1174 => to_unsigned(865, 10), 1175 => to_unsigned(328, 10), 1176 => to_unsigned(475, 10), 1177 => to_unsigned(625, 10), 1178 => to_unsigned(358, 10), 1179 => to_unsigned(322, 10), 1180 => to_unsigned(784, 10), 1181 => to_unsigned(389, 10), 1182 => to_unsigned(272, 10), 1183 => to_unsigned(630, 10), 1184 => to_unsigned(757, 10), 1185 => to_unsigned(443, 10), 1186 => to_unsigned(461, 10), 1187 => to_unsigned(62, 10), 1188 => to_unsigned(118, 10), 1189 => to_unsigned(720, 10), 1190 => to_unsigned(319, 10), 1191 => to_unsigned(442, 10), 1192 => to_unsigned(472, 10), 1193 => to_unsigned(198, 10), 1194 => to_unsigned(903, 10), 1195 => to_unsigned(44, 10), 1196 => to_unsigned(310, 10), 1197 => to_unsigned(468, 10), 1198 => to_unsigned(665, 10), 1199 => to_unsigned(702, 10), 1200 => to_unsigned(599, 10), 1201 => to_unsigned(695, 10), 1202 => to_unsigned(848, 10), 1203 => to_unsigned(922, 10), 1204 => to_unsigned(678, 10), 1205 => to_unsigned(121, 10), 1206 => to_unsigned(980, 10), 1207 => to_unsigned(441, 10), 1208 => to_unsigned(610, 10), 1209 => to_unsigned(140, 10), 1210 => to_unsigned(888, 10), 1211 => to_unsigned(436, 10), 1212 => to_unsigned(562, 10), 1213 => to_unsigned(121, 10), 1214 => to_unsigned(799, 10), 1215 => to_unsigned(193, 10), 1216 => to_unsigned(453, 10), 1217 => to_unsigned(885, 10), 1218 => to_unsigned(1013, 10), 1219 => to_unsigned(483, 10), 1220 => to_unsigned(941, 10), 1221 => to_unsigned(393, 10), 1222 => to_unsigned(178, 10), 1223 => to_unsigned(555, 10), 1224 => to_unsigned(112, 10), 1225 => to_unsigned(601, 10), 1226 => to_unsigned(148, 10), 1227 => to_unsigned(299, 10), 1228 => to_unsigned(858, 10), 1229 => to_unsigned(441, 10), 1230 => to_unsigned(212, 10), 1231 => to_unsigned(125, 10), 1232 => to_unsigned(867, 10), 1233 => to_unsigned(829, 10), 1234 => to_unsigned(492, 10), 1235 => to_unsigned(958, 10), 1236 => to_unsigned(948, 10), 1237 => to_unsigned(834, 10), 1238 => to_unsigned(588, 10), 1239 => to_unsigned(657, 10), 1240 => to_unsigned(277, 10), 1241 => to_unsigned(294, 10), 1242 => to_unsigned(483, 10), 1243 => to_unsigned(125, 10), 1244 => to_unsigned(512, 10), 1245 => to_unsigned(331, 10), 1246 => to_unsigned(207, 10), 1247 => to_unsigned(690, 10), 1248 => to_unsigned(413, 10), 1249 => to_unsigned(603, 10), 1250 => to_unsigned(869, 10), 1251 => to_unsigned(305, 10), 1252 => to_unsigned(644, 10), 1253 => to_unsigned(954, 10), 1254 => to_unsigned(620, 10), 1255 => to_unsigned(641, 10), 1256 => to_unsigned(377, 10), 1257 => to_unsigned(978, 10), 1258 => to_unsigned(398, 10), 1259 => to_unsigned(326, 10), 1260 => to_unsigned(162, 10), 1261 => to_unsigned(194, 10), 1262 => to_unsigned(671, 10), 1263 => to_unsigned(111, 10), 1264 => to_unsigned(129, 10), 1265 => to_unsigned(313, 10), 1266 => to_unsigned(184, 10), 1267 => to_unsigned(140, 10), 1268 => to_unsigned(172, 10), 1269 => to_unsigned(109, 10), 1270 => to_unsigned(226, 10), 1271 => to_unsigned(283, 10), 1272 => to_unsigned(465, 10), 1273 => to_unsigned(244, 10), 1274 => to_unsigned(739, 10), 1275 => to_unsigned(892, 10), 1276 => to_unsigned(207, 10), 1277 => to_unsigned(987, 10), 1278 => to_unsigned(164, 10), 1279 => to_unsigned(525, 10), 1280 => to_unsigned(1003, 10), 1281 => to_unsigned(397, 10), 1282 => to_unsigned(168, 10), 1283 => to_unsigned(344, 10), 1284 => to_unsigned(459, 10), 1285 => to_unsigned(415, 10), 1286 => to_unsigned(488, 10), 1287 => to_unsigned(618, 10), 1288 => to_unsigned(280, 10), 1289 => to_unsigned(790, 10), 1290 => to_unsigned(948, 10), 1291 => to_unsigned(309, 10), 1292 => to_unsigned(930, 10), 1293 => to_unsigned(925, 10), 1294 => to_unsigned(722, 10), 1295 => to_unsigned(463, 10), 1296 => to_unsigned(202, 10), 1297 => to_unsigned(550, 10), 1298 => to_unsigned(458, 10), 1299 => to_unsigned(590, 10), 1300 => to_unsigned(472, 10), 1301 => to_unsigned(751, 10), 1302 => to_unsigned(962, 10), 1303 => to_unsigned(893, 10), 1304 => to_unsigned(884, 10), 1305 => to_unsigned(590, 10), 1306 => to_unsigned(367, 10), 1307 => to_unsigned(123, 10), 1308 => to_unsigned(996, 10), 1309 => to_unsigned(863, 10), 1310 => to_unsigned(249, 10), 1311 => to_unsigned(218, 10), 1312 => to_unsigned(762, 10), 1313 => to_unsigned(875, 10), 1314 => to_unsigned(540, 10), 1315 => to_unsigned(625, 10), 1316 => to_unsigned(286, 10), 1317 => to_unsigned(661, 10), 1318 => to_unsigned(863, 10), 1319 => to_unsigned(209, 10), 1320 => to_unsigned(383, 10), 1321 => to_unsigned(918, 10), 1322 => to_unsigned(133, 10), 1323 => to_unsigned(412, 10), 1324 => to_unsigned(525, 10), 1325 => to_unsigned(979, 10), 1326 => to_unsigned(946, 10), 1327 => to_unsigned(321, 10), 1328 => to_unsigned(0, 10), 1329 => to_unsigned(23, 10), 1330 => to_unsigned(874, 10), 1331 => to_unsigned(845, 10), 1332 => to_unsigned(929, 10), 1333 => to_unsigned(715, 10), 1334 => to_unsigned(203, 10), 1335 => to_unsigned(441, 10), 1336 => to_unsigned(909, 10), 1337 => to_unsigned(195, 10), 1338 => to_unsigned(107, 10), 1339 => to_unsigned(902, 10), 1340 => to_unsigned(446, 10), 1341 => to_unsigned(408, 10), 1342 => to_unsigned(987, 10), 1343 => to_unsigned(499, 10), 1344 => to_unsigned(181, 10), 1345 => to_unsigned(477, 10), 1346 => to_unsigned(337, 10), 1347 => to_unsigned(526, 10), 1348 => to_unsigned(495, 10), 1349 => to_unsigned(477, 10), 1350 => to_unsigned(32, 10), 1351 => to_unsigned(181, 10), 1352 => to_unsigned(5, 10), 1353 => to_unsigned(12, 10), 1354 => to_unsigned(77, 10), 1355 => to_unsigned(15, 10), 1356 => to_unsigned(290, 10), 1357 => to_unsigned(715, 10), 1358 => to_unsigned(239, 10), 1359 => to_unsigned(176, 10), 1360 => to_unsigned(683, 10), 1361 => to_unsigned(367, 10), 1362 => to_unsigned(104, 10), 1363 => to_unsigned(128, 10), 1364 => to_unsigned(66, 10), 1365 => to_unsigned(977, 10), 1366 => to_unsigned(530, 10), 1367 => to_unsigned(859, 10), 1368 => to_unsigned(285, 10), 1369 => to_unsigned(621, 10), 1370 => to_unsigned(644, 10), 1371 => to_unsigned(219, 10), 1372 => to_unsigned(849, 10), 1373 => to_unsigned(79, 10), 1374 => to_unsigned(885, 10), 1375 => to_unsigned(398, 10), 1376 => to_unsigned(1013, 10), 1377 => to_unsigned(677, 10), 1378 => to_unsigned(500, 10), 1379 => to_unsigned(128, 10), 1380 => to_unsigned(709, 10), 1381 => to_unsigned(691, 10), 1382 => to_unsigned(28, 10), 1383 => to_unsigned(126, 10), 1384 => to_unsigned(932, 10), 1385 => to_unsigned(801, 10), 1386 => to_unsigned(957, 10), 1387 => to_unsigned(378, 10), 1388 => to_unsigned(180, 10), 1389 => to_unsigned(989, 10), 1390 => to_unsigned(769, 10), 1391 => to_unsigned(878, 10), 1392 => to_unsigned(985, 10), 1393 => to_unsigned(301, 10), 1394 => to_unsigned(443, 10), 1395 => to_unsigned(683, 10), 1396 => to_unsigned(530, 10), 1397 => to_unsigned(600, 10), 1398 => to_unsigned(645, 10), 1399 => to_unsigned(963, 10), 1400 => to_unsigned(521, 10), 1401 => to_unsigned(954, 10), 1402 => to_unsigned(329, 10), 1403 => to_unsigned(378, 10), 1404 => to_unsigned(110, 10), 1405 => to_unsigned(709, 10), 1406 => to_unsigned(518, 10), 1407 => to_unsigned(2, 10), 1408 => to_unsigned(72, 10), 1409 => to_unsigned(558, 10), 1410 => to_unsigned(32, 10), 1411 => to_unsigned(764, 10), 1412 => to_unsigned(29, 10), 1413 => to_unsigned(614, 10), 1414 => to_unsigned(22, 10), 1415 => to_unsigned(208, 10), 1416 => to_unsigned(310, 10), 1417 => to_unsigned(246, 10), 1418 => to_unsigned(157, 10), 1419 => to_unsigned(854, 10), 1420 => to_unsigned(401, 10), 1421 => to_unsigned(443, 10), 1422 => to_unsigned(829, 10), 1423 => to_unsigned(873, 10), 1424 => to_unsigned(508, 10), 1425 => to_unsigned(34, 10), 1426 => to_unsigned(42, 10), 1427 => to_unsigned(95, 10), 1428 => to_unsigned(692, 10), 1429 => to_unsigned(844, 10), 1430 => to_unsigned(162, 10), 1431 => to_unsigned(214, 10), 1432 => to_unsigned(467, 10), 1433 => to_unsigned(834, 10), 1434 => to_unsigned(983, 10), 1435 => to_unsigned(129, 10), 1436 => to_unsigned(442, 10), 1437 => to_unsigned(986, 10), 1438 => to_unsigned(823, 10), 1439 => to_unsigned(253, 10), 1440 => to_unsigned(162, 10), 1441 => to_unsigned(85, 10), 1442 => to_unsigned(269, 10), 1443 => to_unsigned(183, 10), 1444 => to_unsigned(211, 10), 1445 => to_unsigned(535, 10), 1446 => to_unsigned(549, 10), 1447 => to_unsigned(285, 10), 1448 => to_unsigned(626, 10), 1449 => to_unsigned(961, 10), 1450 => to_unsigned(902, 10), 1451 => to_unsigned(761, 10), 1452 => to_unsigned(66, 10), 1453 => to_unsigned(92, 10), 1454 => to_unsigned(770, 10), 1455 => to_unsigned(562, 10), 1456 => to_unsigned(822, 10), 1457 => to_unsigned(521, 10), 1458 => to_unsigned(965, 10), 1459 => to_unsigned(361, 10), 1460 => to_unsigned(103, 10), 1461 => to_unsigned(601, 10), 1462 => to_unsigned(788, 10), 1463 => to_unsigned(476, 10), 1464 => to_unsigned(992, 10), 1465 => to_unsigned(822, 10), 1466 => to_unsigned(748, 10), 1467 => to_unsigned(682, 10), 1468 => to_unsigned(346, 10), 1469 => to_unsigned(110, 10), 1470 => to_unsigned(913, 10), 1471 => to_unsigned(707, 10), 1472 => to_unsigned(575, 10), 1473 => to_unsigned(538, 10), 1474 => to_unsigned(78, 10), 1475 => to_unsigned(380, 10), 1476 => to_unsigned(728, 10), 1477 => to_unsigned(96, 10), 1478 => to_unsigned(220, 10), 1479 => to_unsigned(573, 10), 1480 => to_unsigned(692, 10), 1481 => to_unsigned(147, 10), 1482 => to_unsigned(932, 10), 1483 => to_unsigned(875, 10), 1484 => to_unsigned(349, 10), 1485 => to_unsigned(518, 10), 1486 => to_unsigned(360, 10), 1487 => to_unsigned(610, 10), 1488 => to_unsigned(1006, 10), 1489 => to_unsigned(544, 10), 1490 => to_unsigned(1022, 10), 1491 => to_unsigned(739, 10), 1492 => to_unsigned(959, 10), 1493 => to_unsigned(894, 10), 1494 => to_unsigned(604, 10), 1495 => to_unsigned(212, 10), 1496 => to_unsigned(405, 10), 1497 => to_unsigned(875, 10), 1498 => to_unsigned(399, 10), 1499 => to_unsigned(668, 10), 1500 => to_unsigned(154, 10), 1501 => to_unsigned(267, 10), 1502 => to_unsigned(779, 10), 1503 => to_unsigned(133, 10), 1504 => to_unsigned(120, 10), 1505 => to_unsigned(271, 10), 1506 => to_unsigned(546, 10), 1507 => to_unsigned(589, 10), 1508 => to_unsigned(843, 10), 1509 => to_unsigned(631, 10), 1510 => to_unsigned(328, 10), 1511 => to_unsigned(874, 10), 1512 => to_unsigned(361, 10), 1513 => to_unsigned(537, 10), 1514 => to_unsigned(19, 10), 1515 => to_unsigned(709, 10), 1516 => to_unsigned(627, 10), 1517 => to_unsigned(64, 10), 1518 => to_unsigned(460, 10), 1519 => to_unsigned(649, 10), 1520 => to_unsigned(128, 10), 1521 => to_unsigned(567, 10), 1522 => to_unsigned(802, 10), 1523 => to_unsigned(772, 10), 1524 => to_unsigned(240, 10), 1525 => to_unsigned(521, 10), 1526 => to_unsigned(747, 10), 1527 => to_unsigned(841, 10), 1528 => to_unsigned(817, 10), 1529 => to_unsigned(878, 10), 1530 => to_unsigned(906, 10), 1531 => to_unsigned(491, 10), 1532 => to_unsigned(231, 10), 1533 => to_unsigned(767, 10), 1534 => to_unsigned(1015, 10), 1535 => to_unsigned(469, 10), 1536 => to_unsigned(699, 10), 1537 => to_unsigned(681, 10), 1538 => to_unsigned(296, 10), 1539 => to_unsigned(880, 10), 1540 => to_unsigned(669, 10), 1541 => to_unsigned(700, 10), 1542 => to_unsigned(478, 10), 1543 => to_unsigned(877, 10), 1544 => to_unsigned(517, 10), 1545 => to_unsigned(852, 10), 1546 => to_unsigned(658, 10), 1547 => to_unsigned(149, 10), 1548 => to_unsigned(119, 10), 1549 => to_unsigned(706, 10), 1550 => to_unsigned(531, 10), 1551 => to_unsigned(769, 10), 1552 => to_unsigned(918, 10), 1553 => to_unsigned(624, 10), 1554 => to_unsigned(809, 10), 1555 => to_unsigned(778, 10), 1556 => to_unsigned(916, 10), 1557 => to_unsigned(702, 10), 1558 => to_unsigned(583, 10), 1559 => to_unsigned(112, 10), 1560 => to_unsigned(311, 10), 1561 => to_unsigned(602, 10), 1562 => to_unsigned(663, 10), 1563 => to_unsigned(40, 10), 1564 => to_unsigned(618, 10), 1565 => to_unsigned(611, 10), 1566 => to_unsigned(239, 10), 1567 => to_unsigned(377, 10), 1568 => to_unsigned(584, 10), 1569 => to_unsigned(418, 10), 1570 => to_unsigned(667, 10), 1571 => to_unsigned(4, 10), 1572 => to_unsigned(452, 10), 1573 => to_unsigned(530, 10), 1574 => to_unsigned(649, 10), 1575 => to_unsigned(232, 10), 1576 => to_unsigned(903, 10), 1577 => to_unsigned(946, 10), 1578 => to_unsigned(30, 10), 1579 => to_unsigned(462, 10), 1580 => to_unsigned(340, 10), 1581 => to_unsigned(189, 10), 1582 => to_unsigned(253, 10), 1583 => to_unsigned(315, 10), 1584 => to_unsigned(1014, 10), 1585 => to_unsigned(213, 10), 1586 => to_unsigned(794, 10), 1587 => to_unsigned(757, 10), 1588 => to_unsigned(99, 10), 1589 => to_unsigned(199, 10), 1590 => to_unsigned(238, 10), 1591 => to_unsigned(198, 10), 1592 => to_unsigned(395, 10), 1593 => to_unsigned(220, 10), 1594 => to_unsigned(762, 10), 1595 => to_unsigned(623, 10), 1596 => to_unsigned(423, 10), 1597 => to_unsigned(839, 10), 1598 => to_unsigned(671, 10), 1599 => to_unsigned(497, 10), 1600 => to_unsigned(635, 10), 1601 => to_unsigned(443, 10), 1602 => to_unsigned(79, 10), 1603 => to_unsigned(906, 10), 1604 => to_unsigned(412, 10), 1605 => to_unsigned(116, 10), 1606 => to_unsigned(390, 10), 1607 => to_unsigned(857, 10), 1608 => to_unsigned(794, 10), 1609 => to_unsigned(54, 10), 1610 => to_unsigned(273, 10), 1611 => to_unsigned(487, 10), 1612 => to_unsigned(12, 10), 1613 => to_unsigned(602, 10), 1614 => to_unsigned(355, 10), 1615 => to_unsigned(578, 10), 1616 => to_unsigned(765, 10), 1617 => to_unsigned(67, 10), 1618 => to_unsigned(668, 10), 1619 => to_unsigned(451, 10), 1620 => to_unsigned(354, 10), 1621 => to_unsigned(891, 10), 1622 => to_unsigned(950, 10), 1623 => to_unsigned(20, 10), 1624 => to_unsigned(240, 10), 1625 => to_unsigned(257, 10), 1626 => to_unsigned(615, 10), 1627 => to_unsigned(212, 10), 1628 => to_unsigned(222, 10), 1629 => to_unsigned(416, 10), 1630 => to_unsigned(669, 10), 1631 => to_unsigned(15, 10), 1632 => to_unsigned(6, 10), 1633 => to_unsigned(809, 10), 1634 => to_unsigned(266, 10), 1635 => to_unsigned(474, 10), 1636 => to_unsigned(773, 10), 1637 => to_unsigned(783, 10), 1638 => to_unsigned(220, 10), 1639 => to_unsigned(835, 10), 1640 => to_unsigned(125, 10), 1641 => to_unsigned(827, 10), 1642 => to_unsigned(565, 10), 1643 => to_unsigned(983, 10), 1644 => to_unsigned(762, 10), 1645 => to_unsigned(200, 10), 1646 => to_unsigned(938, 10), 1647 => to_unsigned(91, 10), 1648 => to_unsigned(632, 10), 1649 => to_unsigned(37, 10), 1650 => to_unsigned(537, 10), 1651 => to_unsigned(114, 10), 1652 => to_unsigned(657, 10), 1653 => to_unsigned(352, 10), 1654 => to_unsigned(983, 10), 1655 => to_unsigned(78, 10), 1656 => to_unsigned(719, 10), 1657 => to_unsigned(71, 10), 1658 => to_unsigned(213, 10), 1659 => to_unsigned(157, 10), 1660 => to_unsigned(636, 10), 1661 => to_unsigned(545, 10), 1662 => to_unsigned(455, 10), 1663 => to_unsigned(983, 10), 1664 => to_unsigned(387, 10), 1665 => to_unsigned(771, 10), 1666 => to_unsigned(258, 10), 1667 => to_unsigned(867, 10), 1668 => to_unsigned(900, 10), 1669 => to_unsigned(190, 10), 1670 => to_unsigned(794, 10), 1671 => to_unsigned(393, 10), 1672 => to_unsigned(591, 10), 1673 => to_unsigned(0, 10), 1674 => to_unsigned(848, 10), 1675 => to_unsigned(472, 10), 1676 => to_unsigned(444, 10), 1677 => to_unsigned(756, 10), 1678 => to_unsigned(840, 10), 1679 => to_unsigned(913, 10), 1680 => to_unsigned(2, 10), 1681 => to_unsigned(36, 10), 1682 => to_unsigned(11, 10), 1683 => to_unsigned(328, 10), 1684 => to_unsigned(439, 10), 1685 => to_unsigned(786, 10), 1686 => to_unsigned(666, 10), 1687 => to_unsigned(919, 10), 1688 => to_unsigned(908, 10), 1689 => to_unsigned(915, 10), 1690 => to_unsigned(935, 10), 1691 => to_unsigned(223, 10), 1692 => to_unsigned(765, 10), 1693 => to_unsigned(774, 10), 1694 => to_unsigned(562, 10), 1695 => to_unsigned(985, 10), 1696 => to_unsigned(761, 10), 1697 => to_unsigned(268, 10), 1698 => to_unsigned(832, 10), 1699 => to_unsigned(570, 10), 1700 => to_unsigned(418, 10), 1701 => to_unsigned(931, 10), 1702 => to_unsigned(246, 10), 1703 => to_unsigned(680, 10), 1704 => to_unsigned(1022, 10), 1705 => to_unsigned(386, 10), 1706 => to_unsigned(230, 10), 1707 => to_unsigned(192, 10), 1708 => to_unsigned(580, 10), 1709 => to_unsigned(69, 10), 1710 => to_unsigned(867, 10), 1711 => to_unsigned(484, 10), 1712 => to_unsigned(73, 10), 1713 => to_unsigned(173, 10), 1714 => to_unsigned(849, 10), 1715 => to_unsigned(733, 10), 1716 => to_unsigned(320, 10), 1717 => to_unsigned(524, 10), 1718 => to_unsigned(180, 10), 1719 => to_unsigned(95, 10), 1720 => to_unsigned(751, 10), 1721 => to_unsigned(18, 10), 1722 => to_unsigned(835, 10), 1723 => to_unsigned(525, 10), 1724 => to_unsigned(514, 10), 1725 => to_unsigned(208, 10), 1726 => to_unsigned(277, 10), 1727 => to_unsigned(169, 10), 1728 => to_unsigned(88, 10), 1729 => to_unsigned(302, 10), 1730 => to_unsigned(392, 10), 1731 => to_unsigned(434, 10), 1732 => to_unsigned(304, 10), 1733 => to_unsigned(495, 10), 1734 => to_unsigned(874, 10), 1735 => to_unsigned(932, 10), 1736 => to_unsigned(59, 10), 1737 => to_unsigned(356, 10), 1738 => to_unsigned(987, 10), 1739 => to_unsigned(602, 10), 1740 => to_unsigned(910, 10), 1741 => to_unsigned(424, 10), 1742 => to_unsigned(644, 10), 1743 => to_unsigned(547, 10), 1744 => to_unsigned(66, 10), 1745 => to_unsigned(403, 10), 1746 => to_unsigned(28, 10), 1747 => to_unsigned(18, 10), 1748 => to_unsigned(588, 10), 1749 => to_unsigned(791, 10), 1750 => to_unsigned(847, 10), 1751 => to_unsigned(110, 10), 1752 => to_unsigned(683, 10), 1753 => to_unsigned(143, 10), 1754 => to_unsigned(382, 10), 1755 => to_unsigned(482, 10), 1756 => to_unsigned(102, 10), 1757 => to_unsigned(813, 10), 1758 => to_unsigned(97, 10), 1759 => to_unsigned(756, 10), 1760 => to_unsigned(443, 10), 1761 => to_unsigned(666, 10), 1762 => to_unsigned(25, 10), 1763 => to_unsigned(167, 10), 1764 => to_unsigned(193, 10), 1765 => to_unsigned(703, 10), 1766 => to_unsigned(170, 10), 1767 => to_unsigned(850, 10), 1768 => to_unsigned(621, 10), 1769 => to_unsigned(971, 10), 1770 => to_unsigned(293, 10), 1771 => to_unsigned(60, 10), 1772 => to_unsigned(720, 10), 1773 => to_unsigned(866, 10), 1774 => to_unsigned(235, 10), 1775 => to_unsigned(284, 10), 1776 => to_unsigned(908, 10), 1777 => to_unsigned(770, 10), 1778 => to_unsigned(302, 10), 1779 => to_unsigned(106, 10), 1780 => to_unsigned(429, 10), 1781 => to_unsigned(266, 10), 1782 => to_unsigned(420, 10), 1783 => to_unsigned(72, 10), 1784 => to_unsigned(435, 10), 1785 => to_unsigned(954, 10), 1786 => to_unsigned(499, 10), 1787 => to_unsigned(1023, 10), 1788 => to_unsigned(887, 10), 1789 => to_unsigned(784, 10), 1790 => to_unsigned(382, 10), 1791 => to_unsigned(816, 10), 1792 => to_unsigned(792, 10), 1793 => to_unsigned(729, 10), 1794 => to_unsigned(228, 10), 1795 => to_unsigned(127, 10), 1796 => to_unsigned(733, 10), 1797 => to_unsigned(768, 10), 1798 => to_unsigned(957, 10), 1799 => to_unsigned(992, 10), 1800 => to_unsigned(170, 10), 1801 => to_unsigned(899, 10), 1802 => to_unsigned(944, 10), 1803 => to_unsigned(936, 10), 1804 => to_unsigned(1000, 10), 1805 => to_unsigned(753, 10), 1806 => to_unsigned(414, 10), 1807 => to_unsigned(425, 10), 1808 => to_unsigned(761, 10), 1809 => to_unsigned(667, 10), 1810 => to_unsigned(458, 10), 1811 => to_unsigned(569, 10), 1812 => to_unsigned(703, 10), 1813 => to_unsigned(201, 10), 1814 => to_unsigned(930, 10), 1815 => to_unsigned(553, 10), 1816 => to_unsigned(152, 10), 1817 => to_unsigned(1018, 10), 1818 => to_unsigned(400, 10), 1819 => to_unsigned(263, 10), 1820 => to_unsigned(304, 10), 1821 => to_unsigned(754, 10), 1822 => to_unsigned(290, 10), 1823 => to_unsigned(335, 10), 1824 => to_unsigned(68, 10), 1825 => to_unsigned(890, 10), 1826 => to_unsigned(870, 10), 1827 => to_unsigned(680, 10), 1828 => to_unsigned(135, 10), 1829 => to_unsigned(426, 10), 1830 => to_unsigned(291, 10), 1831 => to_unsigned(756, 10), 1832 => to_unsigned(971, 10), 1833 => to_unsigned(716, 10), 1834 => to_unsigned(224, 10), 1835 => to_unsigned(883, 10), 1836 => to_unsigned(747, 10), 1837 => to_unsigned(455, 10), 1838 => to_unsigned(680, 10), 1839 => to_unsigned(232, 10), 1840 => to_unsigned(45, 10), 1841 => to_unsigned(207, 10), 1842 => to_unsigned(593, 10), 1843 => to_unsigned(458, 10), 1844 => to_unsigned(378, 10), 1845 => to_unsigned(731, 10), 1846 => to_unsigned(112, 10), 1847 => to_unsigned(146, 10), 1848 => to_unsigned(758, 10), 1849 => to_unsigned(113, 10), 1850 => to_unsigned(374, 10), 1851 => to_unsigned(423, 10), 1852 => to_unsigned(705, 10), 1853 => to_unsigned(911, 10), 1854 => to_unsigned(749, 10), 1855 => to_unsigned(252, 10), 1856 => to_unsigned(501, 10), 1857 => to_unsigned(954, 10), 1858 => to_unsigned(471, 10), 1859 => to_unsigned(582, 10), 1860 => to_unsigned(950, 10), 1861 => to_unsigned(669, 10), 1862 => to_unsigned(205, 10), 1863 => to_unsigned(863, 10), 1864 => to_unsigned(325, 10), 1865 => to_unsigned(78, 10), 1866 => to_unsigned(731, 10), 1867 => to_unsigned(673, 10), 1868 => to_unsigned(797, 10), 1869 => to_unsigned(379, 10), 1870 => to_unsigned(538, 10), 1871 => to_unsigned(547, 10), 1872 => to_unsigned(120, 10), 1873 => to_unsigned(1012, 10), 1874 => to_unsigned(280, 10), 1875 => to_unsigned(699, 10), 1876 => to_unsigned(869, 10), 1877 => to_unsigned(902, 10), 1878 => to_unsigned(766, 10), 1879 => to_unsigned(322, 10), 1880 => to_unsigned(36, 10), 1881 => to_unsigned(497, 10), 1882 => to_unsigned(699, 10), 1883 => to_unsigned(956, 10), 1884 => to_unsigned(750, 10), 1885 => to_unsigned(823, 10), 1886 => to_unsigned(164, 10), 1887 => to_unsigned(271, 10), 1888 => to_unsigned(797, 10), 1889 => to_unsigned(732, 10), 1890 => to_unsigned(422, 10), 1891 => to_unsigned(132, 10), 1892 => to_unsigned(472, 10), 1893 => to_unsigned(893, 10), 1894 => to_unsigned(429, 10), 1895 => to_unsigned(996, 10), 1896 => to_unsigned(257, 10), 1897 => to_unsigned(859, 10), 1898 => to_unsigned(454, 10), 1899 => to_unsigned(672, 10), 1900 => to_unsigned(659, 10), 1901 => to_unsigned(870, 10), 1902 => to_unsigned(545, 10), 1903 => to_unsigned(375, 10), 1904 => to_unsigned(813, 10), 1905 => to_unsigned(880, 10), 1906 => to_unsigned(900, 10), 1907 => to_unsigned(1010, 10), 1908 => to_unsigned(195, 10), 1909 => to_unsigned(770, 10), 1910 => to_unsigned(814, 10), 1911 => to_unsigned(881, 10), 1912 => to_unsigned(505, 10), 1913 => to_unsigned(298, 10), 1914 => to_unsigned(706, 10), 1915 => to_unsigned(892, 10), 1916 => to_unsigned(545, 10), 1917 => to_unsigned(713, 10), 1918 => to_unsigned(654, 10), 1919 => to_unsigned(849, 10), 1920 => to_unsigned(45, 10), 1921 => to_unsigned(973, 10), 1922 => to_unsigned(146, 10), 1923 => to_unsigned(804, 10), 1924 => to_unsigned(378, 10), 1925 => to_unsigned(402, 10), 1926 => to_unsigned(885, 10), 1927 => to_unsigned(470, 10), 1928 => to_unsigned(911, 10), 1929 => to_unsigned(823, 10), 1930 => to_unsigned(630, 10), 1931 => to_unsigned(462, 10), 1932 => to_unsigned(989, 10), 1933 => to_unsigned(636, 10), 1934 => to_unsigned(615, 10), 1935 => to_unsigned(395, 10), 1936 => to_unsigned(83, 10), 1937 => to_unsigned(989, 10), 1938 => to_unsigned(305, 10), 1939 => to_unsigned(828, 10), 1940 => to_unsigned(104, 10), 1941 => to_unsigned(644, 10), 1942 => to_unsigned(923, 10), 1943 => to_unsigned(888, 10), 1944 => to_unsigned(609, 10), 1945 => to_unsigned(346, 10), 1946 => to_unsigned(432, 10), 1947 => to_unsigned(500, 10), 1948 => to_unsigned(718, 10), 1949 => to_unsigned(774, 10), 1950 => to_unsigned(369, 10), 1951 => to_unsigned(322, 10), 1952 => to_unsigned(264, 10), 1953 => to_unsigned(128, 10), 1954 => to_unsigned(44, 10), 1955 => to_unsigned(1008, 10), 1956 => to_unsigned(319, 10), 1957 => to_unsigned(268, 10), 1958 => to_unsigned(915, 10), 1959 => to_unsigned(951, 10), 1960 => to_unsigned(759, 10), 1961 => to_unsigned(107, 10), 1962 => to_unsigned(0, 10), 1963 => to_unsigned(339, 10), 1964 => to_unsigned(389, 10), 1965 => to_unsigned(736, 10), 1966 => to_unsigned(320, 10), 1967 => to_unsigned(186, 10), 1968 => to_unsigned(286, 10), 1969 => to_unsigned(959, 10), 1970 => to_unsigned(723, 10), 1971 => to_unsigned(99, 10), 1972 => to_unsigned(635, 10), 1973 => to_unsigned(887, 10), 1974 => to_unsigned(376, 10), 1975 => to_unsigned(155, 10), 1976 => to_unsigned(205, 10), 1977 => to_unsigned(401, 10), 1978 => to_unsigned(933, 10), 1979 => to_unsigned(177, 10), 1980 => to_unsigned(708, 10), 1981 => to_unsigned(221, 10), 1982 => to_unsigned(529, 10), 1983 => to_unsigned(224, 10), 1984 => to_unsigned(683, 10), 1985 => to_unsigned(851, 10), 1986 => to_unsigned(744, 10), 1987 => to_unsigned(228, 10), 1988 => to_unsigned(491, 10), 1989 => to_unsigned(466, 10), 1990 => to_unsigned(71, 10), 1991 => to_unsigned(486, 10), 1992 => to_unsigned(594, 10), 1993 => to_unsigned(641, 10), 1994 => to_unsigned(830, 10), 1995 => to_unsigned(50, 10), 1996 => to_unsigned(908, 10), 1997 => to_unsigned(898, 10), 1998 => to_unsigned(370, 10), 1999 => to_unsigned(735, 10), 2000 => to_unsigned(86, 10), 2001 => to_unsigned(817, 10), 2002 => to_unsigned(905, 10), 2003 => to_unsigned(942, 10), 2004 => to_unsigned(1012, 10), 2005 => to_unsigned(886, 10), 2006 => to_unsigned(1007, 10), 2007 => to_unsigned(35, 10), 2008 => to_unsigned(218, 10), 2009 => to_unsigned(880, 10), 2010 => to_unsigned(166, 10), 2011 => to_unsigned(230, 10), 2012 => to_unsigned(190, 10), 2013 => to_unsigned(755, 10), 2014 => to_unsigned(298, 10), 2015 => to_unsigned(49, 10), 2016 => to_unsigned(646, 10), 2017 => to_unsigned(888, 10), 2018 => to_unsigned(720, 10), 2019 => to_unsigned(133, 10), 2020 => to_unsigned(57, 10), 2021 => to_unsigned(976, 10), 2022 => to_unsigned(156, 10), 2023 => to_unsigned(328, 10), 2024 => to_unsigned(38, 10), 2025 => to_unsigned(383, 10), 2026 => to_unsigned(591, 10), 2027 => to_unsigned(937, 10), 2028 => to_unsigned(57, 10), 2029 => to_unsigned(247, 10), 2030 => to_unsigned(427, 10), 2031 => to_unsigned(471, 10), 2032 => to_unsigned(924, 10), 2033 => to_unsigned(685, 10), 2034 => to_unsigned(4, 10), 2035 => to_unsigned(720, 10), 2036 => to_unsigned(582, 10), 2037 => to_unsigned(982, 10), 2038 => to_unsigned(475, 10), 2039 => to_unsigned(689, 10), 2040 => to_unsigned(503, 10), 2041 => to_unsigned(815, 10), 2042 => to_unsigned(877, 10), 2043 => to_unsigned(499, 10), 2044 => to_unsigned(748, 10), 2045 => to_unsigned(310, 10), 2046 => to_unsigned(33, 10), 2047 => to_unsigned(127, 10)),
            2 => (0 => to_unsigned(154, 10), 1 => to_unsigned(322, 10), 2 => to_unsigned(505, 10), 3 => to_unsigned(495, 10), 4 => to_unsigned(781, 10), 5 => to_unsigned(703, 10), 6 => to_unsigned(331, 10), 7 => to_unsigned(910, 10), 8 => to_unsigned(764, 10), 9 => to_unsigned(10, 10), 10 => to_unsigned(329, 10), 11 => to_unsigned(409, 10), 12 => to_unsigned(650, 10), 13 => to_unsigned(922, 10), 14 => to_unsigned(764, 10), 15 => to_unsigned(890, 10), 16 => to_unsigned(273, 10), 17 => to_unsigned(341, 10), 18 => to_unsigned(163, 10), 19 => to_unsigned(930, 10), 20 => to_unsigned(928, 10), 21 => to_unsigned(189, 10), 22 => to_unsigned(954, 10), 23 => to_unsigned(448, 10), 24 => to_unsigned(580, 10), 25 => to_unsigned(783, 10), 26 => to_unsigned(617, 10), 27 => to_unsigned(793, 10), 28 => to_unsigned(508, 10), 29 => to_unsigned(316, 10), 30 => to_unsigned(524, 10), 31 => to_unsigned(50, 10), 32 => to_unsigned(835, 10), 33 => to_unsigned(920, 10), 34 => to_unsigned(761, 10), 35 => to_unsigned(579, 10), 36 => to_unsigned(205, 10), 37 => to_unsigned(53, 10), 38 => to_unsigned(902, 10), 39 => to_unsigned(549, 10), 40 => to_unsigned(967, 10), 41 => to_unsigned(199, 10), 42 => to_unsigned(183, 10), 43 => to_unsigned(63, 10), 44 => to_unsigned(817, 10), 45 => to_unsigned(473, 10), 46 => to_unsigned(9, 10), 47 => to_unsigned(441, 10), 48 => to_unsigned(455, 10), 49 => to_unsigned(714, 10), 50 => to_unsigned(166, 10), 51 => to_unsigned(975, 10), 52 => to_unsigned(466, 10), 53 => to_unsigned(597, 10), 54 => to_unsigned(546, 10), 55 => to_unsigned(931, 10), 56 => to_unsigned(81, 10), 57 => to_unsigned(319, 10), 58 => to_unsigned(155, 10), 59 => to_unsigned(599, 10), 60 => to_unsigned(163, 10), 61 => to_unsigned(469, 10), 62 => to_unsigned(745, 10), 63 => to_unsigned(289, 10), 64 => to_unsigned(160, 10), 65 => to_unsigned(848, 10), 66 => to_unsigned(359, 10), 67 => to_unsigned(86, 10), 68 => to_unsigned(75, 10), 69 => to_unsigned(535, 10), 70 => to_unsigned(603, 10), 71 => to_unsigned(838, 10), 72 => to_unsigned(389, 10), 73 => to_unsigned(232, 10), 74 => to_unsigned(886, 10), 75 => to_unsigned(206, 10), 76 => to_unsigned(525, 10), 77 => to_unsigned(305, 10), 78 => to_unsigned(829, 10), 79 => to_unsigned(1007, 10), 80 => to_unsigned(352, 10), 81 => to_unsigned(641, 10), 82 => to_unsigned(356, 10), 83 => to_unsigned(34, 10), 84 => to_unsigned(699, 10), 85 => to_unsigned(122, 10), 86 => to_unsigned(512, 10), 87 => to_unsigned(545, 10), 88 => to_unsigned(266, 10), 89 => to_unsigned(257, 10), 90 => to_unsigned(587, 10), 91 => to_unsigned(431, 10), 92 => to_unsigned(241, 10), 93 => to_unsigned(510, 10), 94 => to_unsigned(699, 10), 95 => to_unsigned(610, 10), 96 => to_unsigned(706, 10), 97 => to_unsigned(684, 10), 98 => to_unsigned(842, 10), 99 => to_unsigned(676, 10), 100 => to_unsigned(62, 10), 101 => to_unsigned(273, 10), 102 => to_unsigned(761, 10), 103 => to_unsigned(233, 10), 104 => to_unsigned(570, 10), 105 => to_unsigned(136, 10), 106 => to_unsigned(896, 10), 107 => to_unsigned(124, 10), 108 => to_unsigned(290, 10), 109 => to_unsigned(724, 10), 110 => to_unsigned(423, 10), 111 => to_unsigned(521, 10), 112 => to_unsigned(674, 10), 113 => to_unsigned(603, 10), 114 => to_unsigned(242, 10), 115 => to_unsigned(4, 10), 116 => to_unsigned(962, 10), 117 => to_unsigned(779, 10), 118 => to_unsigned(765, 10), 119 => to_unsigned(886, 10), 120 => to_unsigned(16, 10), 121 => to_unsigned(718, 10), 122 => to_unsigned(430, 10), 123 => to_unsigned(889, 10), 124 => to_unsigned(290, 10), 125 => to_unsigned(238, 10), 126 => to_unsigned(213, 10), 127 => to_unsigned(777, 10), 128 => to_unsigned(919, 10), 129 => to_unsigned(174, 10), 130 => to_unsigned(30, 10), 131 => to_unsigned(728, 10), 132 => to_unsigned(959, 10), 133 => to_unsigned(129, 10), 134 => to_unsigned(480, 10), 135 => to_unsigned(969, 10), 136 => to_unsigned(193, 10), 137 => to_unsigned(67, 10), 138 => to_unsigned(198, 10), 139 => to_unsigned(502, 10), 140 => to_unsigned(984, 10), 141 => to_unsigned(444, 10), 142 => to_unsigned(771, 10), 143 => to_unsigned(181, 10), 144 => to_unsigned(193, 10), 145 => to_unsigned(470, 10), 146 => to_unsigned(883, 10), 147 => to_unsigned(769, 10), 148 => to_unsigned(256, 10), 149 => to_unsigned(694, 10), 150 => to_unsigned(230, 10), 151 => to_unsigned(76, 10), 152 => to_unsigned(323, 10), 153 => to_unsigned(140, 10), 154 => to_unsigned(439, 10), 155 => to_unsigned(102, 10), 156 => to_unsigned(165, 10), 157 => to_unsigned(782, 10), 158 => to_unsigned(173, 10), 159 => to_unsigned(421, 10), 160 => to_unsigned(951, 10), 161 => to_unsigned(337, 10), 162 => to_unsigned(306, 10), 163 => to_unsigned(870, 10), 164 => to_unsigned(551, 10), 165 => to_unsigned(72, 10), 166 => to_unsigned(173, 10), 167 => to_unsigned(608, 10), 168 => to_unsigned(280, 10), 169 => to_unsigned(161, 10), 170 => to_unsigned(245, 10), 171 => to_unsigned(309, 10), 172 => to_unsigned(443, 10), 173 => to_unsigned(927, 10), 174 => to_unsigned(385, 10), 175 => to_unsigned(861, 10), 176 => to_unsigned(420, 10), 177 => to_unsigned(305, 10), 178 => to_unsigned(446, 10), 179 => to_unsigned(755, 10), 180 => to_unsigned(866, 10), 181 => to_unsigned(746, 10), 182 => to_unsigned(127, 10), 183 => to_unsigned(37, 10), 184 => to_unsigned(186, 10), 185 => to_unsigned(625, 10), 186 => to_unsigned(621, 10), 187 => to_unsigned(644, 10), 188 => to_unsigned(480, 10), 189 => to_unsigned(899, 10), 190 => to_unsigned(382, 10), 191 => to_unsigned(739, 10), 192 => to_unsigned(910, 10), 193 => to_unsigned(1004, 10), 194 => to_unsigned(701, 10), 195 => to_unsigned(113, 10), 196 => to_unsigned(132, 10), 197 => to_unsigned(262, 10), 198 => to_unsigned(243, 10), 199 => to_unsigned(748, 10), 200 => to_unsigned(766, 10), 201 => to_unsigned(547, 10), 202 => to_unsigned(119, 10), 203 => to_unsigned(565, 10), 204 => to_unsigned(636, 10), 205 => to_unsigned(923, 10), 206 => to_unsigned(61, 10), 207 => to_unsigned(301, 10), 208 => to_unsigned(264, 10), 209 => to_unsigned(961, 10), 210 => to_unsigned(555, 10), 211 => to_unsigned(875, 10), 212 => to_unsigned(959, 10), 213 => to_unsigned(32, 10), 214 => to_unsigned(23, 10), 215 => to_unsigned(1000, 10), 216 => to_unsigned(665, 10), 217 => to_unsigned(509, 10), 218 => to_unsigned(369, 10), 219 => to_unsigned(1006, 10), 220 => to_unsigned(578, 10), 221 => to_unsigned(501, 10), 222 => to_unsigned(1016, 10), 223 => to_unsigned(35, 10), 224 => to_unsigned(860, 10), 225 => to_unsigned(715, 10), 226 => to_unsigned(562, 10), 227 => to_unsigned(177, 10), 228 => to_unsigned(577, 10), 229 => to_unsigned(549, 10), 230 => to_unsigned(540, 10), 231 => to_unsigned(901, 10), 232 => to_unsigned(62, 10), 233 => to_unsigned(865, 10), 234 => to_unsigned(561, 10), 235 => to_unsigned(858, 10), 236 => to_unsigned(520, 10), 237 => to_unsigned(294, 10), 238 => to_unsigned(40, 10), 239 => to_unsigned(780, 10), 240 => to_unsigned(1022, 10), 241 => to_unsigned(463, 10), 242 => to_unsigned(175, 10), 243 => to_unsigned(470, 10), 244 => to_unsigned(10, 10), 245 => to_unsigned(119, 10), 246 => to_unsigned(547, 10), 247 => to_unsigned(275, 10), 248 => to_unsigned(674, 10), 249 => to_unsigned(952, 10), 250 => to_unsigned(265, 10), 251 => to_unsigned(89, 10), 252 => to_unsigned(638, 10), 253 => to_unsigned(692, 10), 254 => to_unsigned(454, 10), 255 => to_unsigned(935, 10), 256 => to_unsigned(75, 10), 257 => to_unsigned(140, 10), 258 => to_unsigned(994, 10), 259 => to_unsigned(416, 10), 260 => to_unsigned(565, 10), 261 => to_unsigned(122, 10), 262 => to_unsigned(592, 10), 263 => to_unsigned(963, 10), 264 => to_unsigned(78, 10), 265 => to_unsigned(228, 10), 266 => to_unsigned(55, 10), 267 => to_unsigned(209, 10), 268 => to_unsigned(713, 10), 269 => to_unsigned(61, 10), 270 => to_unsigned(930, 10), 271 => to_unsigned(155, 10), 272 => to_unsigned(156, 10), 273 => to_unsigned(685, 10), 274 => to_unsigned(522, 10), 275 => to_unsigned(517, 10), 276 => to_unsigned(735, 10), 277 => to_unsigned(719, 10), 278 => to_unsigned(556, 10), 279 => to_unsigned(589, 10), 280 => to_unsigned(183, 10), 281 => to_unsigned(198, 10), 282 => to_unsigned(911, 10), 283 => to_unsigned(7, 10), 284 => to_unsigned(108, 10), 285 => to_unsigned(850, 10), 286 => to_unsigned(293, 10), 287 => to_unsigned(793, 10), 288 => to_unsigned(571, 10), 289 => to_unsigned(284, 10), 290 => to_unsigned(818, 10), 291 => to_unsigned(346, 10), 292 => to_unsigned(200, 10), 293 => to_unsigned(303, 10), 294 => to_unsigned(187, 10), 295 => to_unsigned(413, 10), 296 => to_unsigned(147, 10), 297 => to_unsigned(547, 10), 298 => to_unsigned(370, 10), 299 => to_unsigned(57, 10), 300 => to_unsigned(419, 10), 301 => to_unsigned(925, 10), 302 => to_unsigned(336, 10), 303 => to_unsigned(452, 10), 304 => to_unsigned(739, 10), 305 => to_unsigned(50, 10), 306 => to_unsigned(688, 10), 307 => to_unsigned(703, 10), 308 => to_unsigned(164, 10), 309 => to_unsigned(597, 10), 310 => to_unsigned(771, 10), 311 => to_unsigned(265, 10), 312 => to_unsigned(418, 10), 313 => to_unsigned(50, 10), 314 => to_unsigned(975, 10), 315 => to_unsigned(933, 10), 316 => to_unsigned(908, 10), 317 => to_unsigned(458, 10), 318 => to_unsigned(532, 10), 319 => to_unsigned(721, 10), 320 => to_unsigned(980, 10), 321 => to_unsigned(406, 10), 322 => to_unsigned(527, 10), 323 => to_unsigned(995, 10), 324 => to_unsigned(858, 10), 325 => to_unsigned(770, 10), 326 => to_unsigned(787, 10), 327 => to_unsigned(336, 10), 328 => to_unsigned(894, 10), 329 => to_unsigned(563, 10), 330 => to_unsigned(740, 10), 331 => to_unsigned(334, 10), 332 => to_unsigned(102, 10), 333 => to_unsigned(562, 10), 334 => to_unsigned(727, 10), 335 => to_unsigned(187, 10), 336 => to_unsigned(939, 10), 337 => to_unsigned(900, 10), 338 => to_unsigned(818, 10), 339 => to_unsigned(906, 10), 340 => to_unsigned(108, 10), 341 => to_unsigned(30, 10), 342 => to_unsigned(800, 10), 343 => to_unsigned(164, 10), 344 => to_unsigned(402, 10), 345 => to_unsigned(535, 10), 346 => to_unsigned(90, 10), 347 => to_unsigned(229, 10), 348 => to_unsigned(687, 10), 349 => to_unsigned(803, 10), 350 => to_unsigned(560, 10), 351 => to_unsigned(639, 10), 352 => to_unsigned(812, 10), 353 => to_unsigned(61, 10), 354 => to_unsigned(95, 10), 355 => to_unsigned(282, 10), 356 => to_unsigned(997, 10), 357 => to_unsigned(884, 10), 358 => to_unsigned(430, 10), 359 => to_unsigned(545, 10), 360 => to_unsigned(382, 10), 361 => to_unsigned(568, 10), 362 => to_unsigned(888, 10), 363 => to_unsigned(997, 10), 364 => to_unsigned(199, 10), 365 => to_unsigned(936, 10), 366 => to_unsigned(786, 10), 367 => to_unsigned(233, 10), 368 => to_unsigned(671, 10), 369 => to_unsigned(126, 10), 370 => to_unsigned(636, 10), 371 => to_unsigned(831, 10), 372 => to_unsigned(286, 10), 373 => to_unsigned(74, 10), 374 => to_unsigned(925, 10), 375 => to_unsigned(723, 10), 376 => to_unsigned(421, 10), 377 => to_unsigned(913, 10), 378 => to_unsigned(9, 10), 379 => to_unsigned(398, 10), 380 => to_unsigned(647, 10), 381 => to_unsigned(635, 10), 382 => to_unsigned(654, 10), 383 => to_unsigned(433, 10), 384 => to_unsigned(923, 10), 385 => to_unsigned(155, 10), 386 => to_unsigned(544, 10), 387 => to_unsigned(434, 10), 388 => to_unsigned(737, 10), 389 => to_unsigned(480, 10), 390 => to_unsigned(886, 10), 391 => to_unsigned(487, 10), 392 => to_unsigned(503, 10), 393 => to_unsigned(608, 10), 394 => to_unsigned(855, 10), 395 => to_unsigned(453, 10), 396 => to_unsigned(81, 10), 397 => to_unsigned(633, 10), 398 => to_unsigned(995, 10), 399 => to_unsigned(996, 10), 400 => to_unsigned(896, 10), 401 => to_unsigned(796, 10), 402 => to_unsigned(428, 10), 403 => to_unsigned(65, 10), 404 => to_unsigned(240, 10), 405 => to_unsigned(688, 10), 406 => to_unsigned(702, 10), 407 => to_unsigned(580, 10), 408 => to_unsigned(125, 10), 409 => to_unsigned(548, 10), 410 => to_unsigned(894, 10), 411 => to_unsigned(222, 10), 412 => to_unsigned(640, 10), 413 => to_unsigned(565, 10), 414 => to_unsigned(754, 10), 415 => to_unsigned(298, 10), 416 => to_unsigned(789, 10), 417 => to_unsigned(914, 10), 418 => to_unsigned(811, 10), 419 => to_unsigned(502, 10), 420 => to_unsigned(609, 10), 421 => to_unsigned(128, 10), 422 => to_unsigned(126, 10), 423 => to_unsigned(686, 10), 424 => to_unsigned(455, 10), 425 => to_unsigned(556, 10), 426 => to_unsigned(1015, 10), 427 => to_unsigned(590, 10), 428 => to_unsigned(930, 10), 429 => to_unsigned(88, 10), 430 => to_unsigned(499, 10), 431 => to_unsigned(318, 10), 432 => to_unsigned(67, 10), 433 => to_unsigned(191, 10), 434 => to_unsigned(963, 10), 435 => to_unsigned(490, 10), 436 => to_unsigned(267, 10), 437 => to_unsigned(874, 10), 438 => to_unsigned(40, 10), 439 => to_unsigned(617, 10), 440 => to_unsigned(291, 10), 441 => to_unsigned(66, 10), 442 => to_unsigned(740, 10), 443 => to_unsigned(461, 10), 444 => to_unsigned(909, 10), 445 => to_unsigned(737, 10), 446 => to_unsigned(174, 10), 447 => to_unsigned(834, 10), 448 => to_unsigned(476, 10), 449 => to_unsigned(428, 10), 450 => to_unsigned(16, 10), 451 => to_unsigned(505, 10), 452 => to_unsigned(801, 10), 453 => to_unsigned(48, 10), 454 => to_unsigned(696, 10), 455 => to_unsigned(83, 10), 456 => to_unsigned(54, 10), 457 => to_unsigned(195, 10), 458 => to_unsigned(598, 10), 459 => to_unsigned(852, 10), 460 => to_unsigned(838, 10), 461 => to_unsigned(268, 10), 462 => to_unsigned(307, 10), 463 => to_unsigned(164, 10), 464 => to_unsigned(985, 10), 465 => to_unsigned(552, 10), 466 => to_unsigned(70, 10), 467 => to_unsigned(881, 10), 468 => to_unsigned(536, 10), 469 => to_unsigned(439, 10), 470 => to_unsigned(809, 10), 471 => to_unsigned(955, 10), 472 => to_unsigned(1013, 10), 473 => to_unsigned(902, 10), 474 => to_unsigned(302, 10), 475 => to_unsigned(376, 10), 476 => to_unsigned(614, 10), 477 => to_unsigned(577, 10), 478 => to_unsigned(477, 10), 479 => to_unsigned(964, 10), 480 => to_unsigned(281, 10), 481 => to_unsigned(936, 10), 482 => to_unsigned(795, 10), 483 => to_unsigned(336, 10), 484 => to_unsigned(715, 10), 485 => to_unsigned(465, 10), 486 => to_unsigned(882, 10), 487 => to_unsigned(880, 10), 488 => to_unsigned(56, 10), 489 => to_unsigned(462, 10), 490 => to_unsigned(184, 10), 491 => to_unsigned(230, 10), 492 => to_unsigned(529, 10), 493 => to_unsigned(361, 10), 494 => to_unsigned(751, 10), 495 => to_unsigned(170, 10), 496 => to_unsigned(544, 10), 497 => to_unsigned(845, 10), 498 => to_unsigned(119, 10), 499 => to_unsigned(8, 10), 500 => to_unsigned(926, 10), 501 => to_unsigned(1017, 10), 502 => to_unsigned(80, 10), 503 => to_unsigned(577, 10), 504 => to_unsigned(691, 10), 505 => to_unsigned(94, 10), 506 => to_unsigned(384, 10), 507 => to_unsigned(582, 10), 508 => to_unsigned(948, 10), 509 => to_unsigned(84, 10), 510 => to_unsigned(939, 10), 511 => to_unsigned(856, 10), 512 => to_unsigned(101, 10), 513 => to_unsigned(363, 10), 514 => to_unsigned(867, 10), 515 => to_unsigned(694, 10), 516 => to_unsigned(402, 10), 517 => to_unsigned(926, 10), 518 => to_unsigned(390, 10), 519 => to_unsigned(737, 10), 520 => to_unsigned(86, 10), 521 => to_unsigned(831, 10), 522 => to_unsigned(755, 10), 523 => to_unsigned(988, 10), 524 => to_unsigned(216, 10), 525 => to_unsigned(788, 10), 526 => to_unsigned(669, 10), 527 => to_unsigned(258, 10), 528 => to_unsigned(505, 10), 529 => to_unsigned(598, 10), 530 => to_unsigned(321, 10), 531 => to_unsigned(755, 10), 532 => to_unsigned(836, 10), 533 => to_unsigned(247, 10), 534 => to_unsigned(887, 10), 535 => to_unsigned(314, 10), 536 => to_unsigned(892, 10), 537 => to_unsigned(173, 10), 538 => to_unsigned(308, 10), 539 => to_unsigned(439, 10), 540 => to_unsigned(388, 10), 541 => to_unsigned(597, 10), 542 => to_unsigned(634, 10), 543 => to_unsigned(742, 10), 544 => to_unsigned(300, 10), 545 => to_unsigned(433, 10), 546 => to_unsigned(817, 10), 547 => to_unsigned(695, 10), 548 => to_unsigned(975, 10), 549 => to_unsigned(127, 10), 550 => to_unsigned(904, 10), 551 => to_unsigned(156, 10), 552 => to_unsigned(580, 10), 553 => to_unsigned(673, 10), 554 => to_unsigned(628, 10), 555 => to_unsigned(36, 10), 556 => to_unsigned(626, 10), 557 => to_unsigned(66, 10), 558 => to_unsigned(750, 10), 559 => to_unsigned(732, 10), 560 => to_unsigned(49, 10), 561 => to_unsigned(559, 10), 562 => to_unsigned(191, 10), 563 => to_unsigned(832, 10), 564 => to_unsigned(414, 10), 565 => to_unsigned(883, 10), 566 => to_unsigned(901, 10), 567 => to_unsigned(273, 10), 568 => to_unsigned(149, 10), 569 => to_unsigned(96, 10), 570 => to_unsigned(229, 10), 571 => to_unsigned(579, 10), 572 => to_unsigned(816, 10), 573 => to_unsigned(635, 10), 574 => to_unsigned(966, 10), 575 => to_unsigned(537, 10), 576 => to_unsigned(814, 10), 577 => to_unsigned(123, 10), 578 => to_unsigned(1012, 10), 579 => to_unsigned(558, 10), 580 => to_unsigned(901, 10), 581 => to_unsigned(612, 10), 582 => to_unsigned(39, 10), 583 => to_unsigned(245, 10), 584 => to_unsigned(320, 10), 585 => to_unsigned(29, 10), 586 => to_unsigned(56, 10), 587 => to_unsigned(209, 10), 588 => to_unsigned(458, 10), 589 => to_unsigned(895, 10), 590 => to_unsigned(893, 10), 591 => to_unsigned(145, 10), 592 => to_unsigned(642, 10), 593 => to_unsigned(26, 10), 594 => to_unsigned(307, 10), 595 => to_unsigned(428, 10), 596 => to_unsigned(873, 10), 597 => to_unsigned(196, 10), 598 => to_unsigned(344, 10), 599 => to_unsigned(717, 10), 600 => to_unsigned(362, 10), 601 => to_unsigned(771, 10), 602 => to_unsigned(738, 10), 603 => to_unsigned(644, 10), 604 => to_unsigned(430, 10), 605 => to_unsigned(715, 10), 606 => to_unsigned(58, 10), 607 => to_unsigned(726, 10), 608 => to_unsigned(648, 10), 609 => to_unsigned(470, 10), 610 => to_unsigned(398, 10), 611 => to_unsigned(748, 10), 612 => to_unsigned(141, 10), 613 => to_unsigned(649, 10), 614 => to_unsigned(849, 10), 615 => to_unsigned(306, 10), 616 => to_unsigned(8, 10), 617 => to_unsigned(624, 10), 618 => to_unsigned(89, 10), 619 => to_unsigned(329, 10), 620 => to_unsigned(494, 10), 621 => to_unsigned(416, 10), 622 => to_unsigned(161, 10), 623 => to_unsigned(859, 10), 624 => to_unsigned(421, 10), 625 => to_unsigned(807, 10), 626 => to_unsigned(658, 10), 627 => to_unsigned(900, 10), 628 => to_unsigned(693, 10), 629 => to_unsigned(646, 10), 630 => to_unsigned(15, 10), 631 => to_unsigned(944, 10), 632 => to_unsigned(138, 10), 633 => to_unsigned(628, 10), 634 => to_unsigned(58, 10), 635 => to_unsigned(132, 10), 636 => to_unsigned(583, 10), 637 => to_unsigned(51, 10), 638 => to_unsigned(225, 10), 639 => to_unsigned(409, 10), 640 => to_unsigned(701, 10), 641 => to_unsigned(679, 10), 642 => to_unsigned(302, 10), 643 => to_unsigned(118, 10), 644 => to_unsigned(1014, 10), 645 => to_unsigned(133, 10), 646 => to_unsigned(998, 10), 647 => to_unsigned(584, 10), 648 => to_unsigned(660, 10), 649 => to_unsigned(67, 10), 650 => to_unsigned(116, 10), 651 => to_unsigned(97, 10), 652 => to_unsigned(944, 10), 653 => to_unsigned(409, 10), 654 => to_unsigned(347, 10), 655 => to_unsigned(398, 10), 656 => to_unsigned(154, 10), 657 => to_unsigned(612, 10), 658 => to_unsigned(252, 10), 659 => to_unsigned(824, 10), 660 => to_unsigned(616, 10), 661 => to_unsigned(131, 10), 662 => to_unsigned(1006, 10), 663 => to_unsigned(815, 10), 664 => to_unsigned(297, 10), 665 => to_unsigned(676, 10), 666 => to_unsigned(527, 10), 667 => to_unsigned(264, 10), 668 => to_unsigned(607, 10), 669 => to_unsigned(170, 10), 670 => to_unsigned(182, 10), 671 => to_unsigned(27, 10), 672 => to_unsigned(976, 10), 673 => to_unsigned(559, 10), 674 => to_unsigned(175, 10), 675 => to_unsigned(507, 10), 676 => to_unsigned(848, 10), 677 => to_unsigned(922, 10), 678 => to_unsigned(82, 10), 679 => to_unsigned(470, 10), 680 => to_unsigned(0, 10), 681 => to_unsigned(441, 10), 682 => to_unsigned(990, 10), 683 => to_unsigned(452, 10), 684 => to_unsigned(84, 10), 685 => to_unsigned(991, 10), 686 => to_unsigned(555, 10), 687 => to_unsigned(572, 10), 688 => to_unsigned(811, 10), 689 => to_unsigned(202, 10), 690 => to_unsigned(801, 10), 691 => to_unsigned(174, 10), 692 => to_unsigned(147, 10), 693 => to_unsigned(684, 10), 694 => to_unsigned(513, 10), 695 => to_unsigned(523, 10), 696 => to_unsigned(309, 10), 697 => to_unsigned(337, 10), 698 => to_unsigned(775, 10), 699 => to_unsigned(121, 10), 700 => to_unsigned(884, 10), 701 => to_unsigned(5, 10), 702 => to_unsigned(610, 10), 703 => to_unsigned(141, 10), 704 => to_unsigned(117, 10), 705 => to_unsigned(728, 10), 706 => to_unsigned(185, 10), 707 => to_unsigned(352, 10), 708 => to_unsigned(126, 10), 709 => to_unsigned(137, 10), 710 => to_unsigned(204, 10), 711 => to_unsigned(180, 10), 712 => to_unsigned(843, 10), 713 => to_unsigned(125, 10), 714 => to_unsigned(9, 10), 715 => to_unsigned(760, 10), 716 => to_unsigned(919, 10), 717 => to_unsigned(854, 10), 718 => to_unsigned(274, 10), 719 => to_unsigned(898, 10), 720 => to_unsigned(133, 10), 721 => to_unsigned(753, 10), 722 => to_unsigned(144, 10), 723 => to_unsigned(273, 10), 724 => to_unsigned(911, 10), 725 => to_unsigned(146, 10), 726 => to_unsigned(51, 10), 727 => to_unsigned(359, 10), 728 => to_unsigned(362, 10), 729 => to_unsigned(82, 10), 730 => to_unsigned(118, 10), 731 => to_unsigned(266, 10), 732 => to_unsigned(108, 10), 733 => to_unsigned(861, 10), 734 => to_unsigned(615, 10), 735 => to_unsigned(859, 10), 736 => to_unsigned(147, 10), 737 => to_unsigned(721, 10), 738 => to_unsigned(648, 10), 739 => to_unsigned(303, 10), 740 => to_unsigned(897, 10), 741 => to_unsigned(89, 10), 742 => to_unsigned(545, 10), 743 => to_unsigned(26, 10), 744 => to_unsigned(325, 10), 745 => to_unsigned(765, 10), 746 => to_unsigned(776, 10), 747 => to_unsigned(663, 10), 748 => to_unsigned(873, 10), 749 => to_unsigned(87, 10), 750 => to_unsigned(631, 10), 751 => to_unsigned(485, 10), 752 => to_unsigned(272, 10), 753 => to_unsigned(599, 10), 754 => to_unsigned(194, 10), 755 => to_unsigned(707, 10), 756 => to_unsigned(639, 10), 757 => to_unsigned(95, 10), 758 => to_unsigned(10, 10), 759 => to_unsigned(681, 10), 760 => to_unsigned(831, 10), 761 => to_unsigned(117, 10), 762 => to_unsigned(790, 10), 763 => to_unsigned(98, 10), 764 => to_unsigned(823, 10), 765 => to_unsigned(511, 10), 766 => to_unsigned(581, 10), 767 => to_unsigned(562, 10), 768 => to_unsigned(101, 10), 769 => to_unsigned(210, 10), 770 => to_unsigned(372, 10), 771 => to_unsigned(594, 10), 772 => to_unsigned(22, 10), 773 => to_unsigned(320, 10), 774 => to_unsigned(723, 10), 775 => to_unsigned(727, 10), 776 => to_unsigned(594, 10), 777 => to_unsigned(922, 10), 778 => to_unsigned(270, 10), 779 => to_unsigned(888, 10), 780 => to_unsigned(520, 10), 781 => to_unsigned(98, 10), 782 => to_unsigned(941, 10), 783 => to_unsigned(929, 10), 784 => to_unsigned(299, 10), 785 => to_unsigned(80, 10), 786 => to_unsigned(953, 10), 787 => to_unsigned(9, 10), 788 => to_unsigned(257, 10), 789 => to_unsigned(623, 10), 790 => to_unsigned(96, 10), 791 => to_unsigned(300, 10), 792 => to_unsigned(744, 10), 793 => to_unsigned(981, 10), 794 => to_unsigned(713, 10), 795 => to_unsigned(1014, 10), 796 => to_unsigned(576, 10), 797 => to_unsigned(705, 10), 798 => to_unsigned(128, 10), 799 => to_unsigned(272, 10), 800 => to_unsigned(42, 10), 801 => to_unsigned(373, 10), 802 => to_unsigned(222, 10), 803 => to_unsigned(862, 10), 804 => to_unsigned(304, 10), 805 => to_unsigned(302, 10), 806 => to_unsigned(1000, 10), 807 => to_unsigned(60, 10), 808 => to_unsigned(946, 10), 809 => to_unsigned(136, 10), 810 => to_unsigned(680, 10), 811 => to_unsigned(454, 10), 812 => to_unsigned(315, 10), 813 => to_unsigned(213, 10), 814 => to_unsigned(266, 10), 815 => to_unsigned(311, 10), 816 => to_unsigned(388, 10), 817 => to_unsigned(915, 10), 818 => to_unsigned(134, 10), 819 => to_unsigned(113, 10), 820 => to_unsigned(876, 10), 821 => to_unsigned(325, 10), 822 => to_unsigned(353, 10), 823 => to_unsigned(746, 10), 824 => to_unsigned(45, 10), 825 => to_unsigned(4, 10), 826 => to_unsigned(745, 10), 827 => to_unsigned(515, 10), 828 => to_unsigned(73, 10), 829 => to_unsigned(898, 10), 830 => to_unsigned(361, 10), 831 => to_unsigned(651, 10), 832 => to_unsigned(972, 10), 833 => to_unsigned(454, 10), 834 => to_unsigned(754, 10), 835 => to_unsigned(114, 10), 836 => to_unsigned(900, 10), 837 => to_unsigned(296, 10), 838 => to_unsigned(525, 10), 839 => to_unsigned(825, 10), 840 => to_unsigned(74, 10), 841 => to_unsigned(458, 10), 842 => to_unsigned(458, 10), 843 => to_unsigned(524, 10), 844 => to_unsigned(325, 10), 845 => to_unsigned(464, 10), 846 => to_unsigned(555, 10), 847 => to_unsigned(595, 10), 848 => to_unsigned(530, 10), 849 => to_unsigned(326, 10), 850 => to_unsigned(379, 10), 851 => to_unsigned(90, 10), 852 => to_unsigned(1006, 10), 853 => to_unsigned(518, 10), 854 => to_unsigned(2, 10), 855 => to_unsigned(541, 10), 856 => to_unsigned(450, 10), 857 => to_unsigned(181, 10), 858 => to_unsigned(386, 10), 859 => to_unsigned(274, 10), 860 => to_unsigned(919, 10), 861 => to_unsigned(263, 10), 862 => to_unsigned(659, 10), 863 => to_unsigned(357, 10), 864 => to_unsigned(988, 10), 865 => to_unsigned(1009, 10), 866 => to_unsigned(709, 10), 867 => to_unsigned(244, 10), 868 => to_unsigned(635, 10), 869 => to_unsigned(197, 10), 870 => to_unsigned(50, 10), 871 => to_unsigned(313, 10), 872 => to_unsigned(483, 10), 873 => to_unsigned(364, 10), 874 => to_unsigned(287, 10), 875 => to_unsigned(643, 10), 876 => to_unsigned(785, 10), 877 => to_unsigned(686, 10), 878 => to_unsigned(713, 10), 879 => to_unsigned(905, 10), 880 => to_unsigned(837, 10), 881 => to_unsigned(162, 10), 882 => to_unsigned(1021, 10), 883 => to_unsigned(615, 10), 884 => to_unsigned(800, 10), 885 => to_unsigned(863, 10), 886 => to_unsigned(873, 10), 887 => to_unsigned(736, 10), 888 => to_unsigned(153, 10), 889 => to_unsigned(467, 10), 890 => to_unsigned(159, 10), 891 => to_unsigned(691, 10), 892 => to_unsigned(647, 10), 893 => to_unsigned(308, 10), 894 => to_unsigned(982, 10), 895 => to_unsigned(655, 10), 896 => to_unsigned(178, 10), 897 => to_unsigned(944, 10), 898 => to_unsigned(548, 10), 899 => to_unsigned(858, 10), 900 => to_unsigned(294, 10), 901 => to_unsigned(230, 10), 902 => to_unsigned(738, 10), 903 => to_unsigned(152, 10), 904 => to_unsigned(617, 10), 905 => to_unsigned(606, 10), 906 => to_unsigned(769, 10), 907 => to_unsigned(41, 10), 908 => to_unsigned(759, 10), 909 => to_unsigned(504, 10), 910 => to_unsigned(216, 10), 911 => to_unsigned(347, 10), 912 => to_unsigned(171, 10), 913 => to_unsigned(656, 10), 914 => to_unsigned(972, 10), 915 => to_unsigned(73, 10), 916 => to_unsigned(193, 10), 917 => to_unsigned(843, 10), 918 => to_unsigned(686, 10), 919 => to_unsigned(122, 10), 920 => to_unsigned(904, 10), 921 => to_unsigned(530, 10), 922 => to_unsigned(784, 10), 923 => to_unsigned(552, 10), 924 => to_unsigned(874, 10), 925 => to_unsigned(242, 10), 926 => to_unsigned(857, 10), 927 => to_unsigned(136, 10), 928 => to_unsigned(622, 10), 929 => to_unsigned(758, 10), 930 => to_unsigned(218, 10), 931 => to_unsigned(898, 10), 932 => to_unsigned(280, 10), 933 => to_unsigned(318, 10), 934 => to_unsigned(587, 10), 935 => to_unsigned(232, 10), 936 => to_unsigned(710, 10), 937 => to_unsigned(317, 10), 938 => to_unsigned(749, 10), 939 => to_unsigned(514, 10), 940 => to_unsigned(209, 10), 941 => to_unsigned(512, 10), 942 => to_unsigned(661, 10), 943 => to_unsigned(416, 10), 944 => to_unsigned(954, 10), 945 => to_unsigned(236, 10), 946 => to_unsigned(540, 10), 947 => to_unsigned(332, 10), 948 => to_unsigned(187, 10), 949 => to_unsigned(637, 10), 950 => to_unsigned(156, 10), 951 => to_unsigned(229, 10), 952 => to_unsigned(123, 10), 953 => to_unsigned(510, 10), 954 => to_unsigned(983, 10), 955 => to_unsigned(818, 10), 956 => to_unsigned(89, 10), 957 => to_unsigned(438, 10), 958 => to_unsigned(747, 10), 959 => to_unsigned(655, 10), 960 => to_unsigned(204, 10), 961 => to_unsigned(877, 10), 962 => to_unsigned(616, 10), 963 => to_unsigned(719, 10), 964 => to_unsigned(602, 10), 965 => to_unsigned(423, 10), 966 => to_unsigned(132, 10), 967 => to_unsigned(178, 10), 968 => to_unsigned(897, 10), 969 => to_unsigned(495, 10), 970 => to_unsigned(927, 10), 971 => to_unsigned(509, 10), 972 => to_unsigned(112, 10), 973 => to_unsigned(753, 10), 974 => to_unsigned(441, 10), 975 => to_unsigned(639, 10), 976 => to_unsigned(900, 10), 977 => to_unsigned(622, 10), 978 => to_unsigned(213, 10), 979 => to_unsigned(77, 10), 980 => to_unsigned(539, 10), 981 => to_unsigned(324, 10), 982 => to_unsigned(324, 10), 983 => to_unsigned(940, 10), 984 => to_unsigned(125, 10), 985 => to_unsigned(774, 10), 986 => to_unsigned(415, 10), 987 => to_unsigned(634, 10), 988 => to_unsigned(250, 10), 989 => to_unsigned(504, 10), 990 => to_unsigned(260, 10), 991 => to_unsigned(559, 10), 992 => to_unsigned(456, 10), 993 => to_unsigned(544, 10), 994 => to_unsigned(233, 10), 995 => to_unsigned(749, 10), 996 => to_unsigned(520, 10), 997 => to_unsigned(884, 10), 998 => to_unsigned(538, 10), 999 => to_unsigned(958, 10), 1000 => to_unsigned(396, 10), 1001 => to_unsigned(460, 10), 1002 => to_unsigned(439, 10), 1003 => to_unsigned(805, 10), 1004 => to_unsigned(970, 10), 1005 => to_unsigned(263, 10), 1006 => to_unsigned(851, 10), 1007 => to_unsigned(23, 10), 1008 => to_unsigned(256, 10), 1009 => to_unsigned(1004, 10), 1010 => to_unsigned(241, 10), 1011 => to_unsigned(466, 10), 1012 => to_unsigned(612, 10), 1013 => to_unsigned(866, 10), 1014 => to_unsigned(501, 10), 1015 => to_unsigned(385, 10), 1016 => to_unsigned(383, 10), 1017 => to_unsigned(216, 10), 1018 => to_unsigned(1012, 10), 1019 => to_unsigned(680, 10), 1020 => to_unsigned(620, 10), 1021 => to_unsigned(871, 10), 1022 => to_unsigned(407, 10), 1023 => to_unsigned(419, 10), 1024 => to_unsigned(800, 10), 1025 => to_unsigned(702, 10), 1026 => to_unsigned(724, 10), 1027 => to_unsigned(40, 10), 1028 => to_unsigned(861, 10), 1029 => to_unsigned(344, 10), 1030 => to_unsigned(557, 10), 1031 => to_unsigned(197, 10), 1032 => to_unsigned(279, 10), 1033 => to_unsigned(848, 10), 1034 => to_unsigned(362, 10), 1035 => to_unsigned(963, 10), 1036 => to_unsigned(1016, 10), 1037 => to_unsigned(758, 10), 1038 => to_unsigned(653, 10), 1039 => to_unsigned(768, 10), 1040 => to_unsigned(1007, 10), 1041 => to_unsigned(801, 10), 1042 => to_unsigned(699, 10), 1043 => to_unsigned(306, 10), 1044 => to_unsigned(13, 10), 1045 => to_unsigned(712, 10), 1046 => to_unsigned(146, 10), 1047 => to_unsigned(429, 10), 1048 => to_unsigned(708, 10), 1049 => to_unsigned(1010, 10), 1050 => to_unsigned(288, 10), 1051 => to_unsigned(632, 10), 1052 => to_unsigned(733, 10), 1053 => to_unsigned(973, 10), 1054 => to_unsigned(824, 10), 1055 => to_unsigned(717, 10), 1056 => to_unsigned(1016, 10), 1057 => to_unsigned(389, 10), 1058 => to_unsigned(195, 10), 1059 => to_unsigned(856, 10), 1060 => to_unsigned(953, 10), 1061 => to_unsigned(606, 10), 1062 => to_unsigned(453, 10), 1063 => to_unsigned(975, 10), 1064 => to_unsigned(149, 10), 1065 => to_unsigned(504, 10), 1066 => to_unsigned(539, 10), 1067 => to_unsigned(717, 10), 1068 => to_unsigned(27, 10), 1069 => to_unsigned(877, 10), 1070 => to_unsigned(631, 10), 1071 => to_unsigned(604, 10), 1072 => to_unsigned(844, 10), 1073 => to_unsigned(47, 10), 1074 => to_unsigned(677, 10), 1075 => to_unsigned(772, 10), 1076 => to_unsigned(195, 10), 1077 => to_unsigned(1003, 10), 1078 => to_unsigned(858, 10), 1079 => to_unsigned(399, 10), 1080 => to_unsigned(926, 10), 1081 => to_unsigned(949, 10), 1082 => to_unsigned(45, 10), 1083 => to_unsigned(55, 10), 1084 => to_unsigned(642, 10), 1085 => to_unsigned(238, 10), 1086 => to_unsigned(118, 10), 1087 => to_unsigned(664, 10), 1088 => to_unsigned(850, 10), 1089 => to_unsigned(152, 10), 1090 => to_unsigned(404, 10), 1091 => to_unsigned(218, 10), 1092 => to_unsigned(735, 10), 1093 => to_unsigned(75, 10), 1094 => to_unsigned(745, 10), 1095 => to_unsigned(902, 10), 1096 => to_unsigned(1012, 10), 1097 => to_unsigned(202, 10), 1098 => to_unsigned(56, 10), 1099 => to_unsigned(892, 10), 1100 => to_unsigned(688, 10), 1101 => to_unsigned(47, 10), 1102 => to_unsigned(70, 10), 1103 => to_unsigned(437, 10), 1104 => to_unsigned(167, 10), 1105 => to_unsigned(606, 10), 1106 => to_unsigned(486, 10), 1107 => to_unsigned(596, 10), 1108 => to_unsigned(560, 10), 1109 => to_unsigned(645, 10), 1110 => to_unsigned(33, 10), 1111 => to_unsigned(794, 10), 1112 => to_unsigned(732, 10), 1113 => to_unsigned(691, 10), 1114 => to_unsigned(633, 10), 1115 => to_unsigned(206, 10), 1116 => to_unsigned(121, 10), 1117 => to_unsigned(912, 10), 1118 => to_unsigned(621, 10), 1119 => to_unsigned(211, 10), 1120 => to_unsigned(331, 10), 1121 => to_unsigned(525, 10), 1122 => to_unsigned(57, 10), 1123 => to_unsigned(437, 10), 1124 => to_unsigned(805, 10), 1125 => to_unsigned(285, 10), 1126 => to_unsigned(747, 10), 1127 => to_unsigned(168, 10), 1128 => to_unsigned(671, 10), 1129 => to_unsigned(475, 10), 1130 => to_unsigned(347, 10), 1131 => to_unsigned(770, 10), 1132 => to_unsigned(213, 10), 1133 => to_unsigned(766, 10), 1134 => to_unsigned(447, 10), 1135 => to_unsigned(982, 10), 1136 => to_unsigned(510, 10), 1137 => to_unsigned(733, 10), 1138 => to_unsigned(364, 10), 1139 => to_unsigned(38, 10), 1140 => to_unsigned(430, 10), 1141 => to_unsigned(920, 10), 1142 => to_unsigned(332, 10), 1143 => to_unsigned(605, 10), 1144 => to_unsigned(401, 10), 1145 => to_unsigned(460, 10), 1146 => to_unsigned(196, 10), 1147 => to_unsigned(777, 10), 1148 => to_unsigned(914, 10), 1149 => to_unsigned(806, 10), 1150 => to_unsigned(985, 10), 1151 => to_unsigned(591, 10), 1152 => to_unsigned(600, 10), 1153 => to_unsigned(1015, 10), 1154 => to_unsigned(723, 10), 1155 => to_unsigned(663, 10), 1156 => to_unsigned(873, 10), 1157 => to_unsigned(828, 10), 1158 => to_unsigned(52, 10), 1159 => to_unsigned(274, 10), 1160 => to_unsigned(838, 10), 1161 => to_unsigned(328, 10), 1162 => to_unsigned(650, 10), 1163 => to_unsigned(792, 10), 1164 => to_unsigned(749, 10), 1165 => to_unsigned(684, 10), 1166 => to_unsigned(491, 10), 1167 => to_unsigned(769, 10), 1168 => to_unsigned(723, 10), 1169 => to_unsigned(114, 10), 1170 => to_unsigned(178, 10), 1171 => to_unsigned(294, 10), 1172 => to_unsigned(155, 10), 1173 => to_unsigned(659, 10), 1174 => to_unsigned(323, 10), 1175 => to_unsigned(378, 10), 1176 => to_unsigned(72, 10), 1177 => to_unsigned(598, 10), 1178 => to_unsigned(186, 10), 1179 => to_unsigned(574, 10), 1180 => to_unsigned(524, 10), 1181 => to_unsigned(704, 10), 1182 => to_unsigned(784, 10), 1183 => to_unsigned(792, 10), 1184 => to_unsigned(370, 10), 1185 => to_unsigned(351, 10), 1186 => to_unsigned(480, 10), 1187 => to_unsigned(99, 10), 1188 => to_unsigned(581, 10), 1189 => to_unsigned(885, 10), 1190 => to_unsigned(54, 10), 1191 => to_unsigned(122, 10), 1192 => to_unsigned(197, 10), 1193 => to_unsigned(317, 10), 1194 => to_unsigned(641, 10), 1195 => to_unsigned(536, 10), 1196 => to_unsigned(780, 10), 1197 => to_unsigned(945, 10), 1198 => to_unsigned(937, 10), 1199 => to_unsigned(694, 10), 1200 => to_unsigned(339, 10), 1201 => to_unsigned(182, 10), 1202 => to_unsigned(415, 10), 1203 => to_unsigned(490, 10), 1204 => to_unsigned(967, 10), 1205 => to_unsigned(788, 10), 1206 => to_unsigned(538, 10), 1207 => to_unsigned(541, 10), 1208 => to_unsigned(307, 10), 1209 => to_unsigned(461, 10), 1210 => to_unsigned(83, 10), 1211 => to_unsigned(978, 10), 1212 => to_unsigned(64, 10), 1213 => to_unsigned(1001, 10), 1214 => to_unsigned(609, 10), 1215 => to_unsigned(932, 10), 1216 => to_unsigned(218, 10), 1217 => to_unsigned(253, 10), 1218 => to_unsigned(538, 10), 1219 => to_unsigned(254, 10), 1220 => to_unsigned(485, 10), 1221 => to_unsigned(139, 10), 1222 => to_unsigned(123, 10), 1223 => to_unsigned(136, 10), 1224 => to_unsigned(122, 10), 1225 => to_unsigned(602, 10), 1226 => to_unsigned(29, 10), 1227 => to_unsigned(237, 10), 1228 => to_unsigned(191, 10), 1229 => to_unsigned(700, 10), 1230 => to_unsigned(791, 10), 1231 => to_unsigned(978, 10), 1232 => to_unsigned(880, 10), 1233 => to_unsigned(150, 10), 1234 => to_unsigned(867, 10), 1235 => to_unsigned(103, 10), 1236 => to_unsigned(171, 10), 1237 => to_unsigned(401, 10), 1238 => to_unsigned(62, 10), 1239 => to_unsigned(344, 10), 1240 => to_unsigned(660, 10), 1241 => to_unsigned(918, 10), 1242 => to_unsigned(585, 10), 1243 => to_unsigned(810, 10), 1244 => to_unsigned(853, 10), 1245 => to_unsigned(125, 10), 1246 => to_unsigned(573, 10), 1247 => to_unsigned(77, 10), 1248 => to_unsigned(943, 10), 1249 => to_unsigned(1005, 10), 1250 => to_unsigned(625, 10), 1251 => to_unsigned(126, 10), 1252 => to_unsigned(901, 10), 1253 => to_unsigned(669, 10), 1254 => to_unsigned(683, 10), 1255 => to_unsigned(65, 10), 1256 => to_unsigned(475, 10), 1257 => to_unsigned(323, 10), 1258 => to_unsigned(793, 10), 1259 => to_unsigned(144, 10), 1260 => to_unsigned(592, 10), 1261 => to_unsigned(236, 10), 1262 => to_unsigned(687, 10), 1263 => to_unsigned(446, 10), 1264 => to_unsigned(11, 10), 1265 => to_unsigned(584, 10), 1266 => to_unsigned(30, 10), 1267 => to_unsigned(495, 10), 1268 => to_unsigned(174, 10), 1269 => to_unsigned(788, 10), 1270 => to_unsigned(587, 10), 1271 => to_unsigned(796, 10), 1272 => to_unsigned(274, 10), 1273 => to_unsigned(708, 10), 1274 => to_unsigned(70, 10), 1275 => to_unsigned(277, 10), 1276 => to_unsigned(363, 10), 1277 => to_unsigned(888, 10), 1278 => to_unsigned(133, 10), 1279 => to_unsigned(1, 10), 1280 => to_unsigned(862, 10), 1281 => to_unsigned(843, 10), 1282 => to_unsigned(93, 10), 1283 => to_unsigned(875, 10), 1284 => to_unsigned(256, 10), 1285 => to_unsigned(748, 10), 1286 => to_unsigned(402, 10), 1287 => to_unsigned(449, 10), 1288 => to_unsigned(212, 10), 1289 => to_unsigned(185, 10), 1290 => to_unsigned(499, 10), 1291 => to_unsigned(95, 10), 1292 => to_unsigned(115, 10), 1293 => to_unsigned(550, 10), 1294 => to_unsigned(91, 10), 1295 => to_unsigned(237, 10), 1296 => to_unsigned(270, 10), 1297 => to_unsigned(925, 10), 1298 => to_unsigned(124, 10), 1299 => to_unsigned(734, 10), 1300 => to_unsigned(257, 10), 1301 => to_unsigned(571, 10), 1302 => to_unsigned(134, 10), 1303 => to_unsigned(333, 10), 1304 => to_unsigned(37, 10), 1305 => to_unsigned(546, 10), 1306 => to_unsigned(794, 10), 1307 => to_unsigned(180, 10), 1308 => to_unsigned(259, 10), 1309 => to_unsigned(417, 10), 1310 => to_unsigned(725, 10), 1311 => to_unsigned(744, 10), 1312 => to_unsigned(958, 10), 1313 => to_unsigned(886, 10), 1314 => to_unsigned(664, 10), 1315 => to_unsigned(40, 10), 1316 => to_unsigned(894, 10), 1317 => to_unsigned(583, 10), 1318 => to_unsigned(167, 10), 1319 => to_unsigned(617, 10), 1320 => to_unsigned(249, 10), 1321 => to_unsigned(66, 10), 1322 => to_unsigned(682, 10), 1323 => to_unsigned(775, 10), 1324 => to_unsigned(992, 10), 1325 => to_unsigned(191, 10), 1326 => to_unsigned(969, 10), 1327 => to_unsigned(411, 10), 1328 => to_unsigned(908, 10), 1329 => to_unsigned(1021, 10), 1330 => to_unsigned(897, 10), 1331 => to_unsigned(145, 10), 1332 => to_unsigned(669, 10), 1333 => to_unsigned(722, 10), 1334 => to_unsigned(641, 10), 1335 => to_unsigned(826, 10), 1336 => to_unsigned(100, 10), 1337 => to_unsigned(71, 10), 1338 => to_unsigned(758, 10), 1339 => to_unsigned(447, 10), 1340 => to_unsigned(470, 10), 1341 => to_unsigned(887, 10), 1342 => to_unsigned(955, 10), 1343 => to_unsigned(1022, 10), 1344 => to_unsigned(235, 10), 1345 => to_unsigned(533, 10), 1346 => to_unsigned(812, 10), 1347 => to_unsigned(595, 10), 1348 => to_unsigned(996, 10), 1349 => to_unsigned(292, 10), 1350 => to_unsigned(182, 10), 1351 => to_unsigned(158, 10), 1352 => to_unsigned(98, 10), 1353 => to_unsigned(895, 10), 1354 => to_unsigned(1009, 10), 1355 => to_unsigned(572, 10), 1356 => to_unsigned(123, 10), 1357 => to_unsigned(42, 10), 1358 => to_unsigned(606, 10), 1359 => to_unsigned(50, 10), 1360 => to_unsigned(189, 10), 1361 => to_unsigned(328, 10), 1362 => to_unsigned(603, 10), 1363 => to_unsigned(747, 10), 1364 => to_unsigned(964, 10), 1365 => to_unsigned(167, 10), 1366 => to_unsigned(819, 10), 1367 => to_unsigned(298, 10), 1368 => to_unsigned(626, 10), 1369 => to_unsigned(845, 10), 1370 => to_unsigned(36, 10), 1371 => to_unsigned(490, 10), 1372 => to_unsigned(301, 10), 1373 => to_unsigned(747, 10), 1374 => to_unsigned(712, 10), 1375 => to_unsigned(779, 10), 1376 => to_unsigned(785, 10), 1377 => to_unsigned(975, 10), 1378 => to_unsigned(274, 10), 1379 => to_unsigned(448, 10), 1380 => to_unsigned(1015, 10), 1381 => to_unsigned(182, 10), 1382 => to_unsigned(180, 10), 1383 => to_unsigned(209, 10), 1384 => to_unsigned(105, 10), 1385 => to_unsigned(938, 10), 1386 => to_unsigned(855, 10), 1387 => to_unsigned(926, 10), 1388 => to_unsigned(537, 10), 1389 => to_unsigned(829, 10), 1390 => to_unsigned(517, 10), 1391 => to_unsigned(399, 10), 1392 => to_unsigned(873, 10), 1393 => to_unsigned(405, 10), 1394 => to_unsigned(912, 10), 1395 => to_unsigned(786, 10), 1396 => to_unsigned(777, 10), 1397 => to_unsigned(547, 10), 1398 => to_unsigned(41, 10), 1399 => to_unsigned(850, 10), 1400 => to_unsigned(579, 10), 1401 => to_unsigned(578, 10), 1402 => to_unsigned(143, 10), 1403 => to_unsigned(656, 10), 1404 => to_unsigned(138, 10), 1405 => to_unsigned(1001, 10), 1406 => to_unsigned(804, 10), 1407 => to_unsigned(112, 10), 1408 => to_unsigned(195, 10), 1409 => to_unsigned(723, 10), 1410 => to_unsigned(997, 10), 1411 => to_unsigned(793, 10), 1412 => to_unsigned(560, 10), 1413 => to_unsigned(666, 10), 1414 => to_unsigned(905, 10), 1415 => to_unsigned(470, 10), 1416 => to_unsigned(794, 10), 1417 => to_unsigned(121, 10), 1418 => to_unsigned(0, 10), 1419 => to_unsigned(961, 10), 1420 => to_unsigned(465, 10), 1421 => to_unsigned(372, 10), 1422 => to_unsigned(81, 10), 1423 => to_unsigned(111, 10), 1424 => to_unsigned(495, 10), 1425 => to_unsigned(950, 10), 1426 => to_unsigned(624, 10), 1427 => to_unsigned(447, 10), 1428 => to_unsigned(446, 10), 1429 => to_unsigned(54, 10), 1430 => to_unsigned(7, 10), 1431 => to_unsigned(155, 10), 1432 => to_unsigned(250, 10), 1433 => to_unsigned(488, 10), 1434 => to_unsigned(286, 10), 1435 => to_unsigned(99, 10), 1436 => to_unsigned(418, 10), 1437 => to_unsigned(558, 10), 1438 => to_unsigned(803, 10), 1439 => to_unsigned(81, 10), 1440 => to_unsigned(471, 10), 1441 => to_unsigned(1006, 10), 1442 => to_unsigned(820, 10), 1443 => to_unsigned(222, 10), 1444 => to_unsigned(788, 10), 1445 => to_unsigned(1022, 10), 1446 => to_unsigned(82, 10), 1447 => to_unsigned(964, 10), 1448 => to_unsigned(628, 10), 1449 => to_unsigned(292, 10), 1450 => to_unsigned(901, 10), 1451 => to_unsigned(580, 10), 1452 => to_unsigned(320, 10), 1453 => to_unsigned(881, 10), 1454 => to_unsigned(315, 10), 1455 => to_unsigned(799, 10), 1456 => to_unsigned(56, 10), 1457 => to_unsigned(595, 10), 1458 => to_unsigned(848, 10), 1459 => to_unsigned(616, 10), 1460 => to_unsigned(784, 10), 1461 => to_unsigned(909, 10), 1462 => to_unsigned(423, 10), 1463 => to_unsigned(372, 10), 1464 => to_unsigned(495, 10), 1465 => to_unsigned(251, 10), 1466 => to_unsigned(771, 10), 1467 => to_unsigned(484, 10), 1468 => to_unsigned(25, 10), 1469 => to_unsigned(214, 10), 1470 => to_unsigned(797, 10), 1471 => to_unsigned(963, 10), 1472 => to_unsigned(449, 10), 1473 => to_unsigned(798, 10), 1474 => to_unsigned(598, 10), 1475 => to_unsigned(34, 10), 1476 => to_unsigned(744, 10), 1477 => to_unsigned(875, 10), 1478 => to_unsigned(916, 10), 1479 => to_unsigned(493, 10), 1480 => to_unsigned(780, 10), 1481 => to_unsigned(600, 10), 1482 => to_unsigned(2, 10), 1483 => to_unsigned(683, 10), 1484 => to_unsigned(474, 10), 1485 => to_unsigned(540, 10), 1486 => to_unsigned(702, 10), 1487 => to_unsigned(943, 10), 1488 => to_unsigned(228, 10), 1489 => to_unsigned(428, 10), 1490 => to_unsigned(138, 10), 1491 => to_unsigned(707, 10), 1492 => to_unsigned(155, 10), 1493 => to_unsigned(206, 10), 1494 => to_unsigned(78, 10), 1495 => to_unsigned(803, 10), 1496 => to_unsigned(927, 10), 1497 => to_unsigned(171, 10), 1498 => to_unsigned(32, 10), 1499 => to_unsigned(85, 10), 1500 => to_unsigned(935, 10), 1501 => to_unsigned(276, 10), 1502 => to_unsigned(225, 10), 1503 => to_unsigned(751, 10), 1504 => to_unsigned(536, 10), 1505 => to_unsigned(805, 10), 1506 => to_unsigned(774, 10), 1507 => to_unsigned(37, 10), 1508 => to_unsigned(51, 10), 1509 => to_unsigned(62, 10), 1510 => to_unsigned(820, 10), 1511 => to_unsigned(924, 10), 1512 => to_unsigned(554, 10), 1513 => to_unsigned(997, 10), 1514 => to_unsigned(868, 10), 1515 => to_unsigned(193, 10), 1516 => to_unsigned(938, 10), 1517 => to_unsigned(668, 10), 1518 => to_unsigned(185, 10), 1519 => to_unsigned(428, 10), 1520 => to_unsigned(265, 10), 1521 => to_unsigned(86, 10), 1522 => to_unsigned(609, 10), 1523 => to_unsigned(264, 10), 1524 => to_unsigned(207, 10), 1525 => to_unsigned(929, 10), 1526 => to_unsigned(888, 10), 1527 => to_unsigned(121, 10), 1528 => to_unsigned(26, 10), 1529 => to_unsigned(497, 10), 1530 => to_unsigned(124, 10), 1531 => to_unsigned(680, 10), 1532 => to_unsigned(126, 10), 1533 => to_unsigned(283, 10), 1534 => to_unsigned(84, 10), 1535 => to_unsigned(484, 10), 1536 => to_unsigned(855, 10), 1537 => to_unsigned(847, 10), 1538 => to_unsigned(723, 10), 1539 => to_unsigned(899, 10), 1540 => to_unsigned(130, 10), 1541 => to_unsigned(53, 10), 1542 => to_unsigned(1000, 10), 1543 => to_unsigned(274, 10), 1544 => to_unsigned(425, 10), 1545 => to_unsigned(692, 10), 1546 => to_unsigned(839, 10), 1547 => to_unsigned(506, 10), 1548 => to_unsigned(163, 10), 1549 => to_unsigned(634, 10), 1550 => to_unsigned(717, 10), 1551 => to_unsigned(602, 10), 1552 => to_unsigned(554, 10), 1553 => to_unsigned(335, 10), 1554 => to_unsigned(850, 10), 1555 => to_unsigned(221, 10), 1556 => to_unsigned(109, 10), 1557 => to_unsigned(834, 10), 1558 => to_unsigned(355, 10), 1559 => to_unsigned(895, 10), 1560 => to_unsigned(29, 10), 1561 => to_unsigned(910, 10), 1562 => to_unsigned(49, 10), 1563 => to_unsigned(998, 10), 1564 => to_unsigned(676, 10), 1565 => to_unsigned(43, 10), 1566 => to_unsigned(333, 10), 1567 => to_unsigned(524, 10), 1568 => to_unsigned(286, 10), 1569 => to_unsigned(304, 10), 1570 => to_unsigned(990, 10), 1571 => to_unsigned(210, 10), 1572 => to_unsigned(220, 10), 1573 => to_unsigned(396, 10), 1574 => to_unsigned(380, 10), 1575 => to_unsigned(972, 10), 1576 => to_unsigned(684, 10), 1577 => to_unsigned(773, 10), 1578 => to_unsigned(1017, 10), 1579 => to_unsigned(843, 10), 1580 => to_unsigned(889, 10), 1581 => to_unsigned(136, 10), 1582 => to_unsigned(815, 10), 1583 => to_unsigned(168, 10), 1584 => to_unsigned(715, 10), 1585 => to_unsigned(367, 10), 1586 => to_unsigned(438, 10), 1587 => to_unsigned(849, 10), 1588 => to_unsigned(539, 10), 1589 => to_unsigned(389, 10), 1590 => to_unsigned(696, 10), 1591 => to_unsigned(914, 10), 1592 => to_unsigned(315, 10), 1593 => to_unsigned(588, 10), 1594 => to_unsigned(767, 10), 1595 => to_unsigned(944, 10), 1596 => to_unsigned(688, 10), 1597 => to_unsigned(178, 10), 1598 => to_unsigned(431, 10), 1599 => to_unsigned(706, 10), 1600 => to_unsigned(783, 10), 1601 => to_unsigned(456, 10), 1602 => to_unsigned(585, 10), 1603 => to_unsigned(228, 10), 1604 => to_unsigned(233, 10), 1605 => to_unsigned(239, 10), 1606 => to_unsigned(60, 10), 1607 => to_unsigned(255, 10), 1608 => to_unsigned(13, 10), 1609 => to_unsigned(556, 10), 1610 => to_unsigned(176, 10), 1611 => to_unsigned(94, 10), 1612 => to_unsigned(528, 10), 1613 => to_unsigned(408, 10), 1614 => to_unsigned(288, 10), 1615 => to_unsigned(282, 10), 1616 => to_unsigned(516, 10), 1617 => to_unsigned(885, 10), 1618 => to_unsigned(495, 10), 1619 => to_unsigned(968, 10), 1620 => to_unsigned(716, 10), 1621 => to_unsigned(246, 10), 1622 => to_unsigned(940, 10), 1623 => to_unsigned(268, 10), 1624 => to_unsigned(249, 10), 1625 => to_unsigned(540, 10), 1626 => to_unsigned(5, 10), 1627 => to_unsigned(379, 10), 1628 => to_unsigned(268, 10), 1629 => to_unsigned(593, 10), 1630 => to_unsigned(936, 10), 1631 => to_unsigned(497, 10), 1632 => to_unsigned(317, 10), 1633 => to_unsigned(992, 10), 1634 => to_unsigned(834, 10), 1635 => to_unsigned(912, 10), 1636 => to_unsigned(661, 10), 1637 => to_unsigned(856, 10), 1638 => to_unsigned(749, 10), 1639 => to_unsigned(512, 10), 1640 => to_unsigned(590, 10), 1641 => to_unsigned(571, 10), 1642 => to_unsigned(448, 10), 1643 => to_unsigned(612, 10), 1644 => to_unsigned(746, 10), 1645 => to_unsigned(629, 10), 1646 => to_unsigned(711, 10), 1647 => to_unsigned(630, 10), 1648 => to_unsigned(411, 10), 1649 => to_unsigned(945, 10), 1650 => to_unsigned(642, 10), 1651 => to_unsigned(622, 10), 1652 => to_unsigned(180, 10), 1653 => to_unsigned(807, 10), 1654 => to_unsigned(0, 10), 1655 => to_unsigned(737, 10), 1656 => to_unsigned(684, 10), 1657 => to_unsigned(177, 10), 1658 => to_unsigned(658, 10), 1659 => to_unsigned(539, 10), 1660 => to_unsigned(164, 10), 1661 => to_unsigned(514, 10), 1662 => to_unsigned(74, 10), 1663 => to_unsigned(450, 10), 1664 => to_unsigned(913, 10), 1665 => to_unsigned(101, 10), 1666 => to_unsigned(675, 10), 1667 => to_unsigned(268, 10), 1668 => to_unsigned(499, 10), 1669 => to_unsigned(95, 10), 1670 => to_unsigned(415, 10), 1671 => to_unsigned(564, 10), 1672 => to_unsigned(717, 10), 1673 => to_unsigned(333, 10), 1674 => to_unsigned(614, 10), 1675 => to_unsigned(279, 10), 1676 => to_unsigned(336, 10), 1677 => to_unsigned(989, 10), 1678 => to_unsigned(776, 10), 1679 => to_unsigned(726, 10), 1680 => to_unsigned(340, 10), 1681 => to_unsigned(777, 10), 1682 => to_unsigned(969, 10), 1683 => to_unsigned(771, 10), 1684 => to_unsigned(359, 10), 1685 => to_unsigned(31, 10), 1686 => to_unsigned(858, 10), 1687 => to_unsigned(928, 10), 1688 => to_unsigned(647, 10), 1689 => to_unsigned(809, 10), 1690 => to_unsigned(644, 10), 1691 => to_unsigned(877, 10), 1692 => to_unsigned(114, 10), 1693 => to_unsigned(398, 10), 1694 => to_unsigned(783, 10), 1695 => to_unsigned(1002, 10), 1696 => to_unsigned(717, 10), 1697 => to_unsigned(63, 10), 1698 => to_unsigned(182, 10), 1699 => to_unsigned(664, 10), 1700 => to_unsigned(657, 10), 1701 => to_unsigned(364, 10), 1702 => to_unsigned(645, 10), 1703 => to_unsigned(756, 10), 1704 => to_unsigned(1005, 10), 1705 => to_unsigned(957, 10), 1706 => to_unsigned(633, 10), 1707 => to_unsigned(125, 10), 1708 => to_unsigned(294, 10), 1709 => to_unsigned(805, 10), 1710 => to_unsigned(338, 10), 1711 => to_unsigned(428, 10), 1712 => to_unsigned(476, 10), 1713 => to_unsigned(318, 10), 1714 => to_unsigned(369, 10), 1715 => to_unsigned(963, 10), 1716 => to_unsigned(236, 10), 1717 => to_unsigned(934, 10), 1718 => to_unsigned(996, 10), 1719 => to_unsigned(299, 10), 1720 => to_unsigned(259, 10), 1721 => to_unsigned(518, 10), 1722 => to_unsigned(111, 10), 1723 => to_unsigned(689, 10), 1724 => to_unsigned(12, 10), 1725 => to_unsigned(21, 10), 1726 => to_unsigned(400, 10), 1727 => to_unsigned(364, 10), 1728 => to_unsigned(697, 10), 1729 => to_unsigned(882, 10), 1730 => to_unsigned(521, 10), 1731 => to_unsigned(677, 10), 1732 => to_unsigned(389, 10), 1733 => to_unsigned(73, 10), 1734 => to_unsigned(1019, 10), 1735 => to_unsigned(245, 10), 1736 => to_unsigned(839, 10), 1737 => to_unsigned(369, 10), 1738 => to_unsigned(488, 10), 1739 => to_unsigned(578, 10), 1740 => to_unsigned(226, 10), 1741 => to_unsigned(678, 10), 1742 => to_unsigned(637, 10), 1743 => to_unsigned(699, 10), 1744 => to_unsigned(888, 10), 1745 => to_unsigned(276, 10), 1746 => to_unsigned(45, 10), 1747 => to_unsigned(783, 10), 1748 => to_unsigned(785, 10), 1749 => to_unsigned(810, 10), 1750 => to_unsigned(244, 10), 1751 => to_unsigned(704, 10), 1752 => to_unsigned(740, 10), 1753 => to_unsigned(5, 10), 1754 => to_unsigned(986, 10), 1755 => to_unsigned(138, 10), 1756 => to_unsigned(92, 10), 1757 => to_unsigned(654, 10), 1758 => to_unsigned(553, 10), 1759 => to_unsigned(883, 10), 1760 => to_unsigned(751, 10), 1761 => to_unsigned(842, 10), 1762 => to_unsigned(19, 10), 1763 => to_unsigned(798, 10), 1764 => to_unsigned(483, 10), 1765 => to_unsigned(896, 10), 1766 => to_unsigned(489, 10), 1767 => to_unsigned(696, 10), 1768 => to_unsigned(408, 10), 1769 => to_unsigned(197, 10), 1770 => to_unsigned(656, 10), 1771 => to_unsigned(316, 10), 1772 => to_unsigned(890, 10), 1773 => to_unsigned(244, 10), 1774 => to_unsigned(211, 10), 1775 => to_unsigned(492, 10), 1776 => to_unsigned(108, 10), 1777 => to_unsigned(674, 10), 1778 => to_unsigned(561, 10), 1779 => to_unsigned(707, 10), 1780 => to_unsigned(303, 10), 1781 => to_unsigned(46, 10), 1782 => to_unsigned(1000, 10), 1783 => to_unsigned(955, 10), 1784 => to_unsigned(430, 10), 1785 => to_unsigned(986, 10), 1786 => to_unsigned(962, 10), 1787 => to_unsigned(274, 10), 1788 => to_unsigned(19, 10), 1789 => to_unsigned(229, 10), 1790 => to_unsigned(231, 10), 1791 => to_unsigned(953, 10), 1792 => to_unsigned(200, 10), 1793 => to_unsigned(440, 10), 1794 => to_unsigned(618, 10), 1795 => to_unsigned(856, 10), 1796 => to_unsigned(60, 10), 1797 => to_unsigned(872, 10), 1798 => to_unsigned(238, 10), 1799 => to_unsigned(387, 10), 1800 => to_unsigned(987, 10), 1801 => to_unsigned(657, 10), 1802 => to_unsigned(665, 10), 1803 => to_unsigned(911, 10), 1804 => to_unsigned(779, 10), 1805 => to_unsigned(228, 10), 1806 => to_unsigned(1017, 10), 1807 => to_unsigned(203, 10), 1808 => to_unsigned(205, 10), 1809 => to_unsigned(828, 10), 1810 => to_unsigned(469, 10), 1811 => to_unsigned(423, 10), 1812 => to_unsigned(73, 10), 1813 => to_unsigned(228, 10), 1814 => to_unsigned(877, 10), 1815 => to_unsigned(114, 10), 1816 => to_unsigned(811, 10), 1817 => to_unsigned(49, 10), 1818 => to_unsigned(167, 10), 1819 => to_unsigned(640, 10), 1820 => to_unsigned(287, 10), 1821 => to_unsigned(791, 10), 1822 => to_unsigned(621, 10), 1823 => to_unsigned(1005, 10), 1824 => to_unsigned(906, 10), 1825 => to_unsigned(671, 10), 1826 => to_unsigned(336, 10), 1827 => to_unsigned(127, 10), 1828 => to_unsigned(364, 10), 1829 => to_unsigned(882, 10), 1830 => to_unsigned(333, 10), 1831 => to_unsigned(890, 10), 1832 => to_unsigned(219, 10), 1833 => to_unsigned(422, 10), 1834 => to_unsigned(290, 10), 1835 => to_unsigned(395, 10), 1836 => to_unsigned(325, 10), 1837 => to_unsigned(38, 10), 1838 => to_unsigned(248, 10), 1839 => to_unsigned(453, 10), 1840 => to_unsigned(880, 10), 1841 => to_unsigned(504, 10), 1842 => to_unsigned(661, 10), 1843 => to_unsigned(545, 10), 1844 => to_unsigned(693, 10), 1845 => to_unsigned(288, 10), 1846 => to_unsigned(689, 10), 1847 => to_unsigned(682, 10), 1848 => to_unsigned(569, 10), 1849 => to_unsigned(865, 10), 1850 => to_unsigned(142, 10), 1851 => to_unsigned(1021, 10), 1852 => to_unsigned(552, 10), 1853 => to_unsigned(890, 10), 1854 => to_unsigned(152, 10), 1855 => to_unsigned(526, 10), 1856 => to_unsigned(13, 10), 1857 => to_unsigned(116, 10), 1858 => to_unsigned(978, 10), 1859 => to_unsigned(81, 10), 1860 => to_unsigned(869, 10), 1861 => to_unsigned(712, 10), 1862 => to_unsigned(26, 10), 1863 => to_unsigned(82, 10), 1864 => to_unsigned(508, 10), 1865 => to_unsigned(117, 10), 1866 => to_unsigned(282, 10), 1867 => to_unsigned(679, 10), 1868 => to_unsigned(958, 10), 1869 => to_unsigned(288, 10), 1870 => to_unsigned(101, 10), 1871 => to_unsigned(725, 10), 1872 => to_unsigned(775, 10), 1873 => to_unsigned(743, 10), 1874 => to_unsigned(358, 10), 1875 => to_unsigned(273, 10), 1876 => to_unsigned(599, 10), 1877 => to_unsigned(53, 10), 1878 => to_unsigned(763, 10), 1879 => to_unsigned(915, 10), 1880 => to_unsigned(676, 10), 1881 => to_unsigned(456, 10), 1882 => to_unsigned(585, 10), 1883 => to_unsigned(561, 10), 1884 => to_unsigned(893, 10), 1885 => to_unsigned(929, 10), 1886 => to_unsigned(171, 10), 1887 => to_unsigned(645, 10), 1888 => to_unsigned(17, 10), 1889 => to_unsigned(187, 10), 1890 => to_unsigned(1012, 10), 1891 => to_unsigned(591, 10), 1892 => to_unsigned(992, 10), 1893 => to_unsigned(567, 10), 1894 => to_unsigned(266, 10), 1895 => to_unsigned(458, 10), 1896 => to_unsigned(942, 10), 1897 => to_unsigned(1013, 10), 1898 => to_unsigned(165, 10), 1899 => to_unsigned(614, 10), 1900 => to_unsigned(976, 10), 1901 => to_unsigned(4, 10), 1902 => to_unsigned(421, 10), 1903 => to_unsigned(681, 10), 1904 => to_unsigned(310, 10), 1905 => to_unsigned(169, 10), 1906 => to_unsigned(78, 10), 1907 => to_unsigned(153, 10), 1908 => to_unsigned(293, 10), 1909 => to_unsigned(690, 10), 1910 => to_unsigned(628, 10), 1911 => to_unsigned(892, 10), 1912 => to_unsigned(870, 10), 1913 => to_unsigned(48, 10), 1914 => to_unsigned(795, 10), 1915 => to_unsigned(857, 10), 1916 => to_unsigned(756, 10), 1917 => to_unsigned(579, 10), 1918 => to_unsigned(559, 10), 1919 => to_unsigned(179, 10), 1920 => to_unsigned(152, 10), 1921 => to_unsigned(272, 10), 1922 => to_unsigned(25, 10), 1923 => to_unsigned(108, 10), 1924 => to_unsigned(609, 10), 1925 => to_unsigned(180, 10), 1926 => to_unsigned(163, 10), 1927 => to_unsigned(787, 10), 1928 => to_unsigned(1019, 10), 1929 => to_unsigned(642, 10), 1930 => to_unsigned(633, 10), 1931 => to_unsigned(716, 10), 1932 => to_unsigned(882, 10), 1933 => to_unsigned(958, 10), 1934 => to_unsigned(673, 10), 1935 => to_unsigned(952, 10), 1936 => to_unsigned(524, 10), 1937 => to_unsigned(840, 10), 1938 => to_unsigned(59, 10), 1939 => to_unsigned(726, 10), 1940 => to_unsigned(573, 10), 1941 => to_unsigned(367, 10), 1942 => to_unsigned(240, 10), 1943 => to_unsigned(969, 10), 1944 => to_unsigned(680, 10), 1945 => to_unsigned(796, 10), 1946 => to_unsigned(123, 10), 1947 => to_unsigned(857, 10), 1948 => to_unsigned(414, 10), 1949 => to_unsigned(504, 10), 1950 => to_unsigned(806, 10), 1951 => to_unsigned(895, 10), 1952 => to_unsigned(502, 10), 1953 => to_unsigned(579, 10), 1954 => to_unsigned(842, 10), 1955 => to_unsigned(265, 10), 1956 => to_unsigned(63, 10), 1957 => to_unsigned(125, 10), 1958 => to_unsigned(1011, 10), 1959 => to_unsigned(760, 10), 1960 => to_unsigned(29, 10), 1961 => to_unsigned(623, 10), 1962 => to_unsigned(388, 10), 1963 => to_unsigned(162, 10), 1964 => to_unsigned(445, 10), 1965 => to_unsigned(110, 10), 1966 => to_unsigned(103, 10), 1967 => to_unsigned(295, 10), 1968 => to_unsigned(290, 10), 1969 => to_unsigned(1008, 10), 1970 => to_unsigned(8, 10), 1971 => to_unsigned(599, 10), 1972 => to_unsigned(683, 10), 1973 => to_unsigned(602, 10), 1974 => to_unsigned(557, 10), 1975 => to_unsigned(187, 10), 1976 => to_unsigned(642, 10), 1977 => to_unsigned(295, 10), 1978 => to_unsigned(414, 10), 1979 => to_unsigned(65, 10), 1980 => to_unsigned(533, 10), 1981 => to_unsigned(74, 10), 1982 => to_unsigned(171, 10), 1983 => to_unsigned(519, 10), 1984 => to_unsigned(40, 10), 1985 => to_unsigned(737, 10), 1986 => to_unsigned(577, 10), 1987 => to_unsigned(105, 10), 1988 => to_unsigned(970, 10), 1989 => to_unsigned(127, 10), 1990 => to_unsigned(930, 10), 1991 => to_unsigned(26, 10), 1992 => to_unsigned(330, 10), 1993 => to_unsigned(409, 10), 1994 => to_unsigned(408, 10), 1995 => to_unsigned(598, 10), 1996 => to_unsigned(430, 10), 1997 => to_unsigned(510, 10), 1998 => to_unsigned(907, 10), 1999 => to_unsigned(665, 10), 2000 => to_unsigned(284, 10), 2001 => to_unsigned(993, 10), 2002 => to_unsigned(204, 10), 2003 => to_unsigned(573, 10), 2004 => to_unsigned(164, 10), 2005 => to_unsigned(53, 10), 2006 => to_unsigned(817, 10), 2007 => to_unsigned(431, 10), 2008 => to_unsigned(510, 10), 2009 => to_unsigned(310, 10), 2010 => to_unsigned(248, 10), 2011 => to_unsigned(225, 10), 2012 => to_unsigned(468, 10), 2013 => to_unsigned(919, 10), 2014 => to_unsigned(674, 10), 2015 => to_unsigned(710, 10), 2016 => to_unsigned(827, 10), 2017 => to_unsigned(925, 10), 2018 => to_unsigned(166, 10), 2019 => to_unsigned(665, 10), 2020 => to_unsigned(911, 10), 2021 => to_unsigned(202, 10), 2022 => to_unsigned(647, 10), 2023 => to_unsigned(500, 10), 2024 => to_unsigned(195, 10), 2025 => to_unsigned(490, 10), 2026 => to_unsigned(580, 10), 2027 => to_unsigned(823, 10), 2028 => to_unsigned(800, 10), 2029 => to_unsigned(989, 10), 2030 => to_unsigned(868, 10), 2031 => to_unsigned(246, 10), 2032 => to_unsigned(50, 10), 2033 => to_unsigned(250, 10), 2034 => to_unsigned(260, 10), 2035 => to_unsigned(681, 10), 2036 => to_unsigned(873, 10), 2037 => to_unsigned(779, 10), 2038 => to_unsigned(524, 10), 2039 => to_unsigned(262, 10), 2040 => to_unsigned(793, 10), 2041 => to_unsigned(207, 10), 2042 => to_unsigned(864, 10), 2043 => to_unsigned(46, 10), 2044 => to_unsigned(342, 10), 2045 => to_unsigned(439, 10), 2046 => to_unsigned(448, 10), 2047 => to_unsigned(373, 10)),
            3 => (0 => to_unsigned(171, 10), 1 => to_unsigned(649, 10), 2 => to_unsigned(594, 10), 3 => to_unsigned(357, 10), 4 => to_unsigned(237, 10), 5 => to_unsigned(899, 10), 6 => to_unsigned(922, 10), 7 => to_unsigned(548, 10), 8 => to_unsigned(8, 10), 9 => to_unsigned(82, 10), 10 => to_unsigned(222, 10), 11 => to_unsigned(848, 10), 12 => to_unsigned(748, 10), 13 => to_unsigned(424, 10), 14 => to_unsigned(167, 10), 15 => to_unsigned(237, 10), 16 => to_unsigned(436, 10), 17 => to_unsigned(437, 10), 18 => to_unsigned(542, 10), 19 => to_unsigned(167, 10), 20 => to_unsigned(74, 10), 21 => to_unsigned(747, 10), 22 => to_unsigned(498, 10), 23 => to_unsigned(148, 10), 24 => to_unsigned(546, 10), 25 => to_unsigned(873, 10), 26 => to_unsigned(578, 10), 27 => to_unsigned(607, 10), 28 => to_unsigned(518, 10), 29 => to_unsigned(444, 10), 30 => to_unsigned(327, 10), 31 => to_unsigned(864, 10), 32 => to_unsigned(678, 10), 33 => to_unsigned(101, 10), 34 => to_unsigned(812, 10), 35 => to_unsigned(708, 10), 36 => to_unsigned(501, 10), 37 => to_unsigned(444, 10), 38 => to_unsigned(241, 10), 39 => to_unsigned(23, 10), 40 => to_unsigned(941, 10), 41 => to_unsigned(165, 10), 42 => to_unsigned(664, 10), 43 => to_unsigned(186, 10), 44 => to_unsigned(478, 10), 45 => to_unsigned(52, 10), 46 => to_unsigned(101, 10), 47 => to_unsigned(322, 10), 48 => to_unsigned(1022, 10), 49 => to_unsigned(348, 10), 50 => to_unsigned(958, 10), 51 => to_unsigned(202, 10), 52 => to_unsigned(967, 10), 53 => to_unsigned(774, 10), 54 => to_unsigned(984, 10), 55 => to_unsigned(452, 10), 56 => to_unsigned(646, 10), 57 => to_unsigned(906, 10), 58 => to_unsigned(962, 10), 59 => to_unsigned(473, 10), 60 => to_unsigned(754, 10), 61 => to_unsigned(604, 10), 62 => to_unsigned(160, 10), 63 => to_unsigned(591, 10), 64 => to_unsigned(829, 10), 65 => to_unsigned(974, 10), 66 => to_unsigned(769, 10), 67 => to_unsigned(780, 10), 68 => to_unsigned(339, 10), 69 => to_unsigned(25, 10), 70 => to_unsigned(589, 10), 71 => to_unsigned(67, 10), 72 => to_unsigned(1003, 10), 73 => to_unsigned(846, 10), 74 => to_unsigned(790, 10), 75 => to_unsigned(234, 10), 76 => to_unsigned(819, 10), 77 => to_unsigned(799, 10), 78 => to_unsigned(274, 10), 79 => to_unsigned(48, 10), 80 => to_unsigned(389, 10), 81 => to_unsigned(651, 10), 82 => to_unsigned(629, 10), 83 => to_unsigned(707, 10), 84 => to_unsigned(634, 10), 85 => to_unsigned(307, 10), 86 => to_unsigned(295, 10), 87 => to_unsigned(972, 10), 88 => to_unsigned(903, 10), 89 => to_unsigned(888, 10), 90 => to_unsigned(450, 10), 91 => to_unsigned(105, 10), 92 => to_unsigned(697, 10), 93 => to_unsigned(699, 10), 94 => to_unsigned(173, 10), 95 => to_unsigned(169, 10), 96 => to_unsigned(591, 10), 97 => to_unsigned(793, 10), 98 => to_unsigned(440, 10), 99 => to_unsigned(1016, 10), 100 => to_unsigned(27, 10), 101 => to_unsigned(664, 10), 102 => to_unsigned(253, 10), 103 => to_unsigned(582, 10), 104 => to_unsigned(553, 10), 105 => to_unsigned(814, 10), 106 => to_unsigned(489, 10), 107 => to_unsigned(835, 10), 108 => to_unsigned(68, 10), 109 => to_unsigned(565, 10), 110 => to_unsigned(784, 10), 111 => to_unsigned(84, 10), 112 => to_unsigned(938, 10), 113 => to_unsigned(238, 10), 114 => to_unsigned(618, 10), 115 => to_unsigned(224, 10), 116 => to_unsigned(772, 10), 117 => to_unsigned(513, 10), 118 => to_unsigned(851, 10), 119 => to_unsigned(858, 10), 120 => to_unsigned(529, 10), 121 => to_unsigned(909, 10), 122 => to_unsigned(872, 10), 123 => to_unsigned(24, 10), 124 => to_unsigned(237, 10), 125 => to_unsigned(849, 10), 126 => to_unsigned(112, 10), 127 => to_unsigned(263, 10), 128 => to_unsigned(697, 10), 129 => to_unsigned(396, 10), 130 => to_unsigned(932, 10), 131 => to_unsigned(968, 10), 132 => to_unsigned(274, 10), 133 => to_unsigned(206, 10), 134 => to_unsigned(376, 10), 135 => to_unsigned(177, 10), 136 => to_unsigned(453, 10), 137 => to_unsigned(250, 10), 138 => to_unsigned(518, 10), 139 => to_unsigned(983, 10), 140 => to_unsigned(712, 10), 141 => to_unsigned(845, 10), 142 => to_unsigned(916, 10), 143 => to_unsigned(231, 10), 144 => to_unsigned(624, 10), 145 => to_unsigned(715, 10), 146 => to_unsigned(473, 10), 147 => to_unsigned(756, 10), 148 => to_unsigned(77, 10), 149 => to_unsigned(705, 10), 150 => to_unsigned(517, 10), 151 => to_unsigned(707, 10), 152 => to_unsigned(764, 10), 153 => to_unsigned(528, 10), 154 => to_unsigned(878, 10), 155 => to_unsigned(122, 10), 156 => to_unsigned(992, 10), 157 => to_unsigned(84, 10), 158 => to_unsigned(427, 10), 159 => to_unsigned(620, 10), 160 => to_unsigned(225, 10), 161 => to_unsigned(512, 10), 162 => to_unsigned(239, 10), 163 => to_unsigned(301, 10), 164 => to_unsigned(15, 10), 165 => to_unsigned(400, 10), 166 => to_unsigned(938, 10), 167 => to_unsigned(258, 10), 168 => to_unsigned(528, 10), 169 => to_unsigned(468, 10), 170 => to_unsigned(37, 10), 171 => to_unsigned(172, 10), 172 => to_unsigned(165, 10), 173 => to_unsigned(298, 10), 174 => to_unsigned(129, 10), 175 => to_unsigned(870, 10), 176 => to_unsigned(754, 10), 177 => to_unsigned(58, 10), 178 => to_unsigned(642, 10), 179 => to_unsigned(398, 10), 180 => to_unsigned(233, 10), 181 => to_unsigned(716, 10), 182 => to_unsigned(986, 10), 183 => to_unsigned(160, 10), 184 => to_unsigned(879, 10), 185 => to_unsigned(987, 10), 186 => to_unsigned(198, 10), 187 => to_unsigned(426, 10), 188 => to_unsigned(59, 10), 189 => to_unsigned(232, 10), 190 => to_unsigned(477, 10), 191 => to_unsigned(871, 10), 192 => to_unsigned(747, 10), 193 => to_unsigned(295, 10), 194 => to_unsigned(977, 10), 195 => to_unsigned(302, 10), 196 => to_unsigned(232, 10), 197 => to_unsigned(605, 10), 198 => to_unsigned(436, 10), 199 => to_unsigned(560, 10), 200 => to_unsigned(201, 10), 201 => to_unsigned(245, 10), 202 => to_unsigned(849, 10), 203 => to_unsigned(703, 10), 204 => to_unsigned(714, 10), 205 => to_unsigned(396, 10), 206 => to_unsigned(381, 10), 207 => to_unsigned(495, 10), 208 => to_unsigned(638, 10), 209 => to_unsigned(991, 10), 210 => to_unsigned(641, 10), 211 => to_unsigned(281, 10), 212 => to_unsigned(152, 10), 213 => to_unsigned(589, 10), 214 => to_unsigned(233, 10), 215 => to_unsigned(222, 10), 216 => to_unsigned(241, 10), 217 => to_unsigned(812, 10), 218 => to_unsigned(567, 10), 219 => to_unsigned(874, 10), 220 => to_unsigned(936, 10), 221 => to_unsigned(1013, 10), 222 => to_unsigned(236, 10), 223 => to_unsigned(286, 10), 224 => to_unsigned(441, 10), 225 => to_unsigned(531, 10), 226 => to_unsigned(732, 10), 227 => to_unsigned(944, 10), 228 => to_unsigned(262, 10), 229 => to_unsigned(876, 10), 230 => to_unsigned(74, 10), 231 => to_unsigned(246, 10), 232 => to_unsigned(680, 10), 233 => to_unsigned(979, 10), 234 => to_unsigned(624, 10), 235 => to_unsigned(824, 10), 236 => to_unsigned(262, 10), 237 => to_unsigned(549, 10), 238 => to_unsigned(976, 10), 239 => to_unsigned(5, 10), 240 => to_unsigned(418, 10), 241 => to_unsigned(908, 10), 242 => to_unsigned(861, 10), 243 => to_unsigned(882, 10), 244 => to_unsigned(788, 10), 245 => to_unsigned(93, 10), 246 => to_unsigned(266, 10), 247 => to_unsigned(475, 10), 248 => to_unsigned(306, 10), 249 => to_unsigned(764, 10), 250 => to_unsigned(225, 10), 251 => to_unsigned(490, 10), 252 => to_unsigned(458, 10), 253 => to_unsigned(221, 10), 254 => to_unsigned(522, 10), 255 => to_unsigned(911, 10), 256 => to_unsigned(182, 10), 257 => to_unsigned(657, 10), 258 => to_unsigned(349, 10), 259 => to_unsigned(848, 10), 260 => to_unsigned(824, 10), 261 => to_unsigned(76, 10), 262 => to_unsigned(988, 10), 263 => to_unsigned(772, 10), 264 => to_unsigned(262, 10), 265 => to_unsigned(621, 10), 266 => to_unsigned(958, 10), 267 => to_unsigned(375, 10), 268 => to_unsigned(50, 10), 269 => to_unsigned(561, 10), 270 => to_unsigned(812, 10), 271 => to_unsigned(170, 10), 272 => to_unsigned(158, 10), 273 => to_unsigned(339, 10), 274 => to_unsigned(658, 10), 275 => to_unsigned(930, 10), 276 => to_unsigned(285, 10), 277 => to_unsigned(846, 10), 278 => to_unsigned(910, 10), 279 => to_unsigned(492, 10), 280 => to_unsigned(762, 10), 281 => to_unsigned(130, 10), 282 => to_unsigned(250, 10), 283 => to_unsigned(193, 10), 284 => to_unsigned(903, 10), 285 => to_unsigned(369, 10), 286 => to_unsigned(290, 10), 287 => to_unsigned(472, 10), 288 => to_unsigned(927, 10), 289 => to_unsigned(109, 10), 290 => to_unsigned(705, 10), 291 => to_unsigned(380, 10), 292 => to_unsigned(356, 10), 293 => to_unsigned(325, 10), 294 => to_unsigned(164, 10), 295 => to_unsigned(521, 10), 296 => to_unsigned(439, 10), 297 => to_unsigned(71, 10), 298 => to_unsigned(54, 10), 299 => to_unsigned(195, 10), 300 => to_unsigned(401, 10), 301 => to_unsigned(610, 10), 302 => to_unsigned(618, 10), 303 => to_unsigned(856, 10), 304 => to_unsigned(829, 10), 305 => to_unsigned(687, 10), 306 => to_unsigned(862, 10), 307 => to_unsigned(868, 10), 308 => to_unsigned(808, 10), 309 => to_unsigned(671, 10), 310 => to_unsigned(9, 10), 311 => to_unsigned(363, 10), 312 => to_unsigned(16, 10), 313 => to_unsigned(978, 10), 314 => to_unsigned(406, 10), 315 => to_unsigned(585, 10), 316 => to_unsigned(127, 10), 317 => to_unsigned(29, 10), 318 => to_unsigned(835, 10), 319 => to_unsigned(196, 10), 320 => to_unsigned(905, 10), 321 => to_unsigned(757, 10), 322 => to_unsigned(464, 10), 323 => to_unsigned(986, 10), 324 => to_unsigned(671, 10), 325 => to_unsigned(199, 10), 326 => to_unsigned(536, 10), 327 => to_unsigned(81, 10), 328 => to_unsigned(614, 10), 329 => to_unsigned(257, 10), 330 => to_unsigned(741, 10), 331 => to_unsigned(283, 10), 332 => to_unsigned(676, 10), 333 => to_unsigned(838, 10), 334 => to_unsigned(570, 10), 335 => to_unsigned(333, 10), 336 => to_unsigned(5, 10), 337 => to_unsigned(240, 10), 338 => to_unsigned(951, 10), 339 => to_unsigned(792, 10), 340 => to_unsigned(518, 10), 341 => to_unsigned(1006, 10), 342 => to_unsigned(362, 10), 343 => to_unsigned(753, 10), 344 => to_unsigned(886, 10), 345 => to_unsigned(465, 10), 346 => to_unsigned(1020, 10), 347 => to_unsigned(690, 10), 348 => to_unsigned(333, 10), 349 => to_unsigned(486, 10), 350 => to_unsigned(837, 10), 351 => to_unsigned(616, 10), 352 => to_unsigned(262, 10), 353 => to_unsigned(852, 10), 354 => to_unsigned(307, 10), 355 => to_unsigned(412, 10), 356 => to_unsigned(173, 10), 357 => to_unsigned(733, 10), 358 => to_unsigned(433, 10), 359 => to_unsigned(799, 10), 360 => to_unsigned(376, 10), 361 => to_unsigned(1001, 10), 362 => to_unsigned(293, 10), 363 => to_unsigned(383, 10), 364 => to_unsigned(219, 10), 365 => to_unsigned(696, 10), 366 => to_unsigned(960, 10), 367 => to_unsigned(42, 10), 368 => to_unsigned(725, 10), 369 => to_unsigned(680, 10), 370 => to_unsigned(715, 10), 371 => to_unsigned(517, 10), 372 => to_unsigned(873, 10), 373 => to_unsigned(10, 10), 374 => to_unsigned(930, 10), 375 => to_unsigned(984, 10), 376 => to_unsigned(779, 10), 377 => to_unsigned(418, 10), 378 => to_unsigned(671, 10), 379 => to_unsigned(196, 10), 380 => to_unsigned(411, 10), 381 => to_unsigned(39, 10), 382 => to_unsigned(916, 10), 383 => to_unsigned(409, 10), 384 => to_unsigned(450, 10), 385 => to_unsigned(257, 10), 386 => to_unsigned(233, 10), 387 => to_unsigned(911, 10), 388 => to_unsigned(915, 10), 389 => to_unsigned(302, 10), 390 => to_unsigned(340, 10), 391 => to_unsigned(992, 10), 392 => to_unsigned(974, 10), 393 => to_unsigned(44, 10), 394 => to_unsigned(873, 10), 395 => to_unsigned(135, 10), 396 => to_unsigned(137, 10), 397 => to_unsigned(908, 10), 398 => to_unsigned(851, 10), 399 => to_unsigned(312, 10), 400 => to_unsigned(294, 10), 401 => to_unsigned(813, 10), 402 => to_unsigned(739, 10), 403 => to_unsigned(942, 10), 404 => to_unsigned(688, 10), 405 => to_unsigned(825, 10), 406 => to_unsigned(658, 10), 407 => to_unsigned(434, 10), 408 => to_unsigned(163, 10), 409 => to_unsigned(264, 10), 410 => to_unsigned(1022, 10), 411 => to_unsigned(486, 10), 412 => to_unsigned(471, 10), 413 => to_unsigned(16, 10), 414 => to_unsigned(264, 10), 415 => to_unsigned(699, 10), 416 => to_unsigned(373, 10), 417 => to_unsigned(236, 10), 418 => to_unsigned(563, 10), 419 => to_unsigned(280, 10), 420 => to_unsigned(908, 10), 421 => to_unsigned(552, 10), 422 => to_unsigned(533, 10), 423 => to_unsigned(475, 10), 424 => to_unsigned(921, 10), 425 => to_unsigned(929, 10), 426 => to_unsigned(844, 10), 427 => to_unsigned(756, 10), 428 => to_unsigned(363, 10), 429 => to_unsigned(489, 10), 430 => to_unsigned(514, 10), 431 => to_unsigned(35, 10), 432 => to_unsigned(408, 10), 433 => to_unsigned(839, 10), 434 => to_unsigned(267, 10), 435 => to_unsigned(312, 10), 436 => to_unsigned(39, 10), 437 => to_unsigned(335, 10), 438 => to_unsigned(808, 10), 439 => to_unsigned(971, 10), 440 => to_unsigned(226, 10), 441 => to_unsigned(353, 10), 442 => to_unsigned(294, 10), 443 => to_unsigned(496, 10), 444 => to_unsigned(644, 10), 445 => to_unsigned(460, 10), 446 => to_unsigned(674, 10), 447 => to_unsigned(156, 10), 448 => to_unsigned(365, 10), 449 => to_unsigned(973, 10), 450 => to_unsigned(111, 10), 451 => to_unsigned(677, 10), 452 => to_unsigned(330, 10), 453 => to_unsigned(482, 10), 454 => to_unsigned(955, 10), 455 => to_unsigned(227, 10), 456 => to_unsigned(837, 10), 457 => to_unsigned(215, 10), 458 => to_unsigned(114, 10), 459 => to_unsigned(25, 10), 460 => to_unsigned(22, 10), 461 => to_unsigned(414, 10), 462 => to_unsigned(90, 10), 463 => to_unsigned(947, 10), 464 => to_unsigned(941, 10), 465 => to_unsigned(190, 10), 466 => to_unsigned(354, 10), 467 => to_unsigned(407, 10), 468 => to_unsigned(114, 10), 469 => to_unsigned(112, 10), 470 => to_unsigned(419, 10), 471 => to_unsigned(654, 10), 472 => to_unsigned(413, 10), 473 => to_unsigned(334, 10), 474 => to_unsigned(83, 10), 475 => to_unsigned(290, 10), 476 => to_unsigned(45, 10), 477 => to_unsigned(310, 10), 478 => to_unsigned(97, 10), 479 => to_unsigned(829, 10), 480 => to_unsigned(602, 10), 481 => to_unsigned(836, 10), 482 => to_unsigned(467, 10), 483 => to_unsigned(109, 10), 484 => to_unsigned(415, 10), 485 => to_unsigned(886, 10), 486 => to_unsigned(798, 10), 487 => to_unsigned(494, 10), 488 => to_unsigned(418, 10), 489 => to_unsigned(375, 10), 490 => to_unsigned(112, 10), 491 => to_unsigned(545, 10), 492 => to_unsigned(515, 10), 493 => to_unsigned(671, 10), 494 => to_unsigned(914, 10), 495 => to_unsigned(509, 10), 496 => to_unsigned(112, 10), 497 => to_unsigned(669, 10), 498 => to_unsigned(801, 10), 499 => to_unsigned(983, 10), 500 => to_unsigned(189, 10), 501 => to_unsigned(463, 10), 502 => to_unsigned(861, 10), 503 => to_unsigned(325, 10), 504 => to_unsigned(389, 10), 505 => to_unsigned(253, 10), 506 => to_unsigned(644, 10), 507 => to_unsigned(909, 10), 508 => to_unsigned(678, 10), 509 => to_unsigned(481, 10), 510 => to_unsigned(979, 10), 511 => to_unsigned(883, 10), 512 => to_unsigned(414, 10), 513 => to_unsigned(500, 10), 514 => to_unsigned(899, 10), 515 => to_unsigned(637, 10), 516 => to_unsigned(477, 10), 517 => to_unsigned(12, 10), 518 => to_unsigned(275, 10), 519 => to_unsigned(527, 10), 520 => to_unsigned(13, 10), 521 => to_unsigned(354, 10), 522 => to_unsigned(340, 10), 523 => to_unsigned(283, 10), 524 => to_unsigned(467, 10), 525 => to_unsigned(350, 10), 526 => to_unsigned(237, 10), 527 => to_unsigned(83, 10), 528 => to_unsigned(222, 10), 529 => to_unsigned(225, 10), 530 => to_unsigned(499, 10), 531 => to_unsigned(533, 10), 532 => to_unsigned(465, 10), 533 => to_unsigned(323, 10), 534 => to_unsigned(919, 10), 535 => to_unsigned(398, 10), 536 => to_unsigned(116, 10), 537 => to_unsigned(55, 10), 538 => to_unsigned(738, 10), 539 => to_unsigned(785, 10), 540 => to_unsigned(101, 10), 541 => to_unsigned(834, 10), 542 => to_unsigned(726, 10), 543 => to_unsigned(57, 10), 544 => to_unsigned(319, 10), 545 => to_unsigned(15, 10), 546 => to_unsigned(518, 10), 547 => to_unsigned(740, 10), 548 => to_unsigned(469, 10), 549 => to_unsigned(203, 10), 550 => to_unsigned(843, 10), 551 => to_unsigned(819, 10), 552 => to_unsigned(110, 10), 553 => to_unsigned(966, 10), 554 => to_unsigned(343, 10), 555 => to_unsigned(914, 10), 556 => to_unsigned(781, 10), 557 => to_unsigned(627, 10), 558 => to_unsigned(119, 10), 559 => to_unsigned(88, 10), 560 => to_unsigned(327, 10), 561 => to_unsigned(887, 10), 562 => to_unsigned(165, 10), 563 => to_unsigned(226, 10), 564 => to_unsigned(259, 10), 565 => to_unsigned(765, 10), 566 => to_unsigned(690, 10), 567 => to_unsigned(466, 10), 568 => to_unsigned(919, 10), 569 => to_unsigned(993, 10), 570 => to_unsigned(565, 10), 571 => to_unsigned(69, 10), 572 => to_unsigned(431, 10), 573 => to_unsigned(222, 10), 574 => to_unsigned(921, 10), 575 => to_unsigned(693, 10), 576 => to_unsigned(241, 10), 577 => to_unsigned(387, 10), 578 => to_unsigned(136, 10), 579 => to_unsigned(649, 10), 580 => to_unsigned(894, 10), 581 => to_unsigned(88, 10), 582 => to_unsigned(561, 10), 583 => to_unsigned(940, 10), 584 => to_unsigned(30, 10), 585 => to_unsigned(459, 10), 586 => to_unsigned(190, 10), 587 => to_unsigned(386, 10), 588 => to_unsigned(432, 10), 589 => to_unsigned(340, 10), 590 => to_unsigned(175, 10), 591 => to_unsigned(267, 10), 592 => to_unsigned(224, 10), 593 => to_unsigned(796, 10), 594 => to_unsigned(243, 10), 595 => to_unsigned(613, 10), 596 => to_unsigned(235, 10), 597 => to_unsigned(165, 10), 598 => to_unsigned(294, 10), 599 => to_unsigned(950, 10), 600 => to_unsigned(803, 10), 601 => to_unsigned(906, 10), 602 => to_unsigned(447, 10), 603 => to_unsigned(665, 10), 604 => to_unsigned(821, 10), 605 => to_unsigned(91, 10), 606 => to_unsigned(468, 10), 607 => to_unsigned(58, 10), 608 => to_unsigned(1023, 10), 609 => to_unsigned(973, 10), 610 => to_unsigned(90, 10), 611 => to_unsigned(406, 10), 612 => to_unsigned(182, 10), 613 => to_unsigned(451, 10), 614 => to_unsigned(534, 10), 615 => to_unsigned(669, 10), 616 => to_unsigned(831, 10), 617 => to_unsigned(697, 10), 618 => to_unsigned(623, 10), 619 => to_unsigned(754, 10), 620 => to_unsigned(869, 10), 621 => to_unsigned(684, 10), 622 => to_unsigned(768, 10), 623 => to_unsigned(742, 10), 624 => to_unsigned(204, 10), 625 => to_unsigned(207, 10), 626 => to_unsigned(906, 10), 627 => to_unsigned(492, 10), 628 => to_unsigned(459, 10), 629 => to_unsigned(997, 10), 630 => to_unsigned(365, 10), 631 => to_unsigned(503, 10), 632 => to_unsigned(721, 10), 633 => to_unsigned(839, 10), 634 => to_unsigned(277, 10), 635 => to_unsigned(23, 10), 636 => to_unsigned(867, 10), 637 => to_unsigned(522, 10), 638 => to_unsigned(174, 10), 639 => to_unsigned(373, 10), 640 => to_unsigned(785, 10), 641 => to_unsigned(523, 10), 642 => to_unsigned(39, 10), 643 => to_unsigned(552, 10), 644 => to_unsigned(191, 10), 645 => to_unsigned(392, 10), 646 => to_unsigned(183, 10), 647 => to_unsigned(914, 10), 648 => to_unsigned(44, 10), 649 => to_unsigned(902, 10), 650 => to_unsigned(484, 10), 651 => to_unsigned(1005, 10), 652 => to_unsigned(351, 10), 653 => to_unsigned(529, 10), 654 => to_unsigned(364, 10), 655 => to_unsigned(258, 10), 656 => to_unsigned(818, 10), 657 => to_unsigned(135, 10), 658 => to_unsigned(85, 10), 659 => to_unsigned(1, 10), 660 => to_unsigned(271, 10), 661 => to_unsigned(454, 10), 662 => to_unsigned(879, 10), 663 => to_unsigned(394, 10), 664 => to_unsigned(954, 10), 665 => to_unsigned(713, 10), 666 => to_unsigned(936, 10), 667 => to_unsigned(630, 10), 668 => to_unsigned(56, 10), 669 => to_unsigned(845, 10), 670 => to_unsigned(70, 10), 671 => to_unsigned(762, 10), 672 => to_unsigned(664, 10), 673 => to_unsigned(10, 10), 674 => to_unsigned(498, 10), 675 => to_unsigned(122, 10), 676 => to_unsigned(430, 10), 677 => to_unsigned(418, 10), 678 => to_unsigned(704, 10), 679 => to_unsigned(861, 10), 680 => to_unsigned(1009, 10), 681 => to_unsigned(541, 10), 682 => to_unsigned(629, 10), 683 => to_unsigned(459, 10), 684 => to_unsigned(473, 10), 685 => to_unsigned(92, 10), 686 => to_unsigned(664, 10), 687 => to_unsigned(975, 10), 688 => to_unsigned(808, 10), 689 => to_unsigned(798, 10), 690 => to_unsigned(240, 10), 691 => to_unsigned(736, 10), 692 => to_unsigned(124, 10), 693 => to_unsigned(551, 10), 694 => to_unsigned(491, 10), 695 => to_unsigned(957, 10), 696 => to_unsigned(865, 10), 697 => to_unsigned(353, 10), 698 => to_unsigned(861, 10), 699 => to_unsigned(495, 10), 700 => to_unsigned(399, 10), 701 => to_unsigned(885, 10), 702 => to_unsigned(526, 10), 703 => to_unsigned(442, 10), 704 => to_unsigned(246, 10), 705 => to_unsigned(439, 10), 706 => to_unsigned(972, 10), 707 => to_unsigned(277, 10), 708 => to_unsigned(573, 10), 709 => to_unsigned(132, 10), 710 => to_unsigned(897, 10), 711 => to_unsigned(979, 10), 712 => to_unsigned(656, 10), 713 => to_unsigned(279, 10), 714 => to_unsigned(1010, 10), 715 => to_unsigned(658, 10), 716 => to_unsigned(1019, 10), 717 => to_unsigned(684, 10), 718 => to_unsigned(920, 10), 719 => to_unsigned(600, 10), 720 => to_unsigned(208, 10), 721 => to_unsigned(671, 10), 722 => to_unsigned(160, 10), 723 => to_unsigned(863, 10), 724 => to_unsigned(847, 10), 725 => to_unsigned(404, 10), 726 => to_unsigned(36, 10), 727 => to_unsigned(56, 10), 728 => to_unsigned(926, 10), 729 => to_unsigned(232, 10), 730 => to_unsigned(989, 10), 731 => to_unsigned(747, 10), 732 => to_unsigned(885, 10), 733 => to_unsigned(432, 10), 734 => to_unsigned(414, 10), 735 => to_unsigned(340, 10), 736 => to_unsigned(176, 10), 737 => to_unsigned(496, 10), 738 => to_unsigned(307, 10), 739 => to_unsigned(49, 10), 740 => to_unsigned(220, 10), 741 => to_unsigned(760, 10), 742 => to_unsigned(730, 10), 743 => to_unsigned(465, 10), 744 => to_unsigned(70, 10), 745 => to_unsigned(541, 10), 746 => to_unsigned(947, 10), 747 => to_unsigned(897, 10), 748 => to_unsigned(6, 10), 749 => to_unsigned(950, 10), 750 => to_unsigned(821, 10), 751 => to_unsigned(117, 10), 752 => to_unsigned(557, 10), 753 => to_unsigned(503, 10), 754 => to_unsigned(385, 10), 755 => to_unsigned(852, 10), 756 => to_unsigned(701, 10), 757 => to_unsigned(733, 10), 758 => to_unsigned(881, 10), 759 => to_unsigned(233, 10), 760 => to_unsigned(498, 10), 761 => to_unsigned(145, 10), 762 => to_unsigned(541, 10), 763 => to_unsigned(614, 10), 764 => to_unsigned(119, 10), 765 => to_unsigned(699, 10), 766 => to_unsigned(327, 10), 767 => to_unsigned(212, 10), 768 => to_unsigned(987, 10), 769 => to_unsigned(217, 10), 770 => to_unsigned(776, 10), 771 => to_unsigned(204, 10), 772 => to_unsigned(983, 10), 773 => to_unsigned(197, 10), 774 => to_unsigned(509, 10), 775 => to_unsigned(478, 10), 776 => to_unsigned(291, 10), 777 => to_unsigned(539, 10), 778 => to_unsigned(249, 10), 779 => to_unsigned(221, 10), 780 => to_unsigned(495, 10), 781 => to_unsigned(732, 10), 782 => to_unsigned(280, 10), 783 => to_unsigned(458, 10), 784 => to_unsigned(919, 10), 785 => to_unsigned(468, 10), 786 => to_unsigned(764, 10), 787 => to_unsigned(641, 10), 788 => to_unsigned(743, 10), 789 => to_unsigned(262, 10), 790 => to_unsigned(117, 10), 791 => to_unsigned(866, 10), 792 => to_unsigned(217, 10), 793 => to_unsigned(798, 10), 794 => to_unsigned(654, 10), 795 => to_unsigned(364, 10), 796 => to_unsigned(39, 10), 797 => to_unsigned(874, 10), 798 => to_unsigned(926, 10), 799 => to_unsigned(146, 10), 800 => to_unsigned(2, 10), 801 => to_unsigned(147, 10), 802 => to_unsigned(247, 10), 803 => to_unsigned(249, 10), 804 => to_unsigned(829, 10), 805 => to_unsigned(864, 10), 806 => to_unsigned(16, 10), 807 => to_unsigned(743, 10), 808 => to_unsigned(570, 10), 809 => to_unsigned(741, 10), 810 => to_unsigned(40, 10), 811 => to_unsigned(995, 10), 812 => to_unsigned(970, 10), 813 => to_unsigned(47, 10), 814 => to_unsigned(97, 10), 815 => to_unsigned(579, 10), 816 => to_unsigned(853, 10), 817 => to_unsigned(141, 10), 818 => to_unsigned(232, 10), 819 => to_unsigned(292, 10), 820 => to_unsigned(350, 10), 821 => to_unsigned(427, 10), 822 => to_unsigned(593, 10), 823 => to_unsigned(637, 10), 824 => to_unsigned(762, 10), 825 => to_unsigned(169, 10), 826 => to_unsigned(28, 10), 827 => to_unsigned(876, 10), 828 => to_unsigned(546, 10), 829 => to_unsigned(826, 10), 830 => to_unsigned(506, 10), 831 => to_unsigned(462, 10), 832 => to_unsigned(892, 10), 833 => to_unsigned(710, 10), 834 => to_unsigned(983, 10), 835 => to_unsigned(895, 10), 836 => to_unsigned(793, 10), 837 => to_unsigned(796, 10), 838 => to_unsigned(1012, 10), 839 => to_unsigned(163, 10), 840 => to_unsigned(709, 10), 841 => to_unsigned(511, 10), 842 => to_unsigned(757, 10), 843 => to_unsigned(745, 10), 844 => to_unsigned(768, 10), 845 => to_unsigned(388, 10), 846 => to_unsigned(836, 10), 847 => to_unsigned(483, 10), 848 => to_unsigned(713, 10), 849 => to_unsigned(156, 10), 850 => to_unsigned(237, 10), 851 => to_unsigned(514, 10), 852 => to_unsigned(690, 10), 853 => to_unsigned(686, 10), 854 => to_unsigned(914, 10), 855 => to_unsigned(727, 10), 856 => to_unsigned(881, 10), 857 => to_unsigned(375, 10), 858 => to_unsigned(87, 10), 859 => to_unsigned(37, 10), 860 => to_unsigned(815, 10), 861 => to_unsigned(997, 10), 862 => to_unsigned(934, 10), 863 => to_unsigned(48, 10), 864 => to_unsigned(478, 10), 865 => to_unsigned(944, 10), 866 => to_unsigned(261, 10), 867 => to_unsigned(837, 10), 868 => to_unsigned(514, 10), 869 => to_unsigned(402, 10), 870 => to_unsigned(19, 10), 871 => to_unsigned(743, 10), 872 => to_unsigned(28, 10), 873 => to_unsigned(1006, 10), 874 => to_unsigned(265, 10), 875 => to_unsigned(1018, 10), 876 => to_unsigned(334, 10), 877 => to_unsigned(704, 10), 878 => to_unsigned(779, 10), 879 => to_unsigned(137, 10), 880 => to_unsigned(190, 10), 881 => to_unsigned(435, 10), 882 => to_unsigned(731, 10), 883 => to_unsigned(459, 10), 884 => to_unsigned(450, 10), 885 => to_unsigned(483, 10), 886 => to_unsigned(716, 10), 887 => to_unsigned(146, 10), 888 => to_unsigned(135, 10), 889 => to_unsigned(65, 10), 890 => to_unsigned(889, 10), 891 => to_unsigned(286, 10), 892 => to_unsigned(903, 10), 893 => to_unsigned(78, 10), 894 => to_unsigned(160, 10), 895 => to_unsigned(871, 10), 896 => to_unsigned(353, 10), 897 => to_unsigned(714, 10), 898 => to_unsigned(860, 10), 899 => to_unsigned(999, 10), 900 => to_unsigned(17, 10), 901 => to_unsigned(258, 10), 902 => to_unsigned(119, 10), 903 => to_unsigned(407, 10), 904 => to_unsigned(804, 10), 905 => to_unsigned(362, 10), 906 => to_unsigned(847, 10), 907 => to_unsigned(262, 10), 908 => to_unsigned(662, 10), 909 => to_unsigned(461, 10), 910 => to_unsigned(890, 10), 911 => to_unsigned(216, 10), 912 => to_unsigned(191, 10), 913 => to_unsigned(825, 10), 914 => to_unsigned(90, 10), 915 => to_unsigned(252, 10), 916 => to_unsigned(287, 10), 917 => to_unsigned(277, 10), 918 => to_unsigned(520, 10), 919 => to_unsigned(232, 10), 920 => to_unsigned(69, 10), 921 => to_unsigned(246, 10), 922 => to_unsigned(537, 10), 923 => to_unsigned(59, 10), 924 => to_unsigned(585, 10), 925 => to_unsigned(1009, 10), 926 => to_unsigned(906, 10), 927 => to_unsigned(527, 10), 928 => to_unsigned(935, 10), 929 => to_unsigned(798, 10), 930 => to_unsigned(964, 10), 931 => to_unsigned(744, 10), 932 => to_unsigned(780, 10), 933 => to_unsigned(499, 10), 934 => to_unsigned(837, 10), 935 => to_unsigned(744, 10), 936 => to_unsigned(520, 10), 937 => to_unsigned(861, 10), 938 => to_unsigned(593, 10), 939 => to_unsigned(397, 10), 940 => to_unsigned(970, 10), 941 => to_unsigned(525, 10), 942 => to_unsigned(259, 10), 943 => to_unsigned(684, 10), 944 => to_unsigned(327, 10), 945 => to_unsigned(842, 10), 946 => to_unsigned(604, 10), 947 => to_unsigned(946, 10), 948 => to_unsigned(669, 10), 949 => to_unsigned(339, 10), 950 => to_unsigned(402, 10), 951 => to_unsigned(544, 10), 952 => to_unsigned(739, 10), 953 => to_unsigned(500, 10), 954 => to_unsigned(57, 10), 955 => to_unsigned(722, 10), 956 => to_unsigned(259, 10), 957 => to_unsigned(211, 10), 958 => to_unsigned(684, 10), 959 => to_unsigned(242, 10), 960 => to_unsigned(641, 10), 961 => to_unsigned(283, 10), 962 => to_unsigned(859, 10), 963 => to_unsigned(280, 10), 964 => to_unsigned(308, 10), 965 => to_unsigned(931, 10), 966 => to_unsigned(733, 10), 967 => to_unsigned(40, 10), 968 => to_unsigned(83, 10), 969 => to_unsigned(19, 10), 970 => to_unsigned(634, 10), 971 => to_unsigned(156, 10), 972 => to_unsigned(140, 10), 973 => to_unsigned(46, 10), 974 => to_unsigned(221, 10), 975 => to_unsigned(68, 10), 976 => to_unsigned(155, 10), 977 => to_unsigned(118, 10), 978 => to_unsigned(829, 10), 979 => to_unsigned(987, 10), 980 => to_unsigned(300, 10), 981 => to_unsigned(720, 10), 982 => to_unsigned(88, 10), 983 => to_unsigned(169, 10), 984 => to_unsigned(837, 10), 985 => to_unsigned(605, 10), 986 => to_unsigned(966, 10), 987 => to_unsigned(264, 10), 988 => to_unsigned(374, 10), 989 => to_unsigned(995, 10), 990 => to_unsigned(1007, 10), 991 => to_unsigned(446, 10), 992 => to_unsigned(393, 10), 993 => to_unsigned(163, 10), 994 => to_unsigned(589, 10), 995 => to_unsigned(154, 10), 996 => to_unsigned(712, 10), 997 => to_unsigned(828, 10), 998 => to_unsigned(637, 10), 999 => to_unsigned(996, 10), 1000 => to_unsigned(903, 10), 1001 => to_unsigned(42, 10), 1002 => to_unsigned(674, 10), 1003 => to_unsigned(111, 10), 1004 => to_unsigned(987, 10), 1005 => to_unsigned(311, 10), 1006 => to_unsigned(1012, 10), 1007 => to_unsigned(590, 10), 1008 => to_unsigned(407, 10), 1009 => to_unsigned(985, 10), 1010 => to_unsigned(293, 10), 1011 => to_unsigned(712, 10), 1012 => to_unsigned(341, 10), 1013 => to_unsigned(804, 10), 1014 => to_unsigned(663, 10), 1015 => to_unsigned(487, 10), 1016 => to_unsigned(925, 10), 1017 => to_unsigned(140, 10), 1018 => to_unsigned(320, 10), 1019 => to_unsigned(998, 10), 1020 => to_unsigned(552, 10), 1021 => to_unsigned(120, 10), 1022 => to_unsigned(93, 10), 1023 => to_unsigned(771, 10), 1024 => to_unsigned(1023, 10), 1025 => to_unsigned(583, 10), 1026 => to_unsigned(418, 10), 1027 => to_unsigned(191, 10), 1028 => to_unsigned(647, 10), 1029 => to_unsigned(436, 10), 1030 => to_unsigned(629, 10), 1031 => to_unsigned(528, 10), 1032 => to_unsigned(114, 10), 1033 => to_unsigned(592, 10), 1034 => to_unsigned(289, 10), 1035 => to_unsigned(298, 10), 1036 => to_unsigned(290, 10), 1037 => to_unsigned(254, 10), 1038 => to_unsigned(256, 10), 1039 => to_unsigned(974, 10), 1040 => to_unsigned(559, 10), 1041 => to_unsigned(38, 10), 1042 => to_unsigned(256, 10), 1043 => to_unsigned(137, 10), 1044 => to_unsigned(123, 10), 1045 => to_unsigned(497, 10), 1046 => to_unsigned(265, 10), 1047 => to_unsigned(682, 10), 1048 => to_unsigned(640, 10), 1049 => to_unsigned(632, 10), 1050 => to_unsigned(574, 10), 1051 => to_unsigned(823, 10), 1052 => to_unsigned(386, 10), 1053 => to_unsigned(972, 10), 1054 => to_unsigned(670, 10), 1055 => to_unsigned(44, 10), 1056 => to_unsigned(206, 10), 1057 => to_unsigned(669, 10), 1058 => to_unsigned(771, 10), 1059 => to_unsigned(420, 10), 1060 => to_unsigned(428, 10), 1061 => to_unsigned(84, 10), 1062 => to_unsigned(872, 10), 1063 => to_unsigned(203, 10), 1064 => to_unsigned(1015, 10), 1065 => to_unsigned(396, 10), 1066 => to_unsigned(723, 10), 1067 => to_unsigned(383, 10), 1068 => to_unsigned(458, 10), 1069 => to_unsigned(412, 10), 1070 => to_unsigned(962, 10), 1071 => to_unsigned(540, 10), 1072 => to_unsigned(602, 10), 1073 => to_unsigned(190, 10), 1074 => to_unsigned(893, 10), 1075 => to_unsigned(397, 10), 1076 => to_unsigned(7, 10), 1077 => to_unsigned(736, 10), 1078 => to_unsigned(481, 10), 1079 => to_unsigned(252, 10), 1080 => to_unsigned(452, 10), 1081 => to_unsigned(818, 10), 1082 => to_unsigned(113, 10), 1083 => to_unsigned(514, 10), 1084 => to_unsigned(193, 10), 1085 => to_unsigned(497, 10), 1086 => to_unsigned(954, 10), 1087 => to_unsigned(947, 10), 1088 => to_unsigned(296, 10), 1089 => to_unsigned(767, 10), 1090 => to_unsigned(577, 10), 1091 => to_unsigned(95, 10), 1092 => to_unsigned(528, 10), 1093 => to_unsigned(471, 10), 1094 => to_unsigned(383, 10), 1095 => to_unsigned(604, 10), 1096 => to_unsigned(413, 10), 1097 => to_unsigned(554, 10), 1098 => to_unsigned(777, 10), 1099 => to_unsigned(473, 10), 1100 => to_unsigned(363, 10), 1101 => to_unsigned(628, 10), 1102 => to_unsigned(616, 10), 1103 => to_unsigned(377, 10), 1104 => to_unsigned(839, 10), 1105 => to_unsigned(996, 10), 1106 => to_unsigned(882, 10), 1107 => to_unsigned(294, 10), 1108 => to_unsigned(335, 10), 1109 => to_unsigned(657, 10), 1110 => to_unsigned(681, 10), 1111 => to_unsigned(703, 10), 1112 => to_unsigned(274, 10), 1113 => to_unsigned(139, 10), 1114 => to_unsigned(383, 10), 1115 => to_unsigned(474, 10), 1116 => to_unsigned(684, 10), 1117 => to_unsigned(437, 10), 1118 => to_unsigned(213, 10), 1119 => to_unsigned(361, 10), 1120 => to_unsigned(353, 10), 1121 => to_unsigned(869, 10), 1122 => to_unsigned(662, 10), 1123 => to_unsigned(623, 10), 1124 => to_unsigned(535, 10), 1125 => to_unsigned(491, 10), 1126 => to_unsigned(658, 10), 1127 => to_unsigned(837, 10), 1128 => to_unsigned(249, 10), 1129 => to_unsigned(898, 10), 1130 => to_unsigned(179, 10), 1131 => to_unsigned(117, 10), 1132 => to_unsigned(884, 10), 1133 => to_unsigned(430, 10), 1134 => to_unsigned(89, 10), 1135 => to_unsigned(851, 10), 1136 => to_unsigned(485, 10), 1137 => to_unsigned(73, 10), 1138 => to_unsigned(152, 10), 1139 => to_unsigned(546, 10), 1140 => to_unsigned(944, 10), 1141 => to_unsigned(703, 10), 1142 => to_unsigned(727, 10), 1143 => to_unsigned(212, 10), 1144 => to_unsigned(353, 10), 1145 => to_unsigned(721, 10), 1146 => to_unsigned(246, 10), 1147 => to_unsigned(210, 10), 1148 => to_unsigned(706, 10), 1149 => to_unsigned(709, 10), 1150 => to_unsigned(979, 10), 1151 => to_unsigned(55, 10), 1152 => to_unsigned(341, 10), 1153 => to_unsigned(177, 10), 1154 => to_unsigned(502, 10), 1155 => to_unsigned(608, 10), 1156 => to_unsigned(589, 10), 1157 => to_unsigned(694, 10), 1158 => to_unsigned(107, 10), 1159 => to_unsigned(584, 10), 1160 => to_unsigned(44, 10), 1161 => to_unsigned(383, 10), 1162 => to_unsigned(856, 10), 1163 => to_unsigned(750, 10), 1164 => to_unsigned(399, 10), 1165 => to_unsigned(646, 10), 1166 => to_unsigned(693, 10), 1167 => to_unsigned(138, 10), 1168 => to_unsigned(986, 10), 1169 => to_unsigned(887, 10), 1170 => to_unsigned(487, 10), 1171 => to_unsigned(464, 10), 1172 => to_unsigned(964, 10), 1173 => to_unsigned(604, 10), 1174 => to_unsigned(137, 10), 1175 => to_unsigned(757, 10), 1176 => to_unsigned(110, 10), 1177 => to_unsigned(312, 10), 1178 => to_unsigned(308, 10), 1179 => to_unsigned(216, 10), 1180 => to_unsigned(407, 10), 1181 => to_unsigned(555, 10), 1182 => to_unsigned(139, 10), 1183 => to_unsigned(708, 10), 1184 => to_unsigned(244, 10), 1185 => to_unsigned(796, 10), 1186 => to_unsigned(866, 10), 1187 => to_unsigned(406, 10), 1188 => to_unsigned(223, 10), 1189 => to_unsigned(551, 10), 1190 => to_unsigned(978, 10), 1191 => to_unsigned(856, 10), 1192 => to_unsigned(508, 10), 1193 => to_unsigned(172, 10), 1194 => to_unsigned(932, 10), 1195 => to_unsigned(960, 10), 1196 => to_unsigned(1002, 10), 1197 => to_unsigned(636, 10), 1198 => to_unsigned(908, 10), 1199 => to_unsigned(331, 10), 1200 => to_unsigned(110, 10), 1201 => to_unsigned(618, 10), 1202 => to_unsigned(760, 10), 1203 => to_unsigned(952, 10), 1204 => to_unsigned(380, 10), 1205 => to_unsigned(996, 10), 1206 => to_unsigned(105, 10), 1207 => to_unsigned(168, 10), 1208 => to_unsigned(587, 10), 1209 => to_unsigned(227, 10), 1210 => to_unsigned(741, 10), 1211 => to_unsigned(371, 10), 1212 => to_unsigned(520, 10), 1213 => to_unsigned(653, 10), 1214 => to_unsigned(236, 10), 1215 => to_unsigned(34, 10), 1216 => to_unsigned(799, 10), 1217 => to_unsigned(45, 10), 1218 => to_unsigned(66, 10), 1219 => to_unsigned(797, 10), 1220 => to_unsigned(880, 10), 1221 => to_unsigned(198, 10), 1222 => to_unsigned(889, 10), 1223 => to_unsigned(832, 10), 1224 => to_unsigned(1021, 10), 1225 => to_unsigned(1021, 10), 1226 => to_unsigned(497, 10), 1227 => to_unsigned(575, 10), 1228 => to_unsigned(211, 10), 1229 => to_unsigned(792, 10), 1230 => to_unsigned(507, 10), 1231 => to_unsigned(928, 10), 1232 => to_unsigned(546, 10), 1233 => to_unsigned(123, 10), 1234 => to_unsigned(315, 10), 1235 => to_unsigned(380, 10), 1236 => to_unsigned(950, 10), 1237 => to_unsigned(683, 10), 1238 => to_unsigned(727, 10), 1239 => to_unsigned(77, 10), 1240 => to_unsigned(678, 10), 1241 => to_unsigned(427, 10), 1242 => to_unsigned(244, 10), 1243 => to_unsigned(632, 10), 1244 => to_unsigned(929, 10), 1245 => to_unsigned(17, 10), 1246 => to_unsigned(769, 10), 1247 => to_unsigned(933, 10), 1248 => to_unsigned(829, 10), 1249 => to_unsigned(976, 10), 1250 => to_unsigned(598, 10), 1251 => to_unsigned(121, 10), 1252 => to_unsigned(690, 10), 1253 => to_unsigned(224, 10), 1254 => to_unsigned(731, 10), 1255 => to_unsigned(142, 10), 1256 => to_unsigned(586, 10), 1257 => to_unsigned(150, 10), 1258 => to_unsigned(140, 10), 1259 => to_unsigned(316, 10), 1260 => to_unsigned(110, 10), 1261 => to_unsigned(74, 10), 1262 => to_unsigned(291, 10), 1263 => to_unsigned(101, 10), 1264 => to_unsigned(474, 10), 1265 => to_unsigned(209, 10), 1266 => to_unsigned(935, 10), 1267 => to_unsigned(255, 10), 1268 => to_unsigned(549, 10), 1269 => to_unsigned(225, 10), 1270 => to_unsigned(533, 10), 1271 => to_unsigned(721, 10), 1272 => to_unsigned(437, 10), 1273 => to_unsigned(104, 10), 1274 => to_unsigned(627, 10), 1275 => to_unsigned(337, 10), 1276 => to_unsigned(140, 10), 1277 => to_unsigned(998, 10), 1278 => to_unsigned(847, 10), 1279 => to_unsigned(519, 10), 1280 => to_unsigned(289, 10), 1281 => to_unsigned(1023, 10), 1282 => to_unsigned(540, 10), 1283 => to_unsigned(261, 10), 1284 => to_unsigned(549, 10), 1285 => to_unsigned(611, 10), 1286 => to_unsigned(175, 10), 1287 => to_unsigned(62, 10), 1288 => to_unsigned(233, 10), 1289 => to_unsigned(921, 10), 1290 => to_unsigned(273, 10), 1291 => to_unsigned(266, 10), 1292 => to_unsigned(538, 10), 1293 => to_unsigned(541, 10), 1294 => to_unsigned(657, 10), 1295 => to_unsigned(874, 10), 1296 => to_unsigned(67, 10), 1297 => to_unsigned(261, 10), 1298 => to_unsigned(213, 10), 1299 => to_unsigned(833, 10), 1300 => to_unsigned(179, 10), 1301 => to_unsigned(878, 10), 1302 => to_unsigned(1007, 10), 1303 => to_unsigned(167, 10), 1304 => to_unsigned(351, 10), 1305 => to_unsigned(1016, 10), 1306 => to_unsigned(486, 10), 1307 => to_unsigned(433, 10), 1308 => to_unsigned(148, 10), 1309 => to_unsigned(519, 10), 1310 => to_unsigned(88, 10), 1311 => to_unsigned(360, 10), 1312 => to_unsigned(739, 10), 1313 => to_unsigned(451, 10), 1314 => to_unsigned(567, 10), 1315 => to_unsigned(334, 10), 1316 => to_unsigned(795, 10), 1317 => to_unsigned(19, 10), 1318 => to_unsigned(229, 10), 1319 => to_unsigned(69, 10), 1320 => to_unsigned(157, 10), 1321 => to_unsigned(574, 10), 1322 => to_unsigned(351, 10), 1323 => to_unsigned(176, 10), 1324 => to_unsigned(488, 10), 1325 => to_unsigned(835, 10), 1326 => to_unsigned(60, 10), 1327 => to_unsigned(34, 10), 1328 => to_unsigned(29, 10), 1329 => to_unsigned(560, 10), 1330 => to_unsigned(936, 10), 1331 => to_unsigned(307, 10), 1332 => to_unsigned(725, 10), 1333 => to_unsigned(1, 10), 1334 => to_unsigned(369, 10), 1335 => to_unsigned(820, 10), 1336 => to_unsigned(459, 10), 1337 => to_unsigned(993, 10), 1338 => to_unsigned(993, 10), 1339 => to_unsigned(717, 10), 1340 => to_unsigned(38, 10), 1341 => to_unsigned(742, 10), 1342 => to_unsigned(236, 10), 1343 => to_unsigned(5, 10), 1344 => to_unsigned(903, 10), 1345 => to_unsigned(794, 10), 1346 => to_unsigned(459, 10), 1347 => to_unsigned(497, 10), 1348 => to_unsigned(596, 10), 1349 => to_unsigned(503, 10), 1350 => to_unsigned(485, 10), 1351 => to_unsigned(515, 10), 1352 => to_unsigned(88, 10), 1353 => to_unsigned(888, 10), 1354 => to_unsigned(170, 10), 1355 => to_unsigned(343, 10), 1356 => to_unsigned(139, 10), 1357 => to_unsigned(58, 10), 1358 => to_unsigned(796, 10), 1359 => to_unsigned(354, 10), 1360 => to_unsigned(702, 10), 1361 => to_unsigned(569, 10), 1362 => to_unsigned(356, 10), 1363 => to_unsigned(797, 10), 1364 => to_unsigned(872, 10), 1365 => to_unsigned(571, 10), 1366 => to_unsigned(425, 10), 1367 => to_unsigned(290, 10), 1368 => to_unsigned(0, 10), 1369 => to_unsigned(39, 10), 1370 => to_unsigned(601, 10), 1371 => to_unsigned(508, 10), 1372 => to_unsigned(930, 10), 1373 => to_unsigned(564, 10), 1374 => to_unsigned(489, 10), 1375 => to_unsigned(454, 10), 1376 => to_unsigned(771, 10), 1377 => to_unsigned(196, 10), 1378 => to_unsigned(251, 10), 1379 => to_unsigned(806, 10), 1380 => to_unsigned(138, 10), 1381 => to_unsigned(398, 10), 1382 => to_unsigned(95, 10), 1383 => to_unsigned(369, 10), 1384 => to_unsigned(676, 10), 1385 => to_unsigned(840, 10), 1386 => to_unsigned(238, 10), 1387 => to_unsigned(927, 10), 1388 => to_unsigned(96, 10), 1389 => to_unsigned(57, 10), 1390 => to_unsigned(470, 10), 1391 => to_unsigned(782, 10), 1392 => to_unsigned(541, 10), 1393 => to_unsigned(15, 10), 1394 => to_unsigned(498, 10), 1395 => to_unsigned(533, 10), 1396 => to_unsigned(938, 10), 1397 => to_unsigned(157, 10), 1398 => to_unsigned(0, 10), 1399 => to_unsigned(610, 10), 1400 => to_unsigned(435, 10), 1401 => to_unsigned(337, 10), 1402 => to_unsigned(78, 10), 1403 => to_unsigned(1009, 10), 1404 => to_unsigned(444, 10), 1405 => to_unsigned(660, 10), 1406 => to_unsigned(935, 10), 1407 => to_unsigned(257, 10), 1408 => to_unsigned(605, 10), 1409 => to_unsigned(615, 10), 1410 => to_unsigned(671, 10), 1411 => to_unsigned(667, 10), 1412 => to_unsigned(970, 10), 1413 => to_unsigned(63, 10), 1414 => to_unsigned(582, 10), 1415 => to_unsigned(704, 10), 1416 => to_unsigned(42, 10), 1417 => to_unsigned(283, 10), 1418 => to_unsigned(102, 10), 1419 => to_unsigned(146, 10), 1420 => to_unsigned(562, 10), 1421 => to_unsigned(166, 10), 1422 => to_unsigned(543, 10), 1423 => to_unsigned(306, 10), 1424 => to_unsigned(1008, 10), 1425 => to_unsigned(437, 10), 1426 => to_unsigned(52, 10), 1427 => to_unsigned(349, 10), 1428 => to_unsigned(449, 10), 1429 => to_unsigned(683, 10), 1430 => to_unsigned(426, 10), 1431 => to_unsigned(932, 10), 1432 => to_unsigned(210, 10), 1433 => to_unsigned(153, 10), 1434 => to_unsigned(1013, 10), 1435 => to_unsigned(318, 10), 1436 => to_unsigned(64, 10), 1437 => to_unsigned(169, 10), 1438 => to_unsigned(347, 10), 1439 => to_unsigned(374, 10), 1440 => to_unsigned(954, 10), 1441 => to_unsigned(89, 10), 1442 => to_unsigned(103, 10), 1443 => to_unsigned(802, 10), 1444 => to_unsigned(386, 10), 1445 => to_unsigned(760, 10), 1446 => to_unsigned(921, 10), 1447 => to_unsigned(32, 10), 1448 => to_unsigned(955, 10), 1449 => to_unsigned(725, 10), 1450 => to_unsigned(637, 10), 1451 => to_unsigned(901, 10), 1452 => to_unsigned(297, 10), 1453 => to_unsigned(481, 10), 1454 => to_unsigned(706, 10), 1455 => to_unsigned(248, 10), 1456 => to_unsigned(848, 10), 1457 => to_unsigned(773, 10), 1458 => to_unsigned(809, 10), 1459 => to_unsigned(635, 10), 1460 => to_unsigned(772, 10), 1461 => to_unsigned(19, 10), 1462 => to_unsigned(704, 10), 1463 => to_unsigned(56, 10), 1464 => to_unsigned(599, 10), 1465 => to_unsigned(456, 10), 1466 => to_unsigned(398, 10), 1467 => to_unsigned(890, 10), 1468 => to_unsigned(702, 10), 1469 => to_unsigned(822, 10), 1470 => to_unsigned(932, 10), 1471 => to_unsigned(593, 10), 1472 => to_unsigned(697, 10), 1473 => to_unsigned(505, 10), 1474 => to_unsigned(533, 10), 1475 => to_unsigned(714, 10), 1476 => to_unsigned(997, 10), 1477 => to_unsigned(898, 10), 1478 => to_unsigned(540, 10), 1479 => to_unsigned(1012, 10), 1480 => to_unsigned(621, 10), 1481 => to_unsigned(927, 10), 1482 => to_unsigned(417, 10), 1483 => to_unsigned(377, 10), 1484 => to_unsigned(71, 10), 1485 => to_unsigned(865, 10), 1486 => to_unsigned(196, 10), 1487 => to_unsigned(520, 10), 1488 => to_unsigned(464, 10), 1489 => to_unsigned(467, 10), 1490 => to_unsigned(41, 10), 1491 => to_unsigned(474, 10), 1492 => to_unsigned(374, 10), 1493 => to_unsigned(324, 10), 1494 => to_unsigned(45, 10), 1495 => to_unsigned(188, 10), 1496 => to_unsigned(540, 10), 1497 => to_unsigned(778, 10), 1498 => to_unsigned(25, 10), 1499 => to_unsigned(121, 10), 1500 => to_unsigned(214, 10), 1501 => to_unsigned(337, 10), 1502 => to_unsigned(113, 10), 1503 => to_unsigned(339, 10), 1504 => to_unsigned(811, 10), 1505 => to_unsigned(1019, 10), 1506 => to_unsigned(691, 10), 1507 => to_unsigned(660, 10), 1508 => to_unsigned(985, 10), 1509 => to_unsigned(287, 10), 1510 => to_unsigned(576, 10), 1511 => to_unsigned(577, 10), 1512 => to_unsigned(116, 10), 1513 => to_unsigned(963, 10), 1514 => to_unsigned(424, 10), 1515 => to_unsigned(9, 10), 1516 => to_unsigned(440, 10), 1517 => to_unsigned(475, 10), 1518 => to_unsigned(880, 10), 1519 => to_unsigned(868, 10), 1520 => to_unsigned(592, 10), 1521 => to_unsigned(925, 10), 1522 => to_unsigned(517, 10), 1523 => to_unsigned(10, 10), 1524 => to_unsigned(567, 10), 1525 => to_unsigned(778, 10), 1526 => to_unsigned(513, 10), 1527 => to_unsigned(403, 10), 1528 => to_unsigned(289, 10), 1529 => to_unsigned(377, 10), 1530 => to_unsigned(296, 10), 1531 => to_unsigned(576, 10), 1532 => to_unsigned(431, 10), 1533 => to_unsigned(26, 10), 1534 => to_unsigned(756, 10), 1535 => to_unsigned(436, 10), 1536 => to_unsigned(153, 10), 1537 => to_unsigned(563, 10), 1538 => to_unsigned(985, 10), 1539 => to_unsigned(711, 10), 1540 => to_unsigned(307, 10), 1541 => to_unsigned(156, 10), 1542 => to_unsigned(656, 10), 1543 => to_unsigned(288, 10), 1544 => to_unsigned(512, 10), 1545 => to_unsigned(407, 10), 1546 => to_unsigned(88, 10), 1547 => to_unsigned(694, 10), 1548 => to_unsigned(49, 10), 1549 => to_unsigned(247, 10), 1550 => to_unsigned(832, 10), 1551 => to_unsigned(473, 10), 1552 => to_unsigned(271, 10), 1553 => to_unsigned(304, 10), 1554 => to_unsigned(928, 10), 1555 => to_unsigned(315, 10), 1556 => to_unsigned(923, 10), 1557 => to_unsigned(812, 10), 1558 => to_unsigned(54, 10), 1559 => to_unsigned(535, 10), 1560 => to_unsigned(931, 10), 1561 => to_unsigned(589, 10), 1562 => to_unsigned(48, 10), 1563 => to_unsigned(260, 10), 1564 => to_unsigned(185, 10), 1565 => to_unsigned(378, 10), 1566 => to_unsigned(185, 10), 1567 => to_unsigned(90, 10), 1568 => to_unsigned(77, 10), 1569 => to_unsigned(632, 10), 1570 => to_unsigned(791, 10), 1571 => to_unsigned(301, 10), 1572 => to_unsigned(731, 10), 1573 => to_unsigned(327, 10), 1574 => to_unsigned(418, 10), 1575 => to_unsigned(110, 10), 1576 => to_unsigned(316, 10), 1577 => to_unsigned(575, 10), 1578 => to_unsigned(500, 10), 1579 => to_unsigned(354, 10), 1580 => to_unsigned(854, 10), 1581 => to_unsigned(191, 10), 1582 => to_unsigned(140, 10), 1583 => to_unsigned(750, 10), 1584 => to_unsigned(208, 10), 1585 => to_unsigned(734, 10), 1586 => to_unsigned(649, 10), 1587 => to_unsigned(291, 10), 1588 => to_unsigned(924, 10), 1589 => to_unsigned(655, 10), 1590 => to_unsigned(442, 10), 1591 => to_unsigned(571, 10), 1592 => to_unsigned(928, 10), 1593 => to_unsigned(829, 10), 1594 => to_unsigned(973, 10), 1595 => to_unsigned(646, 10), 1596 => to_unsigned(416, 10), 1597 => to_unsigned(706, 10), 1598 => to_unsigned(985, 10), 1599 => to_unsigned(422, 10), 1600 => to_unsigned(132, 10), 1601 => to_unsigned(126, 10), 1602 => to_unsigned(214, 10), 1603 => to_unsigned(121, 10), 1604 => to_unsigned(96, 10), 1605 => to_unsigned(93, 10), 1606 => to_unsigned(928, 10), 1607 => to_unsigned(426, 10), 1608 => to_unsigned(792, 10), 1609 => to_unsigned(725, 10), 1610 => to_unsigned(896, 10), 1611 => to_unsigned(585, 10), 1612 => to_unsigned(22, 10), 1613 => to_unsigned(992, 10), 1614 => to_unsigned(998, 10), 1615 => to_unsigned(411, 10), 1616 => to_unsigned(362, 10), 1617 => to_unsigned(379, 10), 1618 => to_unsigned(583, 10), 1619 => to_unsigned(886, 10), 1620 => to_unsigned(282, 10), 1621 => to_unsigned(250, 10), 1622 => to_unsigned(316, 10), 1623 => to_unsigned(900, 10), 1624 => to_unsigned(590, 10), 1625 => to_unsigned(439, 10), 1626 => to_unsigned(824, 10), 1627 => to_unsigned(495, 10), 1628 => to_unsigned(149, 10), 1629 => to_unsigned(951, 10), 1630 => to_unsigned(482, 10), 1631 => to_unsigned(371, 10), 1632 => to_unsigned(605, 10), 1633 => to_unsigned(623, 10), 1634 => to_unsigned(555, 10), 1635 => to_unsigned(309, 10), 1636 => to_unsigned(672, 10), 1637 => to_unsigned(861, 10), 1638 => to_unsigned(763, 10), 1639 => to_unsigned(547, 10), 1640 => to_unsigned(463, 10), 1641 => to_unsigned(37, 10), 1642 => to_unsigned(182, 10), 1643 => to_unsigned(726, 10), 1644 => to_unsigned(292, 10), 1645 => to_unsigned(548, 10), 1646 => to_unsigned(411, 10), 1647 => to_unsigned(973, 10), 1648 => to_unsigned(895, 10), 1649 => to_unsigned(762, 10), 1650 => to_unsigned(643, 10), 1651 => to_unsigned(166, 10), 1652 => to_unsigned(498, 10), 1653 => to_unsigned(928, 10), 1654 => to_unsigned(350, 10), 1655 => to_unsigned(716, 10), 1656 => to_unsigned(163, 10), 1657 => to_unsigned(201, 10), 1658 => to_unsigned(434, 10), 1659 => to_unsigned(686, 10), 1660 => to_unsigned(478, 10), 1661 => to_unsigned(116, 10), 1662 => to_unsigned(601, 10), 1663 => to_unsigned(375, 10), 1664 => to_unsigned(318, 10), 1665 => to_unsigned(781, 10), 1666 => to_unsigned(771, 10), 1667 => to_unsigned(32, 10), 1668 => to_unsigned(942, 10), 1669 => to_unsigned(588, 10), 1670 => to_unsigned(623, 10), 1671 => to_unsigned(183, 10), 1672 => to_unsigned(1000, 10), 1673 => to_unsigned(764, 10), 1674 => to_unsigned(892, 10), 1675 => to_unsigned(59, 10), 1676 => to_unsigned(433, 10), 1677 => to_unsigned(929, 10), 1678 => to_unsigned(426, 10), 1679 => to_unsigned(34, 10), 1680 => to_unsigned(347, 10), 1681 => to_unsigned(862, 10), 1682 => to_unsigned(29, 10), 1683 => to_unsigned(799, 10), 1684 => to_unsigned(588, 10), 1685 => to_unsigned(40, 10), 1686 => to_unsigned(353, 10), 1687 => to_unsigned(7, 10), 1688 => to_unsigned(425, 10), 1689 => to_unsigned(756, 10), 1690 => to_unsigned(536, 10), 1691 => to_unsigned(544, 10), 1692 => to_unsigned(905, 10), 1693 => to_unsigned(743, 10), 1694 => to_unsigned(673, 10), 1695 => to_unsigned(945, 10), 1696 => to_unsigned(747, 10), 1697 => to_unsigned(608, 10), 1698 => to_unsigned(324, 10), 1699 => to_unsigned(1004, 10), 1700 => to_unsigned(730, 10), 1701 => to_unsigned(327, 10), 1702 => to_unsigned(498, 10), 1703 => to_unsigned(947, 10), 1704 => to_unsigned(838, 10), 1705 => to_unsigned(405, 10), 1706 => to_unsigned(557, 10), 1707 => to_unsigned(155, 10), 1708 => to_unsigned(8, 10), 1709 => to_unsigned(317, 10), 1710 => to_unsigned(1020, 10), 1711 => to_unsigned(94, 10), 1712 => to_unsigned(515, 10), 1713 => to_unsigned(68, 10), 1714 => to_unsigned(780, 10), 1715 => to_unsigned(645, 10), 1716 => to_unsigned(181, 10), 1717 => to_unsigned(278, 10), 1718 => to_unsigned(501, 10), 1719 => to_unsigned(622, 10), 1720 => to_unsigned(34, 10), 1721 => to_unsigned(59, 10), 1722 => to_unsigned(289, 10), 1723 => to_unsigned(1020, 10), 1724 => to_unsigned(823, 10), 1725 => to_unsigned(310, 10), 1726 => to_unsigned(485, 10), 1727 => to_unsigned(545, 10), 1728 => to_unsigned(889, 10), 1729 => to_unsigned(458, 10), 1730 => to_unsigned(517, 10), 1731 => to_unsigned(123, 10), 1732 => to_unsigned(479, 10), 1733 => to_unsigned(820, 10), 1734 => to_unsigned(118, 10), 1735 => to_unsigned(866, 10), 1736 => to_unsigned(690, 10), 1737 => to_unsigned(993, 10), 1738 => to_unsigned(234, 10), 1739 => to_unsigned(187, 10), 1740 => to_unsigned(411, 10), 1741 => to_unsigned(4, 10), 1742 => to_unsigned(993, 10), 1743 => to_unsigned(608, 10), 1744 => to_unsigned(907, 10), 1745 => to_unsigned(49, 10), 1746 => to_unsigned(615, 10), 1747 => to_unsigned(505, 10), 1748 => to_unsigned(1003, 10), 1749 => to_unsigned(869, 10), 1750 => to_unsigned(1023, 10), 1751 => to_unsigned(747, 10), 1752 => to_unsigned(267, 10), 1753 => to_unsigned(548, 10), 1754 => to_unsigned(704, 10), 1755 => to_unsigned(871, 10), 1756 => to_unsigned(964, 10), 1757 => to_unsigned(641, 10), 1758 => to_unsigned(557, 10), 1759 => to_unsigned(1021, 10), 1760 => to_unsigned(152, 10), 1761 => to_unsigned(677, 10), 1762 => to_unsigned(856, 10), 1763 => to_unsigned(47, 10), 1764 => to_unsigned(277, 10), 1765 => to_unsigned(56, 10), 1766 => to_unsigned(630, 10), 1767 => to_unsigned(690, 10), 1768 => to_unsigned(256, 10), 1769 => to_unsigned(664, 10), 1770 => to_unsigned(736, 10), 1771 => to_unsigned(981, 10), 1772 => to_unsigned(158, 10), 1773 => to_unsigned(210, 10), 1774 => to_unsigned(571, 10), 1775 => to_unsigned(111, 10), 1776 => to_unsigned(700, 10), 1777 => to_unsigned(913, 10), 1778 => to_unsigned(704, 10), 1779 => to_unsigned(402, 10), 1780 => to_unsigned(1012, 10), 1781 => to_unsigned(698, 10), 1782 => to_unsigned(333, 10), 1783 => to_unsigned(842, 10), 1784 => to_unsigned(839, 10), 1785 => to_unsigned(849, 10), 1786 => to_unsigned(264, 10), 1787 => to_unsigned(554, 10), 1788 => to_unsigned(603, 10), 1789 => to_unsigned(74, 10), 1790 => to_unsigned(958, 10), 1791 => to_unsigned(48, 10), 1792 => to_unsigned(552, 10), 1793 => to_unsigned(541, 10), 1794 => to_unsigned(747, 10), 1795 => to_unsigned(26, 10), 1796 => to_unsigned(1022, 10), 1797 => to_unsigned(217, 10), 1798 => to_unsigned(880, 10), 1799 => to_unsigned(822, 10), 1800 => to_unsigned(715, 10), 1801 => to_unsigned(293, 10), 1802 => to_unsigned(666, 10), 1803 => to_unsigned(420, 10), 1804 => to_unsigned(144, 10), 1805 => to_unsigned(621, 10), 1806 => to_unsigned(200, 10), 1807 => to_unsigned(901, 10), 1808 => to_unsigned(460, 10), 1809 => to_unsigned(261, 10), 1810 => to_unsigned(165, 10), 1811 => to_unsigned(515, 10), 1812 => to_unsigned(378, 10), 1813 => to_unsigned(911, 10), 1814 => to_unsigned(951, 10), 1815 => to_unsigned(355, 10), 1816 => to_unsigned(362, 10), 1817 => to_unsigned(845, 10), 1818 => to_unsigned(412, 10), 1819 => to_unsigned(855, 10), 1820 => to_unsigned(565, 10), 1821 => to_unsigned(230, 10), 1822 => to_unsigned(761, 10), 1823 => to_unsigned(870, 10), 1824 => to_unsigned(108, 10), 1825 => to_unsigned(152, 10), 1826 => to_unsigned(183, 10), 1827 => to_unsigned(365, 10), 1828 => to_unsigned(557, 10), 1829 => to_unsigned(829, 10), 1830 => to_unsigned(578, 10), 1831 => to_unsigned(809, 10), 1832 => to_unsigned(50, 10), 1833 => to_unsigned(410, 10), 1834 => to_unsigned(331, 10), 1835 => to_unsigned(42, 10), 1836 => to_unsigned(769, 10), 1837 => to_unsigned(613, 10), 1838 => to_unsigned(89, 10), 1839 => to_unsigned(988, 10), 1840 => to_unsigned(703, 10), 1841 => to_unsigned(556, 10), 1842 => to_unsigned(184, 10), 1843 => to_unsigned(861, 10), 1844 => to_unsigned(805, 10), 1845 => to_unsigned(104, 10), 1846 => to_unsigned(863, 10), 1847 => to_unsigned(741, 10), 1848 => to_unsigned(821, 10), 1849 => to_unsigned(724, 10), 1850 => to_unsigned(575, 10), 1851 => to_unsigned(71, 10), 1852 => to_unsigned(5, 10), 1853 => to_unsigned(451, 10), 1854 => to_unsigned(272, 10), 1855 => to_unsigned(532, 10), 1856 => to_unsigned(451, 10), 1857 => to_unsigned(610, 10), 1858 => to_unsigned(378, 10), 1859 => to_unsigned(157, 10), 1860 => to_unsigned(379, 10), 1861 => to_unsigned(730, 10), 1862 => to_unsigned(843, 10), 1863 => to_unsigned(687, 10), 1864 => to_unsigned(891, 10), 1865 => to_unsigned(19, 10), 1866 => to_unsigned(999, 10), 1867 => to_unsigned(939, 10), 1868 => to_unsigned(379, 10), 1869 => to_unsigned(168, 10), 1870 => to_unsigned(160, 10), 1871 => to_unsigned(959, 10), 1872 => to_unsigned(757, 10), 1873 => to_unsigned(137, 10), 1874 => to_unsigned(692, 10), 1875 => to_unsigned(433, 10), 1876 => to_unsigned(836, 10), 1877 => to_unsigned(842, 10), 1878 => to_unsigned(980, 10), 1879 => to_unsigned(189, 10), 1880 => to_unsigned(851, 10), 1881 => to_unsigned(235, 10), 1882 => to_unsigned(968, 10), 1883 => to_unsigned(958, 10), 1884 => to_unsigned(413, 10), 1885 => to_unsigned(1007, 10), 1886 => to_unsigned(179, 10), 1887 => to_unsigned(67, 10), 1888 => to_unsigned(692, 10), 1889 => to_unsigned(776, 10), 1890 => to_unsigned(243, 10), 1891 => to_unsigned(679, 10), 1892 => to_unsigned(315, 10), 1893 => to_unsigned(893, 10), 1894 => to_unsigned(578, 10), 1895 => to_unsigned(59, 10), 1896 => to_unsigned(101, 10), 1897 => to_unsigned(408, 10), 1898 => to_unsigned(356, 10), 1899 => to_unsigned(29, 10), 1900 => to_unsigned(350, 10), 1901 => to_unsigned(336, 10), 1902 => to_unsigned(649, 10), 1903 => to_unsigned(391, 10), 1904 => to_unsigned(569, 10), 1905 => to_unsigned(497, 10), 1906 => to_unsigned(897, 10), 1907 => to_unsigned(223, 10), 1908 => to_unsigned(522, 10), 1909 => to_unsigned(393, 10), 1910 => to_unsigned(168, 10), 1911 => to_unsigned(31, 10), 1912 => to_unsigned(855, 10), 1913 => to_unsigned(134, 10), 1914 => to_unsigned(891, 10), 1915 => to_unsigned(860, 10), 1916 => to_unsigned(761, 10), 1917 => to_unsigned(641, 10), 1918 => to_unsigned(15, 10), 1919 => to_unsigned(862, 10), 1920 => to_unsigned(779, 10), 1921 => to_unsigned(116, 10), 1922 => to_unsigned(956, 10), 1923 => to_unsigned(223, 10), 1924 => to_unsigned(558, 10), 1925 => to_unsigned(693, 10), 1926 => to_unsigned(232, 10), 1927 => to_unsigned(593, 10), 1928 => to_unsigned(322, 10), 1929 => to_unsigned(911, 10), 1930 => to_unsigned(48, 10), 1931 => to_unsigned(489, 10), 1932 => to_unsigned(977, 10), 1933 => to_unsigned(754, 10), 1934 => to_unsigned(171, 10), 1935 => to_unsigned(893, 10), 1936 => to_unsigned(692, 10), 1937 => to_unsigned(910, 10), 1938 => to_unsigned(552, 10), 1939 => to_unsigned(699, 10), 1940 => to_unsigned(484, 10), 1941 => to_unsigned(86, 10), 1942 => to_unsigned(573, 10), 1943 => to_unsigned(409, 10), 1944 => to_unsigned(70, 10), 1945 => to_unsigned(950, 10), 1946 => to_unsigned(495, 10), 1947 => to_unsigned(823, 10), 1948 => to_unsigned(113, 10), 1949 => to_unsigned(148, 10), 1950 => to_unsigned(732, 10), 1951 => to_unsigned(876, 10), 1952 => to_unsigned(518, 10), 1953 => to_unsigned(517, 10), 1954 => to_unsigned(538, 10), 1955 => to_unsigned(938, 10), 1956 => to_unsigned(1005, 10), 1957 => to_unsigned(570, 10), 1958 => to_unsigned(497, 10), 1959 => to_unsigned(754, 10), 1960 => to_unsigned(656, 10), 1961 => to_unsigned(343, 10), 1962 => to_unsigned(539, 10), 1963 => to_unsigned(121, 10), 1964 => to_unsigned(537, 10), 1965 => to_unsigned(677, 10), 1966 => to_unsigned(217, 10), 1967 => to_unsigned(314, 10), 1968 => to_unsigned(626, 10), 1969 => to_unsigned(758, 10), 1970 => to_unsigned(871, 10), 1971 => to_unsigned(192, 10), 1972 => to_unsigned(338, 10), 1973 => to_unsigned(985, 10), 1974 => to_unsigned(226, 10), 1975 => to_unsigned(847, 10), 1976 => to_unsigned(780, 10), 1977 => to_unsigned(521, 10), 1978 => to_unsigned(839, 10), 1979 => to_unsigned(474, 10), 1980 => to_unsigned(409, 10), 1981 => to_unsigned(258, 10), 1982 => to_unsigned(876, 10), 1983 => to_unsigned(1011, 10), 1984 => to_unsigned(1021, 10), 1985 => to_unsigned(184, 10), 1986 => to_unsigned(867, 10), 1987 => to_unsigned(552, 10), 1988 => to_unsigned(967, 10), 1989 => to_unsigned(543, 10), 1990 => to_unsigned(466, 10), 1991 => to_unsigned(971, 10), 1992 => to_unsigned(1019, 10), 1993 => to_unsigned(895, 10), 1994 => to_unsigned(940, 10), 1995 => to_unsigned(383, 10), 1996 => to_unsigned(172, 10), 1997 => to_unsigned(76, 10), 1998 => to_unsigned(555, 10), 1999 => to_unsigned(367, 10), 2000 => to_unsigned(236, 10), 2001 => to_unsigned(506, 10), 2002 => to_unsigned(434, 10), 2003 => to_unsigned(454, 10), 2004 => to_unsigned(46, 10), 2005 => to_unsigned(878, 10), 2006 => to_unsigned(975, 10), 2007 => to_unsigned(607, 10), 2008 => to_unsigned(456, 10), 2009 => to_unsigned(25, 10), 2010 => to_unsigned(367, 10), 2011 => to_unsigned(884, 10), 2012 => to_unsigned(124, 10), 2013 => to_unsigned(807, 10), 2014 => to_unsigned(174, 10), 2015 => to_unsigned(787, 10), 2016 => to_unsigned(965, 10), 2017 => to_unsigned(714, 10), 2018 => to_unsigned(220, 10), 2019 => to_unsigned(70, 10), 2020 => to_unsigned(732, 10), 2021 => to_unsigned(633, 10), 2022 => to_unsigned(42, 10), 2023 => to_unsigned(835, 10), 2024 => to_unsigned(314, 10), 2025 => to_unsigned(599, 10), 2026 => to_unsigned(706, 10), 2027 => to_unsigned(459, 10), 2028 => to_unsigned(674, 10), 2029 => to_unsigned(181, 10), 2030 => to_unsigned(199, 10), 2031 => to_unsigned(421, 10), 2032 => to_unsigned(828, 10), 2033 => to_unsigned(488, 10), 2034 => to_unsigned(997, 10), 2035 => to_unsigned(952, 10), 2036 => to_unsigned(462, 10), 2037 => to_unsigned(196, 10), 2038 => to_unsigned(568, 10), 2039 => to_unsigned(935, 10), 2040 => to_unsigned(760, 10), 2041 => to_unsigned(124, 10), 2042 => to_unsigned(463, 10), 2043 => to_unsigned(958, 10), 2044 => to_unsigned(301, 10), 2045 => to_unsigned(539, 10), 2046 => to_unsigned(268, 10), 2047 => to_unsigned(360, 10)),
            4 => (0 => to_unsigned(202, 10), 1 => to_unsigned(164, 10), 2 => to_unsigned(635, 10), 3 => to_unsigned(834, 10), 4 => to_unsigned(135, 10), 5 => to_unsigned(741, 10), 6 => to_unsigned(302, 10), 7 => to_unsigned(417, 10), 8 => to_unsigned(293, 10), 9 => to_unsigned(745, 10), 10 => to_unsigned(535, 10), 11 => to_unsigned(849, 10), 12 => to_unsigned(664, 10), 13 => to_unsigned(697, 10), 14 => to_unsigned(185, 10), 15 => to_unsigned(308, 10), 16 => to_unsigned(305, 10), 17 => to_unsigned(332, 10), 18 => to_unsigned(614, 10), 19 => to_unsigned(981, 10), 20 => to_unsigned(349, 10), 21 => to_unsigned(157, 10), 22 => to_unsigned(569, 10), 23 => to_unsigned(740, 10), 24 => to_unsigned(44, 10), 25 => to_unsigned(170, 10), 26 => to_unsigned(846, 10), 27 => to_unsigned(226, 10), 28 => to_unsigned(382, 10), 29 => to_unsigned(837, 10), 30 => to_unsigned(266, 10), 31 => to_unsigned(795, 10), 32 => to_unsigned(477, 10), 33 => to_unsigned(143, 10), 34 => to_unsigned(731, 10), 35 => to_unsigned(24, 10), 36 => to_unsigned(175, 10), 37 => to_unsigned(349, 10), 38 => to_unsigned(693, 10), 39 => to_unsigned(1004, 10), 40 => to_unsigned(909, 10), 41 => to_unsigned(858, 10), 42 => to_unsigned(687, 10), 43 => to_unsigned(945, 10), 44 => to_unsigned(29, 10), 45 => to_unsigned(892, 10), 46 => to_unsigned(905, 10), 47 => to_unsigned(505, 10), 48 => to_unsigned(83, 10), 49 => to_unsigned(427, 10), 50 => to_unsigned(710, 10), 51 => to_unsigned(434, 10), 52 => to_unsigned(545, 10), 53 => to_unsigned(51, 10), 54 => to_unsigned(154, 10), 55 => to_unsigned(342, 10), 56 => to_unsigned(949, 10), 57 => to_unsigned(45, 10), 58 => to_unsigned(108, 10), 59 => to_unsigned(728, 10), 60 => to_unsigned(91, 10), 61 => to_unsigned(977, 10), 62 => to_unsigned(908, 10), 63 => to_unsigned(652, 10), 64 => to_unsigned(748, 10), 65 => to_unsigned(673, 10), 66 => to_unsigned(205, 10), 67 => to_unsigned(923, 10), 68 => to_unsigned(268, 10), 69 => to_unsigned(865, 10), 70 => to_unsigned(580, 10), 71 => to_unsigned(743, 10), 72 => to_unsigned(969, 10), 73 => to_unsigned(355, 10), 74 => to_unsigned(133, 10), 75 => to_unsigned(1010, 10), 76 => to_unsigned(84, 10), 77 => to_unsigned(866, 10), 78 => to_unsigned(783, 10), 79 => to_unsigned(127, 10), 80 => to_unsigned(531, 10), 81 => to_unsigned(829, 10), 82 => to_unsigned(670, 10), 83 => to_unsigned(964, 10), 84 => to_unsigned(133, 10), 85 => to_unsigned(705, 10), 86 => to_unsigned(806, 10), 87 => to_unsigned(213, 10), 88 => to_unsigned(330, 10), 89 => to_unsigned(78, 10), 90 => to_unsigned(51, 10), 91 => to_unsigned(716, 10), 92 => to_unsigned(288, 10), 93 => to_unsigned(252, 10), 94 => to_unsigned(301, 10), 95 => to_unsigned(13, 10), 96 => to_unsigned(486, 10), 97 => to_unsigned(833, 10), 98 => to_unsigned(502, 10), 99 => to_unsigned(265, 10), 100 => to_unsigned(178, 10), 101 => to_unsigned(233, 10), 102 => to_unsigned(157, 10), 103 => to_unsigned(735, 10), 104 => to_unsigned(968, 10), 105 => to_unsigned(47, 10), 106 => to_unsigned(15, 10), 107 => to_unsigned(38, 10), 108 => to_unsigned(132, 10), 109 => to_unsigned(813, 10), 110 => to_unsigned(206, 10), 111 => to_unsigned(771, 10), 112 => to_unsigned(215, 10), 113 => to_unsigned(956, 10), 114 => to_unsigned(856, 10), 115 => to_unsigned(740, 10), 116 => to_unsigned(407, 10), 117 => to_unsigned(681, 10), 118 => to_unsigned(780, 10), 119 => to_unsigned(531, 10), 120 => to_unsigned(260, 10), 121 => to_unsigned(434, 10), 122 => to_unsigned(244, 10), 123 => to_unsigned(467, 10), 124 => to_unsigned(913, 10), 125 => to_unsigned(230, 10), 126 => to_unsigned(304, 10), 127 => to_unsigned(194, 10), 128 => to_unsigned(242, 10), 129 => to_unsigned(939, 10), 130 => to_unsigned(606, 10), 131 => to_unsigned(989, 10), 132 => to_unsigned(104, 10), 133 => to_unsigned(535, 10), 134 => to_unsigned(184, 10), 135 => to_unsigned(318, 10), 136 => to_unsigned(886, 10), 137 => to_unsigned(324, 10), 138 => to_unsigned(211, 10), 139 => to_unsigned(759, 10), 140 => to_unsigned(23, 10), 141 => to_unsigned(400, 10), 142 => to_unsigned(71, 10), 143 => to_unsigned(532, 10), 144 => to_unsigned(973, 10), 145 => to_unsigned(758, 10), 146 => to_unsigned(241, 10), 147 => to_unsigned(485, 10), 148 => to_unsigned(799, 10), 149 => to_unsigned(675, 10), 150 => to_unsigned(59, 10), 151 => to_unsigned(103, 10), 152 => to_unsigned(835, 10), 153 => to_unsigned(376, 10), 154 => to_unsigned(212, 10), 155 => to_unsigned(792, 10), 156 => to_unsigned(364, 10), 157 => to_unsigned(960, 10), 158 => to_unsigned(814, 10), 159 => to_unsigned(652, 10), 160 => to_unsigned(655, 10), 161 => to_unsigned(476, 10), 162 => to_unsigned(422, 10), 163 => to_unsigned(253, 10), 164 => to_unsigned(604, 10), 165 => to_unsigned(523, 10), 166 => to_unsigned(542, 10), 167 => to_unsigned(339, 10), 168 => to_unsigned(572, 10), 169 => to_unsigned(738, 10), 170 => to_unsigned(488, 10), 171 => to_unsigned(475, 10), 172 => to_unsigned(610, 10), 173 => to_unsigned(184, 10), 174 => to_unsigned(860, 10), 175 => to_unsigned(875, 10), 176 => to_unsigned(678, 10), 177 => to_unsigned(604, 10), 178 => to_unsigned(481, 10), 179 => to_unsigned(841, 10), 180 => to_unsigned(100, 10), 181 => to_unsigned(815, 10), 182 => to_unsigned(947, 10), 183 => to_unsigned(774, 10), 184 => to_unsigned(392, 10), 185 => to_unsigned(271, 10), 186 => to_unsigned(247, 10), 187 => to_unsigned(916, 10), 188 => to_unsigned(845, 10), 189 => to_unsigned(897, 10), 190 => to_unsigned(630, 10), 191 => to_unsigned(561, 10), 192 => to_unsigned(601, 10), 193 => to_unsigned(609, 10), 194 => to_unsigned(174, 10), 195 => to_unsigned(304, 10), 196 => to_unsigned(209, 10), 197 => to_unsigned(971, 10), 198 => to_unsigned(305, 10), 199 => to_unsigned(466, 10), 200 => to_unsigned(227, 10), 201 => to_unsigned(741, 10), 202 => to_unsigned(527, 10), 203 => to_unsigned(173, 10), 204 => to_unsigned(391, 10), 205 => to_unsigned(72, 10), 206 => to_unsigned(195, 10), 207 => to_unsigned(163, 10), 208 => to_unsigned(374, 10), 209 => to_unsigned(366, 10), 210 => to_unsigned(613, 10), 211 => to_unsigned(829, 10), 212 => to_unsigned(560, 10), 213 => to_unsigned(624, 10), 214 => to_unsigned(684, 10), 215 => to_unsigned(755, 10), 216 => to_unsigned(707, 10), 217 => to_unsigned(711, 10), 218 => to_unsigned(106, 10), 219 => to_unsigned(6, 10), 220 => to_unsigned(130, 10), 221 => to_unsigned(567, 10), 222 => to_unsigned(0, 10), 223 => to_unsigned(771, 10), 224 => to_unsigned(703, 10), 225 => to_unsigned(448, 10), 226 => to_unsigned(365, 10), 227 => to_unsigned(489, 10), 228 => to_unsigned(187, 10), 229 => to_unsigned(569, 10), 230 => to_unsigned(421, 10), 231 => to_unsigned(356, 10), 232 => to_unsigned(523, 10), 233 => to_unsigned(361, 10), 234 => to_unsigned(393, 10), 235 => to_unsigned(942, 10), 236 => to_unsigned(629, 10), 237 => to_unsigned(0, 10), 238 => to_unsigned(1, 10), 239 => to_unsigned(395, 10), 240 => to_unsigned(870, 10), 241 => to_unsigned(495, 10), 242 => to_unsigned(547, 10), 243 => to_unsigned(518, 10), 244 => to_unsigned(187, 10), 245 => to_unsigned(504, 10), 246 => to_unsigned(741, 10), 247 => to_unsigned(216, 10), 248 => to_unsigned(66, 10), 249 => to_unsigned(57, 10), 250 => to_unsigned(282, 10), 251 => to_unsigned(113, 10), 252 => to_unsigned(215, 10), 253 => to_unsigned(346, 10), 254 => to_unsigned(389, 10), 255 => to_unsigned(408, 10), 256 => to_unsigned(375, 10), 257 => to_unsigned(106, 10), 258 => to_unsigned(990, 10), 259 => to_unsigned(427, 10), 260 => to_unsigned(392, 10), 261 => to_unsigned(632, 10), 262 => to_unsigned(230, 10), 263 => to_unsigned(759, 10), 264 => to_unsigned(189, 10), 265 => to_unsigned(412, 10), 266 => to_unsigned(77, 10), 267 => to_unsigned(867, 10), 268 => to_unsigned(113, 10), 269 => to_unsigned(220, 10), 270 => to_unsigned(106, 10), 271 => to_unsigned(552, 10), 272 => to_unsigned(677, 10), 273 => to_unsigned(597, 10), 274 => to_unsigned(523, 10), 275 => to_unsigned(295, 10), 276 => to_unsigned(944, 10), 277 => to_unsigned(89, 10), 278 => to_unsigned(237, 10), 279 => to_unsigned(411, 10), 280 => to_unsigned(852, 10), 281 => to_unsigned(474, 10), 282 => to_unsigned(224, 10), 283 => to_unsigned(954, 10), 284 => to_unsigned(732, 10), 285 => to_unsigned(1014, 10), 286 => to_unsigned(575, 10), 287 => to_unsigned(535, 10), 288 => to_unsigned(31, 10), 289 => to_unsigned(325, 10), 290 => to_unsigned(955, 10), 291 => to_unsigned(538, 10), 292 => to_unsigned(975, 10), 293 => to_unsigned(99, 10), 294 => to_unsigned(174, 10), 295 => to_unsigned(605, 10), 296 => to_unsigned(206, 10), 297 => to_unsigned(187, 10), 298 => to_unsigned(391, 10), 299 => to_unsigned(566, 10), 300 => to_unsigned(414, 10), 301 => to_unsigned(520, 10), 302 => to_unsigned(489, 10), 303 => to_unsigned(183, 10), 304 => to_unsigned(532, 10), 305 => to_unsigned(678, 10), 306 => to_unsigned(870, 10), 307 => to_unsigned(952, 10), 308 => to_unsigned(42, 10), 309 => to_unsigned(467, 10), 310 => to_unsigned(601, 10), 311 => to_unsigned(741, 10), 312 => to_unsigned(234, 10), 313 => to_unsigned(1016, 10), 314 => to_unsigned(717, 10), 315 => to_unsigned(435, 10), 316 => to_unsigned(691, 10), 317 => to_unsigned(815, 10), 318 => to_unsigned(680, 10), 319 => to_unsigned(566, 10), 320 => to_unsigned(532, 10), 321 => to_unsigned(948, 10), 322 => to_unsigned(884, 10), 323 => to_unsigned(274, 10), 324 => to_unsigned(893, 10), 325 => to_unsigned(61, 10), 326 => to_unsigned(909, 10), 327 => to_unsigned(887, 10), 328 => to_unsigned(264, 10), 329 => to_unsigned(297, 10), 330 => to_unsigned(249, 10), 331 => to_unsigned(67, 10), 332 => to_unsigned(319, 10), 333 => to_unsigned(918, 10), 334 => to_unsigned(85, 10), 335 => to_unsigned(723, 10), 336 => to_unsigned(274, 10), 337 => to_unsigned(82, 10), 338 => to_unsigned(726, 10), 339 => to_unsigned(286, 10), 340 => to_unsigned(179, 10), 341 => to_unsigned(893, 10), 342 => to_unsigned(507, 10), 343 => to_unsigned(749, 10), 344 => to_unsigned(124, 10), 345 => to_unsigned(594, 10), 346 => to_unsigned(939, 10), 347 => to_unsigned(595, 10), 348 => to_unsigned(374, 10), 349 => to_unsigned(153, 10), 350 => to_unsigned(837, 10), 351 => to_unsigned(411, 10), 352 => to_unsigned(296, 10), 353 => to_unsigned(190, 10), 354 => to_unsigned(117, 10), 355 => to_unsigned(451, 10), 356 => to_unsigned(880, 10), 357 => to_unsigned(107, 10), 358 => to_unsigned(72, 10), 359 => to_unsigned(816, 10), 360 => to_unsigned(525, 10), 361 => to_unsigned(286, 10), 362 => to_unsigned(318, 10), 363 => to_unsigned(372, 10), 364 => to_unsigned(668, 10), 365 => to_unsigned(624, 10), 366 => to_unsigned(21, 10), 367 => to_unsigned(892, 10), 368 => to_unsigned(1015, 10), 369 => to_unsigned(572, 10), 370 => to_unsigned(72, 10), 371 => to_unsigned(63, 10), 372 => to_unsigned(906, 10), 373 => to_unsigned(638, 10), 374 => to_unsigned(152, 10), 375 => to_unsigned(161, 10), 376 => to_unsigned(613, 10), 377 => to_unsigned(324, 10), 378 => to_unsigned(686, 10), 379 => to_unsigned(214, 10), 380 => to_unsigned(533, 10), 381 => to_unsigned(164, 10), 382 => to_unsigned(42, 10), 383 => to_unsigned(878, 10), 384 => to_unsigned(70, 10), 385 => to_unsigned(839, 10), 386 => to_unsigned(566, 10), 387 => to_unsigned(714, 10), 388 => to_unsigned(552, 10), 389 => to_unsigned(865, 10), 390 => to_unsigned(283, 10), 391 => to_unsigned(778, 10), 392 => to_unsigned(377, 10), 393 => to_unsigned(241, 10), 394 => to_unsigned(1022, 10), 395 => to_unsigned(160, 10), 396 => to_unsigned(85, 10), 397 => to_unsigned(601, 10), 398 => to_unsigned(645, 10), 399 => to_unsigned(581, 10), 400 => to_unsigned(466, 10), 401 => to_unsigned(845, 10), 402 => to_unsigned(226, 10), 403 => to_unsigned(495, 10), 404 => to_unsigned(46, 10), 405 => to_unsigned(228, 10), 406 => to_unsigned(640, 10), 407 => to_unsigned(407, 10), 408 => to_unsigned(199, 10), 409 => to_unsigned(440, 10), 410 => to_unsigned(704, 10), 411 => to_unsigned(252, 10), 412 => to_unsigned(912, 10), 413 => to_unsigned(429, 10), 414 => to_unsigned(739, 10), 415 => to_unsigned(874, 10), 416 => to_unsigned(1010, 10), 417 => to_unsigned(65, 10), 418 => to_unsigned(528, 10), 419 => to_unsigned(776, 10), 420 => to_unsigned(1001, 10), 421 => to_unsigned(124, 10), 422 => to_unsigned(281, 10), 423 => to_unsigned(745, 10), 424 => to_unsigned(389, 10), 425 => to_unsigned(389, 10), 426 => to_unsigned(626, 10), 427 => to_unsigned(80, 10), 428 => to_unsigned(547, 10), 429 => to_unsigned(955, 10), 430 => to_unsigned(716, 10), 431 => to_unsigned(548, 10), 432 => to_unsigned(616, 10), 433 => to_unsigned(743, 10), 434 => to_unsigned(189, 10), 435 => to_unsigned(969, 10), 436 => to_unsigned(506, 10), 437 => to_unsigned(66, 10), 438 => to_unsigned(413, 10), 439 => to_unsigned(909, 10), 440 => to_unsigned(280, 10), 441 => to_unsigned(1020, 10), 442 => to_unsigned(1011, 10), 443 => to_unsigned(196, 10), 444 => to_unsigned(317, 10), 445 => to_unsigned(511, 10), 446 => to_unsigned(338, 10), 447 => to_unsigned(7, 10), 448 => to_unsigned(820, 10), 449 => to_unsigned(61, 10), 450 => to_unsigned(983, 10), 451 => to_unsigned(37, 10), 452 => to_unsigned(147, 10), 453 => to_unsigned(1001, 10), 454 => to_unsigned(512, 10), 455 => to_unsigned(646, 10), 456 => to_unsigned(412, 10), 457 => to_unsigned(823, 10), 458 => to_unsigned(252, 10), 459 => to_unsigned(297, 10), 460 => to_unsigned(232, 10), 461 => to_unsigned(383, 10), 462 => to_unsigned(349, 10), 463 => to_unsigned(927, 10), 464 => to_unsigned(431, 10), 465 => to_unsigned(77, 10), 466 => to_unsigned(254, 10), 467 => to_unsigned(728, 10), 468 => to_unsigned(1016, 10), 469 => to_unsigned(209, 10), 470 => to_unsigned(905, 10), 471 => to_unsigned(917, 10), 472 => to_unsigned(972, 10), 473 => to_unsigned(607, 10), 474 => to_unsigned(628, 10), 475 => to_unsigned(834, 10), 476 => to_unsigned(811, 10), 477 => to_unsigned(657, 10), 478 => to_unsigned(480, 10), 479 => to_unsigned(213, 10), 480 => to_unsigned(604, 10), 481 => to_unsigned(627, 10), 482 => to_unsigned(746, 10), 483 => to_unsigned(184, 10), 484 => to_unsigned(3, 10), 485 => to_unsigned(604, 10), 486 => to_unsigned(657, 10), 487 => to_unsigned(128, 10), 488 => to_unsigned(519, 10), 489 => to_unsigned(542, 10), 490 => to_unsigned(494, 10), 491 => to_unsigned(617, 10), 492 => to_unsigned(724, 10), 493 => to_unsigned(101, 10), 494 => to_unsigned(712, 10), 495 => to_unsigned(624, 10), 496 => to_unsigned(300, 10), 497 => to_unsigned(851, 10), 498 => to_unsigned(470, 10), 499 => to_unsigned(391, 10), 500 => to_unsigned(73, 10), 501 => to_unsigned(556, 10), 502 => to_unsigned(531, 10), 503 => to_unsigned(963, 10), 504 => to_unsigned(918, 10), 505 => to_unsigned(736, 10), 506 => to_unsigned(177, 10), 507 => to_unsigned(257, 10), 508 => to_unsigned(933, 10), 509 => to_unsigned(529, 10), 510 => to_unsigned(183, 10), 511 => to_unsigned(844, 10), 512 => to_unsigned(817, 10), 513 => to_unsigned(650, 10), 514 => to_unsigned(568, 10), 515 => to_unsigned(787, 10), 516 => to_unsigned(129, 10), 517 => to_unsigned(179, 10), 518 => to_unsigned(940, 10), 519 => to_unsigned(780, 10), 520 => to_unsigned(975, 10), 521 => to_unsigned(498, 10), 522 => to_unsigned(22, 10), 523 => to_unsigned(58, 10), 524 => to_unsigned(237, 10), 525 => to_unsigned(434, 10), 526 => to_unsigned(475, 10), 527 => to_unsigned(180, 10), 528 => to_unsigned(140, 10), 529 => to_unsigned(25, 10), 530 => to_unsigned(613, 10), 531 => to_unsigned(771, 10), 532 => to_unsigned(512, 10), 533 => to_unsigned(509, 10), 534 => to_unsigned(468, 10), 535 => to_unsigned(280, 10), 536 => to_unsigned(376, 10), 537 => to_unsigned(754, 10), 538 => to_unsigned(439, 10), 539 => to_unsigned(653, 10), 540 => to_unsigned(818, 10), 541 => to_unsigned(819, 10), 542 => to_unsigned(922, 10), 543 => to_unsigned(230, 10), 544 => to_unsigned(894, 10), 545 => to_unsigned(64, 10), 546 => to_unsigned(118, 10), 547 => to_unsigned(346, 10), 548 => to_unsigned(96, 10), 549 => to_unsigned(896, 10), 550 => to_unsigned(516, 10), 551 => to_unsigned(676, 10), 552 => to_unsigned(829, 10), 553 => to_unsigned(609, 10), 554 => to_unsigned(102, 10), 555 => to_unsigned(132, 10), 556 => to_unsigned(435, 10), 557 => to_unsigned(785, 10), 558 => to_unsigned(480, 10), 559 => to_unsigned(202, 10), 560 => to_unsigned(547, 10), 561 => to_unsigned(51, 10), 562 => to_unsigned(1023, 10), 563 => to_unsigned(957, 10), 564 => to_unsigned(59, 10), 565 => to_unsigned(165, 10), 566 => to_unsigned(52, 10), 567 => to_unsigned(164, 10), 568 => to_unsigned(214, 10), 569 => to_unsigned(789, 10), 570 => to_unsigned(216, 10), 571 => to_unsigned(940, 10), 572 => to_unsigned(48, 10), 573 => to_unsigned(765, 10), 574 => to_unsigned(844, 10), 575 => to_unsigned(482, 10), 576 => to_unsigned(179, 10), 577 => to_unsigned(508, 10), 578 => to_unsigned(444, 10), 579 => to_unsigned(173, 10), 580 => to_unsigned(235, 10), 581 => to_unsigned(179, 10), 582 => to_unsigned(102, 10), 583 => to_unsigned(449, 10), 584 => to_unsigned(820, 10), 585 => to_unsigned(464, 10), 586 => to_unsigned(800, 10), 587 => to_unsigned(82, 10), 588 => to_unsigned(31, 10), 589 => to_unsigned(616, 10), 590 => to_unsigned(181, 10), 591 => to_unsigned(346, 10), 592 => to_unsigned(183, 10), 593 => to_unsigned(910, 10), 594 => to_unsigned(887, 10), 595 => to_unsigned(348, 10), 596 => to_unsigned(50, 10), 597 => to_unsigned(928, 10), 598 => to_unsigned(451, 10), 599 => to_unsigned(491, 10), 600 => to_unsigned(562, 10), 601 => to_unsigned(516, 10), 602 => to_unsigned(375, 10), 603 => to_unsigned(192, 10), 604 => to_unsigned(54, 10), 605 => to_unsigned(210, 10), 606 => to_unsigned(710, 10), 607 => to_unsigned(635, 10), 608 => to_unsigned(762, 10), 609 => to_unsigned(738, 10), 610 => to_unsigned(75, 10), 611 => to_unsigned(219, 10), 612 => to_unsigned(911, 10), 613 => to_unsigned(513, 10), 614 => to_unsigned(868, 10), 615 => to_unsigned(631, 10), 616 => to_unsigned(993, 10), 617 => to_unsigned(169, 10), 618 => to_unsigned(785, 10), 619 => to_unsigned(757, 10), 620 => to_unsigned(196, 10), 621 => to_unsigned(456, 10), 622 => to_unsigned(659, 10), 623 => to_unsigned(835, 10), 624 => to_unsigned(464, 10), 625 => to_unsigned(931, 10), 626 => to_unsigned(392, 10), 627 => to_unsigned(906, 10), 628 => to_unsigned(546, 10), 629 => to_unsigned(930, 10), 630 => to_unsigned(690, 10), 631 => to_unsigned(222, 10), 632 => to_unsigned(478, 10), 633 => to_unsigned(278, 10), 634 => to_unsigned(65, 10), 635 => to_unsigned(137, 10), 636 => to_unsigned(554, 10), 637 => to_unsigned(273, 10), 638 => to_unsigned(705, 10), 639 => to_unsigned(888, 10), 640 => to_unsigned(854, 10), 641 => to_unsigned(749, 10), 642 => to_unsigned(392, 10), 643 => to_unsigned(20, 10), 644 => to_unsigned(190, 10), 645 => to_unsigned(397, 10), 646 => to_unsigned(160, 10), 647 => to_unsigned(99, 10), 648 => to_unsigned(681, 10), 649 => to_unsigned(205, 10), 650 => to_unsigned(754, 10), 651 => to_unsigned(679, 10), 652 => to_unsigned(175, 10), 653 => to_unsigned(459, 10), 654 => to_unsigned(918, 10), 655 => to_unsigned(45, 10), 656 => to_unsigned(495, 10), 657 => to_unsigned(937, 10), 658 => to_unsigned(56, 10), 659 => to_unsigned(441, 10), 660 => to_unsigned(48, 10), 661 => to_unsigned(737, 10), 662 => to_unsigned(975, 10), 663 => to_unsigned(525, 10), 664 => to_unsigned(528, 10), 665 => to_unsigned(739, 10), 666 => to_unsigned(367, 10), 667 => to_unsigned(315, 10), 668 => to_unsigned(886, 10), 669 => to_unsigned(889, 10), 670 => to_unsigned(11, 10), 671 => to_unsigned(606, 10), 672 => to_unsigned(917, 10), 673 => to_unsigned(996, 10), 674 => to_unsigned(743, 10), 675 => to_unsigned(845, 10), 676 => to_unsigned(134, 10), 677 => to_unsigned(923, 10), 678 => to_unsigned(530, 10), 679 => to_unsigned(813, 10), 680 => to_unsigned(977, 10), 681 => to_unsigned(957, 10), 682 => to_unsigned(159, 10), 683 => to_unsigned(858, 10), 684 => to_unsigned(21, 10), 685 => to_unsigned(607, 10), 686 => to_unsigned(584, 10), 687 => to_unsigned(939, 10), 688 => to_unsigned(389, 10), 689 => to_unsigned(69, 10), 690 => to_unsigned(272, 10), 691 => to_unsigned(768, 10), 692 => to_unsigned(983, 10), 693 => to_unsigned(961, 10), 694 => to_unsigned(312, 10), 695 => to_unsigned(677, 10), 696 => to_unsigned(310, 10), 697 => to_unsigned(967, 10), 698 => to_unsigned(957, 10), 699 => to_unsigned(587, 10), 700 => to_unsigned(483, 10), 701 => to_unsigned(621, 10), 702 => to_unsigned(932, 10), 703 => to_unsigned(989, 10), 704 => to_unsigned(851, 10), 705 => to_unsigned(553, 10), 706 => to_unsigned(698, 10), 707 => to_unsigned(587, 10), 708 => to_unsigned(903, 10), 709 => to_unsigned(142, 10), 710 => to_unsigned(155, 10), 711 => to_unsigned(50, 10), 712 => to_unsigned(613, 10), 713 => to_unsigned(325, 10), 714 => to_unsigned(776, 10), 715 => to_unsigned(436, 10), 716 => to_unsigned(324, 10), 717 => to_unsigned(46, 10), 718 => to_unsigned(208, 10), 719 => to_unsigned(205, 10), 720 => to_unsigned(726, 10), 721 => to_unsigned(697, 10), 722 => to_unsigned(938, 10), 723 => to_unsigned(210, 10), 724 => to_unsigned(785, 10), 725 => to_unsigned(893, 10), 726 => to_unsigned(745, 10), 727 => to_unsigned(899, 10), 728 => to_unsigned(213, 10), 729 => to_unsigned(760, 10), 730 => to_unsigned(79, 10), 731 => to_unsigned(556, 10), 732 => to_unsigned(188, 10), 733 => to_unsigned(973, 10), 734 => to_unsigned(19, 10), 735 => to_unsigned(857, 10), 736 => to_unsigned(388, 10), 737 => to_unsigned(7, 10), 738 => to_unsigned(359, 10), 739 => to_unsigned(981, 10), 740 => to_unsigned(146, 10), 741 => to_unsigned(373, 10), 742 => to_unsigned(319, 10), 743 => to_unsigned(355, 10), 744 => to_unsigned(607, 10), 745 => to_unsigned(244, 10), 746 => to_unsigned(409, 10), 747 => to_unsigned(32, 10), 748 => to_unsigned(209, 10), 749 => to_unsigned(461, 10), 750 => to_unsigned(765, 10), 751 => to_unsigned(119, 10), 752 => to_unsigned(119, 10), 753 => to_unsigned(499, 10), 754 => to_unsigned(27, 10), 755 => to_unsigned(1013, 10), 756 => to_unsigned(336, 10), 757 => to_unsigned(860, 10), 758 => to_unsigned(302, 10), 759 => to_unsigned(767, 10), 760 => to_unsigned(658, 10), 761 => to_unsigned(866, 10), 762 => to_unsigned(951, 10), 763 => to_unsigned(64, 10), 764 => to_unsigned(283, 10), 765 => to_unsigned(795, 10), 766 => to_unsigned(795, 10), 767 => to_unsigned(32, 10), 768 => to_unsigned(426, 10), 769 => to_unsigned(530, 10), 770 => to_unsigned(340, 10), 771 => to_unsigned(369, 10), 772 => to_unsigned(10, 10), 773 => to_unsigned(1019, 10), 774 => to_unsigned(691, 10), 775 => to_unsigned(584, 10), 776 => to_unsigned(44, 10), 777 => to_unsigned(79, 10), 778 => to_unsigned(290, 10), 779 => to_unsigned(235, 10), 780 => to_unsigned(120, 10), 781 => to_unsigned(962, 10), 782 => to_unsigned(161, 10), 783 => to_unsigned(198, 10), 784 => to_unsigned(159, 10), 785 => to_unsigned(549, 10), 786 => to_unsigned(257, 10), 787 => to_unsigned(908, 10), 788 => to_unsigned(732, 10), 789 => to_unsigned(248, 10), 790 => to_unsigned(1012, 10), 791 => to_unsigned(93, 10), 792 => to_unsigned(371, 10), 793 => to_unsigned(933, 10), 794 => to_unsigned(1020, 10), 795 => to_unsigned(622, 10), 796 => to_unsigned(565, 10), 797 => to_unsigned(272, 10), 798 => to_unsigned(312, 10), 799 => to_unsigned(1023, 10), 800 => to_unsigned(835, 10), 801 => to_unsigned(596, 10), 802 => to_unsigned(442, 10), 803 => to_unsigned(498, 10), 804 => to_unsigned(201, 10), 805 => to_unsigned(61, 10), 806 => to_unsigned(133, 10), 807 => to_unsigned(855, 10), 808 => to_unsigned(739, 10), 809 => to_unsigned(1021, 10), 810 => to_unsigned(975, 10), 811 => to_unsigned(227, 10), 812 => to_unsigned(638, 10), 813 => to_unsigned(127, 10), 814 => to_unsigned(728, 10), 815 => to_unsigned(657, 10), 816 => to_unsigned(14, 10), 817 => to_unsigned(347, 10), 818 => to_unsigned(250, 10), 819 => to_unsigned(216, 10), 820 => to_unsigned(237, 10), 821 => to_unsigned(972, 10), 822 => to_unsigned(246, 10), 823 => to_unsigned(658, 10), 824 => to_unsigned(287, 10), 825 => to_unsigned(766, 10), 826 => to_unsigned(113, 10), 827 => to_unsigned(684, 10), 828 => to_unsigned(883, 10), 829 => to_unsigned(56, 10), 830 => to_unsigned(631, 10), 831 => to_unsigned(22, 10), 832 => to_unsigned(864, 10), 833 => to_unsigned(959, 10), 834 => to_unsigned(14, 10), 835 => to_unsigned(124, 10), 836 => to_unsigned(113, 10), 837 => to_unsigned(369, 10), 838 => to_unsigned(1011, 10), 839 => to_unsigned(921, 10), 840 => to_unsigned(804, 10), 841 => to_unsigned(489, 10), 842 => to_unsigned(829, 10), 843 => to_unsigned(960, 10), 844 => to_unsigned(113, 10), 845 => to_unsigned(536, 10), 846 => to_unsigned(37, 10), 847 => to_unsigned(912, 10), 848 => to_unsigned(559, 10), 849 => to_unsigned(526, 10), 850 => to_unsigned(489, 10), 851 => to_unsigned(97, 10), 852 => to_unsigned(54, 10), 853 => to_unsigned(124, 10), 854 => to_unsigned(97, 10), 855 => to_unsigned(708, 10), 856 => to_unsigned(466, 10), 857 => to_unsigned(809, 10), 858 => to_unsigned(416, 10), 859 => to_unsigned(579, 10), 860 => to_unsigned(371, 10), 861 => to_unsigned(756, 10), 862 => to_unsigned(385, 10), 863 => to_unsigned(236, 10), 864 => to_unsigned(493, 10), 865 => to_unsigned(474, 10), 866 => to_unsigned(824, 10), 867 => to_unsigned(917, 10), 868 => to_unsigned(763, 10), 869 => to_unsigned(275, 10), 870 => to_unsigned(858, 10), 871 => to_unsigned(391, 10), 872 => to_unsigned(849, 10), 873 => to_unsigned(139, 10), 874 => to_unsigned(618, 10), 875 => to_unsigned(366, 10), 876 => to_unsigned(1, 10), 877 => to_unsigned(687, 10), 878 => to_unsigned(303, 10), 879 => to_unsigned(267, 10), 880 => to_unsigned(377, 10), 881 => to_unsigned(698, 10), 882 => to_unsigned(15, 10), 883 => to_unsigned(483, 10), 884 => to_unsigned(858, 10), 885 => to_unsigned(127, 10), 886 => to_unsigned(85, 10), 887 => to_unsigned(419, 10), 888 => to_unsigned(222, 10), 889 => to_unsigned(9, 10), 890 => to_unsigned(111, 10), 891 => to_unsigned(1012, 10), 892 => to_unsigned(322, 10), 893 => to_unsigned(760, 10), 894 => to_unsigned(381, 10), 895 => to_unsigned(490, 10), 896 => to_unsigned(832, 10), 897 => to_unsigned(894, 10), 898 => to_unsigned(375, 10), 899 => to_unsigned(522, 10), 900 => to_unsigned(269, 10), 901 => to_unsigned(269, 10), 902 => to_unsigned(660, 10), 903 => to_unsigned(168, 10), 904 => to_unsigned(672, 10), 905 => to_unsigned(79, 10), 906 => to_unsigned(750, 10), 907 => to_unsigned(417, 10), 908 => to_unsigned(25, 10), 909 => to_unsigned(501, 10), 910 => to_unsigned(749, 10), 911 => to_unsigned(255, 10), 912 => to_unsigned(889, 10), 913 => to_unsigned(710, 10), 914 => to_unsigned(289, 10), 915 => to_unsigned(486, 10), 916 => to_unsigned(952, 10), 917 => to_unsigned(667, 10), 918 => to_unsigned(497, 10), 919 => to_unsigned(847, 10), 920 => to_unsigned(944, 10), 921 => to_unsigned(363, 10), 922 => to_unsigned(557, 10), 923 => to_unsigned(66, 10), 924 => to_unsigned(667, 10), 925 => to_unsigned(184, 10), 926 => to_unsigned(487, 10), 927 => to_unsigned(609, 10), 928 => to_unsigned(456, 10), 929 => to_unsigned(521, 10), 930 => to_unsigned(547, 10), 931 => to_unsigned(219, 10), 932 => to_unsigned(690, 10), 933 => to_unsigned(658, 10), 934 => to_unsigned(706, 10), 935 => to_unsigned(905, 10), 936 => to_unsigned(971, 10), 937 => to_unsigned(353, 10), 938 => to_unsigned(937, 10), 939 => to_unsigned(162, 10), 940 => to_unsigned(205, 10), 941 => to_unsigned(37, 10), 942 => to_unsigned(590, 10), 943 => to_unsigned(67, 10), 944 => to_unsigned(648, 10), 945 => to_unsigned(324, 10), 946 => to_unsigned(288, 10), 947 => to_unsigned(507, 10), 948 => to_unsigned(422, 10), 949 => to_unsigned(739, 10), 950 => to_unsigned(138, 10), 951 => to_unsigned(915, 10), 952 => to_unsigned(990, 10), 953 => to_unsigned(927, 10), 954 => to_unsigned(837, 10), 955 => to_unsigned(144, 10), 956 => to_unsigned(383, 10), 957 => to_unsigned(844, 10), 958 => to_unsigned(741, 10), 959 => to_unsigned(599, 10), 960 => to_unsigned(502, 10), 961 => to_unsigned(612, 10), 962 => to_unsigned(940, 10), 963 => to_unsigned(916, 10), 964 => to_unsigned(175, 10), 965 => to_unsigned(841, 10), 966 => to_unsigned(926, 10), 967 => to_unsigned(555, 10), 968 => to_unsigned(46, 10), 969 => to_unsigned(838, 10), 970 => to_unsigned(115, 10), 971 => to_unsigned(583, 10), 972 => to_unsigned(955, 10), 973 => to_unsigned(113, 10), 974 => to_unsigned(993, 10), 975 => to_unsigned(495, 10), 976 => to_unsigned(60, 10), 977 => to_unsigned(692, 10), 978 => to_unsigned(170, 10), 979 => to_unsigned(244, 10), 980 => to_unsigned(545, 10), 981 => to_unsigned(68, 10), 982 => to_unsigned(186, 10), 983 => to_unsigned(451, 10), 984 => to_unsigned(404, 10), 985 => to_unsigned(511, 10), 986 => to_unsigned(124, 10), 987 => to_unsigned(487, 10), 988 => to_unsigned(1018, 10), 989 => to_unsigned(252, 10), 990 => to_unsigned(653, 10), 991 => to_unsigned(377, 10), 992 => to_unsigned(703, 10), 993 => to_unsigned(491, 10), 994 => to_unsigned(933, 10), 995 => to_unsigned(443, 10), 996 => to_unsigned(910, 10), 997 => to_unsigned(803, 10), 998 => to_unsigned(440, 10), 999 => to_unsigned(151, 10), 1000 => to_unsigned(698, 10), 1001 => to_unsigned(66, 10), 1002 => to_unsigned(484, 10), 1003 => to_unsigned(47, 10), 1004 => to_unsigned(933, 10), 1005 => to_unsigned(337, 10), 1006 => to_unsigned(465, 10), 1007 => to_unsigned(537, 10), 1008 => to_unsigned(722, 10), 1009 => to_unsigned(342, 10), 1010 => to_unsigned(841, 10), 1011 => to_unsigned(690, 10), 1012 => to_unsigned(893, 10), 1013 => to_unsigned(44, 10), 1014 => to_unsigned(186, 10), 1015 => to_unsigned(872, 10), 1016 => to_unsigned(16, 10), 1017 => to_unsigned(25, 10), 1018 => to_unsigned(261, 10), 1019 => to_unsigned(739, 10), 1020 => to_unsigned(124, 10), 1021 => to_unsigned(368, 10), 1022 => to_unsigned(839, 10), 1023 => to_unsigned(997, 10), 1024 => to_unsigned(604, 10), 1025 => to_unsigned(639, 10), 1026 => to_unsigned(706, 10), 1027 => to_unsigned(262, 10), 1028 => to_unsigned(1022, 10), 1029 => to_unsigned(150, 10), 1030 => to_unsigned(232, 10), 1031 => to_unsigned(1008, 10), 1032 => to_unsigned(0, 10), 1033 => to_unsigned(673, 10), 1034 => to_unsigned(200, 10), 1035 => to_unsigned(1008, 10), 1036 => to_unsigned(113, 10), 1037 => to_unsigned(329, 10), 1038 => to_unsigned(166, 10), 1039 => to_unsigned(33, 10), 1040 => to_unsigned(753, 10), 1041 => to_unsigned(927, 10), 1042 => to_unsigned(112, 10), 1043 => to_unsigned(333, 10), 1044 => to_unsigned(358, 10), 1045 => to_unsigned(80, 10), 1046 => to_unsigned(246, 10), 1047 => to_unsigned(500, 10), 1048 => to_unsigned(849, 10), 1049 => to_unsigned(193, 10), 1050 => to_unsigned(328, 10), 1051 => to_unsigned(979, 10), 1052 => to_unsigned(951, 10), 1053 => to_unsigned(115, 10), 1054 => to_unsigned(271, 10), 1055 => to_unsigned(1022, 10), 1056 => to_unsigned(96, 10), 1057 => to_unsigned(939, 10), 1058 => to_unsigned(396, 10), 1059 => to_unsigned(333, 10), 1060 => to_unsigned(877, 10), 1061 => to_unsigned(473, 10), 1062 => to_unsigned(426, 10), 1063 => to_unsigned(892, 10), 1064 => to_unsigned(243, 10), 1065 => to_unsigned(893, 10), 1066 => to_unsigned(644, 10), 1067 => to_unsigned(325, 10), 1068 => to_unsigned(480, 10), 1069 => to_unsigned(461, 10), 1070 => to_unsigned(192, 10), 1071 => to_unsigned(121, 10), 1072 => to_unsigned(928, 10), 1073 => to_unsigned(928, 10), 1074 => to_unsigned(791, 10), 1075 => to_unsigned(835, 10), 1076 => to_unsigned(780, 10), 1077 => to_unsigned(394, 10), 1078 => to_unsigned(94, 10), 1079 => to_unsigned(568, 10), 1080 => to_unsigned(405, 10), 1081 => to_unsigned(938, 10), 1082 => to_unsigned(501, 10), 1083 => to_unsigned(125, 10), 1084 => to_unsigned(707, 10), 1085 => to_unsigned(539, 10), 1086 => to_unsigned(161, 10), 1087 => to_unsigned(731, 10), 1088 => to_unsigned(421, 10), 1089 => to_unsigned(363, 10), 1090 => to_unsigned(515, 10), 1091 => to_unsigned(868, 10), 1092 => to_unsigned(793, 10), 1093 => to_unsigned(610, 10), 1094 => to_unsigned(312, 10), 1095 => to_unsigned(960, 10), 1096 => to_unsigned(844, 10), 1097 => to_unsigned(12, 10), 1098 => to_unsigned(107, 10), 1099 => to_unsigned(525, 10), 1100 => to_unsigned(259, 10), 1101 => to_unsigned(205, 10), 1102 => to_unsigned(968, 10), 1103 => to_unsigned(785, 10), 1104 => to_unsigned(927, 10), 1105 => to_unsigned(32, 10), 1106 => to_unsigned(744, 10), 1107 => to_unsigned(593, 10), 1108 => to_unsigned(114, 10), 1109 => to_unsigned(262, 10), 1110 => to_unsigned(1009, 10), 1111 => to_unsigned(322, 10), 1112 => to_unsigned(802, 10), 1113 => to_unsigned(588, 10), 1114 => to_unsigned(465, 10), 1115 => to_unsigned(535, 10), 1116 => to_unsigned(680, 10), 1117 => to_unsigned(882, 10), 1118 => to_unsigned(591, 10), 1119 => to_unsigned(162, 10), 1120 => to_unsigned(803, 10), 1121 => to_unsigned(988, 10), 1122 => to_unsigned(670, 10), 1123 => to_unsigned(37, 10), 1124 => to_unsigned(297, 10), 1125 => to_unsigned(231, 10), 1126 => to_unsigned(637, 10), 1127 => to_unsigned(690, 10), 1128 => to_unsigned(856, 10), 1129 => to_unsigned(453, 10), 1130 => to_unsigned(161, 10), 1131 => to_unsigned(472, 10), 1132 => to_unsigned(215, 10), 1133 => to_unsigned(617, 10), 1134 => to_unsigned(862, 10), 1135 => to_unsigned(873, 10), 1136 => to_unsigned(689, 10), 1137 => to_unsigned(987, 10), 1138 => to_unsigned(155, 10), 1139 => to_unsigned(509, 10), 1140 => to_unsigned(609, 10), 1141 => to_unsigned(860, 10), 1142 => to_unsigned(938, 10), 1143 => to_unsigned(743, 10), 1144 => to_unsigned(822, 10), 1145 => to_unsigned(722, 10), 1146 => to_unsigned(627, 10), 1147 => to_unsigned(152, 10), 1148 => to_unsigned(620, 10), 1149 => to_unsigned(971, 10), 1150 => to_unsigned(590, 10), 1151 => to_unsigned(58, 10), 1152 => to_unsigned(1012, 10), 1153 => to_unsigned(325, 10), 1154 => to_unsigned(114, 10), 1155 => to_unsigned(371, 10), 1156 => to_unsigned(612, 10), 1157 => to_unsigned(321, 10), 1158 => to_unsigned(145, 10), 1159 => to_unsigned(829, 10), 1160 => to_unsigned(81, 10), 1161 => to_unsigned(233, 10), 1162 => to_unsigned(570, 10), 1163 => to_unsigned(132, 10), 1164 => to_unsigned(992, 10), 1165 => to_unsigned(951, 10), 1166 => to_unsigned(955, 10), 1167 => to_unsigned(364, 10), 1168 => to_unsigned(593, 10), 1169 => to_unsigned(547, 10), 1170 => to_unsigned(68, 10), 1171 => to_unsigned(161, 10), 1172 => to_unsigned(7, 10), 1173 => to_unsigned(524, 10), 1174 => to_unsigned(749, 10), 1175 => to_unsigned(784, 10), 1176 => to_unsigned(363, 10), 1177 => to_unsigned(754, 10), 1178 => to_unsigned(613, 10), 1179 => to_unsigned(210, 10), 1180 => to_unsigned(409, 10), 1181 => to_unsigned(343, 10), 1182 => to_unsigned(487, 10), 1183 => to_unsigned(19, 10), 1184 => to_unsigned(86, 10), 1185 => to_unsigned(48, 10), 1186 => to_unsigned(111, 10), 1187 => to_unsigned(988, 10), 1188 => to_unsigned(494, 10), 1189 => to_unsigned(336, 10), 1190 => to_unsigned(502, 10), 1191 => to_unsigned(540, 10), 1192 => to_unsigned(91, 10), 1193 => to_unsigned(96, 10), 1194 => to_unsigned(894, 10), 1195 => to_unsigned(100, 10), 1196 => to_unsigned(39, 10), 1197 => to_unsigned(979, 10), 1198 => to_unsigned(193, 10), 1199 => to_unsigned(377, 10), 1200 => to_unsigned(477, 10), 1201 => to_unsigned(551, 10), 1202 => to_unsigned(652, 10), 1203 => to_unsigned(289, 10), 1204 => to_unsigned(1017, 10), 1205 => to_unsigned(521, 10), 1206 => to_unsigned(611, 10), 1207 => to_unsigned(760, 10), 1208 => to_unsigned(807, 10), 1209 => to_unsigned(837, 10), 1210 => to_unsigned(397, 10), 1211 => to_unsigned(75, 10), 1212 => to_unsigned(601, 10), 1213 => to_unsigned(747, 10), 1214 => to_unsigned(821, 10), 1215 => to_unsigned(673, 10), 1216 => to_unsigned(178, 10), 1217 => to_unsigned(796, 10), 1218 => to_unsigned(238, 10), 1219 => to_unsigned(538, 10), 1220 => to_unsigned(207, 10), 1221 => to_unsigned(770, 10), 1222 => to_unsigned(621, 10), 1223 => to_unsigned(986, 10), 1224 => to_unsigned(47, 10), 1225 => to_unsigned(582, 10), 1226 => to_unsigned(533, 10), 1227 => to_unsigned(265, 10), 1228 => to_unsigned(720, 10), 1229 => to_unsigned(549, 10), 1230 => to_unsigned(757, 10), 1231 => to_unsigned(535, 10), 1232 => to_unsigned(493, 10), 1233 => to_unsigned(602, 10), 1234 => to_unsigned(518, 10), 1235 => to_unsigned(706, 10), 1236 => to_unsigned(285, 10), 1237 => to_unsigned(805, 10), 1238 => to_unsigned(423, 10), 1239 => to_unsigned(25, 10), 1240 => to_unsigned(619, 10), 1241 => to_unsigned(432, 10), 1242 => to_unsigned(786, 10), 1243 => to_unsigned(442, 10), 1244 => to_unsigned(592, 10), 1245 => to_unsigned(946, 10), 1246 => to_unsigned(430, 10), 1247 => to_unsigned(849, 10), 1248 => to_unsigned(749, 10), 1249 => to_unsigned(638, 10), 1250 => to_unsigned(507, 10), 1251 => to_unsigned(400, 10), 1252 => to_unsigned(280, 10), 1253 => to_unsigned(812, 10), 1254 => to_unsigned(140, 10), 1255 => to_unsigned(169, 10), 1256 => to_unsigned(724, 10), 1257 => to_unsigned(58, 10), 1258 => to_unsigned(155, 10), 1259 => to_unsigned(272, 10), 1260 => to_unsigned(292, 10), 1261 => to_unsigned(479, 10), 1262 => to_unsigned(252, 10), 1263 => to_unsigned(268, 10), 1264 => to_unsigned(261, 10), 1265 => to_unsigned(269, 10), 1266 => to_unsigned(429, 10), 1267 => to_unsigned(873, 10), 1268 => to_unsigned(370, 10), 1269 => to_unsigned(994, 10), 1270 => to_unsigned(79, 10), 1271 => to_unsigned(113, 10), 1272 => to_unsigned(293, 10), 1273 => to_unsigned(547, 10), 1274 => to_unsigned(224, 10), 1275 => to_unsigned(104, 10), 1276 => to_unsigned(1023, 10), 1277 => to_unsigned(777, 10), 1278 => to_unsigned(367, 10), 1279 => to_unsigned(381, 10), 1280 => to_unsigned(40, 10), 1281 => to_unsigned(14, 10), 1282 => to_unsigned(771, 10), 1283 => to_unsigned(913, 10), 1284 => to_unsigned(427, 10), 1285 => to_unsigned(710, 10), 1286 => to_unsigned(983, 10), 1287 => to_unsigned(282, 10), 1288 => to_unsigned(300, 10), 1289 => to_unsigned(924, 10), 1290 => to_unsigned(229, 10), 1291 => to_unsigned(892, 10), 1292 => to_unsigned(650, 10), 1293 => to_unsigned(434, 10), 1294 => to_unsigned(253, 10), 1295 => to_unsigned(530, 10), 1296 => to_unsigned(492, 10), 1297 => to_unsigned(723, 10), 1298 => to_unsigned(861, 10), 1299 => to_unsigned(899, 10), 1300 => to_unsigned(772, 10), 1301 => to_unsigned(687, 10), 1302 => to_unsigned(686, 10), 1303 => to_unsigned(847, 10), 1304 => to_unsigned(976, 10), 1305 => to_unsigned(587, 10), 1306 => to_unsigned(941, 10), 1307 => to_unsigned(875, 10), 1308 => to_unsigned(779, 10), 1309 => to_unsigned(767, 10), 1310 => to_unsigned(639, 10), 1311 => to_unsigned(156, 10), 1312 => to_unsigned(2, 10), 1313 => to_unsigned(37, 10), 1314 => to_unsigned(327, 10), 1315 => to_unsigned(582, 10), 1316 => to_unsigned(492, 10), 1317 => to_unsigned(15, 10), 1318 => to_unsigned(603, 10), 1319 => to_unsigned(93, 10), 1320 => to_unsigned(739, 10), 1321 => to_unsigned(133, 10), 1322 => to_unsigned(516, 10), 1323 => to_unsigned(556, 10), 1324 => to_unsigned(998, 10), 1325 => to_unsigned(82, 10), 1326 => to_unsigned(761, 10), 1327 => to_unsigned(221, 10), 1328 => to_unsigned(270, 10), 1329 => to_unsigned(936, 10), 1330 => to_unsigned(90, 10), 1331 => to_unsigned(871, 10), 1332 => to_unsigned(34, 10), 1333 => to_unsigned(24, 10), 1334 => to_unsigned(395, 10), 1335 => to_unsigned(166, 10), 1336 => to_unsigned(52, 10), 1337 => to_unsigned(281, 10), 1338 => to_unsigned(692, 10), 1339 => to_unsigned(558, 10), 1340 => to_unsigned(440, 10), 1341 => to_unsigned(1001, 10), 1342 => to_unsigned(46, 10), 1343 => to_unsigned(190, 10), 1344 => to_unsigned(378, 10), 1345 => to_unsigned(958, 10), 1346 => to_unsigned(342, 10), 1347 => to_unsigned(936, 10), 1348 => to_unsigned(723, 10), 1349 => to_unsigned(1017, 10), 1350 => to_unsigned(892, 10), 1351 => to_unsigned(847, 10), 1352 => to_unsigned(902, 10), 1353 => to_unsigned(128, 10), 1354 => to_unsigned(890, 10), 1355 => to_unsigned(743, 10), 1356 => to_unsigned(865, 10), 1357 => to_unsigned(780, 10), 1358 => to_unsigned(97, 10), 1359 => to_unsigned(27, 10), 1360 => to_unsigned(924, 10), 1361 => to_unsigned(710, 10), 1362 => to_unsigned(750, 10), 1363 => to_unsigned(524, 10), 1364 => to_unsigned(887, 10), 1365 => to_unsigned(191, 10), 1366 => to_unsigned(800, 10), 1367 => to_unsigned(1009, 10), 1368 => to_unsigned(577, 10), 1369 => to_unsigned(998, 10), 1370 => to_unsigned(827, 10), 1371 => to_unsigned(401, 10), 1372 => to_unsigned(725, 10), 1373 => to_unsigned(882, 10), 1374 => to_unsigned(783, 10), 1375 => to_unsigned(630, 10), 1376 => to_unsigned(676, 10), 1377 => to_unsigned(1011, 10), 1378 => to_unsigned(91, 10), 1379 => to_unsigned(405, 10), 1380 => to_unsigned(820, 10), 1381 => to_unsigned(109, 10), 1382 => to_unsigned(63, 10), 1383 => to_unsigned(550, 10), 1384 => to_unsigned(226, 10), 1385 => to_unsigned(870, 10), 1386 => to_unsigned(469, 10), 1387 => to_unsigned(431, 10), 1388 => to_unsigned(443, 10), 1389 => to_unsigned(199, 10), 1390 => to_unsigned(294, 10), 1391 => to_unsigned(751, 10), 1392 => to_unsigned(342, 10), 1393 => to_unsigned(76, 10), 1394 => to_unsigned(272, 10), 1395 => to_unsigned(137, 10), 1396 => to_unsigned(746, 10), 1397 => to_unsigned(281, 10), 1398 => to_unsigned(93, 10), 1399 => to_unsigned(88, 10), 1400 => to_unsigned(159, 10), 1401 => to_unsigned(644, 10), 1402 => to_unsigned(8, 10), 1403 => to_unsigned(953, 10), 1404 => to_unsigned(882, 10), 1405 => to_unsigned(992, 10), 1406 => to_unsigned(716, 10), 1407 => to_unsigned(24, 10), 1408 => to_unsigned(539, 10), 1409 => to_unsigned(254, 10), 1410 => to_unsigned(531, 10), 1411 => to_unsigned(805, 10), 1412 => to_unsigned(201, 10), 1413 => to_unsigned(706, 10), 1414 => to_unsigned(491, 10), 1415 => to_unsigned(429, 10), 1416 => to_unsigned(846, 10), 1417 => to_unsigned(487, 10), 1418 => to_unsigned(283, 10), 1419 => to_unsigned(540, 10), 1420 => to_unsigned(782, 10), 1421 => to_unsigned(703, 10), 1422 => to_unsigned(369, 10), 1423 => to_unsigned(808, 10), 1424 => to_unsigned(575, 10), 1425 => to_unsigned(80, 10), 1426 => to_unsigned(876, 10), 1427 => to_unsigned(672, 10), 1428 => to_unsigned(1007, 10), 1429 => to_unsigned(583, 10), 1430 => to_unsigned(359, 10), 1431 => to_unsigned(494, 10), 1432 => to_unsigned(901, 10), 1433 => to_unsigned(991, 10), 1434 => to_unsigned(657, 10), 1435 => to_unsigned(628, 10), 1436 => to_unsigned(638, 10), 1437 => to_unsigned(239, 10), 1438 => to_unsigned(129, 10), 1439 => to_unsigned(358, 10), 1440 => to_unsigned(330, 10), 1441 => to_unsigned(603, 10), 1442 => to_unsigned(482, 10), 1443 => to_unsigned(929, 10), 1444 => to_unsigned(66, 10), 1445 => to_unsigned(1015, 10), 1446 => to_unsigned(542, 10), 1447 => to_unsigned(881, 10), 1448 => to_unsigned(111, 10), 1449 => to_unsigned(906, 10), 1450 => to_unsigned(774, 10), 1451 => to_unsigned(640, 10), 1452 => to_unsigned(395, 10), 1453 => to_unsigned(832, 10), 1454 => to_unsigned(951, 10), 1455 => to_unsigned(265, 10), 1456 => to_unsigned(530, 10), 1457 => to_unsigned(819, 10), 1458 => to_unsigned(76, 10), 1459 => to_unsigned(434, 10), 1460 => to_unsigned(562, 10), 1461 => to_unsigned(590, 10), 1462 => to_unsigned(745, 10), 1463 => to_unsigned(780, 10), 1464 => to_unsigned(993, 10), 1465 => to_unsigned(288, 10), 1466 => to_unsigned(281, 10), 1467 => to_unsigned(221, 10), 1468 => to_unsigned(407, 10), 1469 => to_unsigned(791, 10), 1470 => to_unsigned(940, 10), 1471 => to_unsigned(639, 10), 1472 => to_unsigned(602, 10), 1473 => to_unsigned(875, 10), 1474 => to_unsigned(741, 10), 1475 => to_unsigned(341, 10), 1476 => to_unsigned(691, 10), 1477 => to_unsigned(117, 10), 1478 => to_unsigned(227, 10), 1479 => to_unsigned(46, 10), 1480 => to_unsigned(141, 10), 1481 => to_unsigned(939, 10), 1482 => to_unsigned(910, 10), 1483 => to_unsigned(405, 10), 1484 => to_unsigned(252, 10), 1485 => to_unsigned(804, 10), 1486 => to_unsigned(751, 10), 1487 => to_unsigned(175, 10), 1488 => to_unsigned(277, 10), 1489 => to_unsigned(1001, 10), 1490 => to_unsigned(811, 10), 1491 => to_unsigned(239, 10), 1492 => to_unsigned(258, 10), 1493 => to_unsigned(515, 10), 1494 => to_unsigned(708, 10), 1495 => to_unsigned(165, 10), 1496 => to_unsigned(545, 10), 1497 => to_unsigned(925, 10), 1498 => to_unsigned(494, 10), 1499 => to_unsigned(171, 10), 1500 => to_unsigned(340, 10), 1501 => to_unsigned(806, 10), 1502 => to_unsigned(168, 10), 1503 => to_unsigned(460, 10), 1504 => to_unsigned(131, 10), 1505 => to_unsigned(851, 10), 1506 => to_unsigned(952, 10), 1507 => to_unsigned(215, 10), 1508 => to_unsigned(919, 10), 1509 => to_unsigned(732, 10), 1510 => to_unsigned(770, 10), 1511 => to_unsigned(199, 10), 1512 => to_unsigned(605, 10), 1513 => to_unsigned(72, 10), 1514 => to_unsigned(228, 10), 1515 => to_unsigned(946, 10), 1516 => to_unsigned(96, 10), 1517 => to_unsigned(983, 10), 1518 => to_unsigned(330, 10), 1519 => to_unsigned(788, 10), 1520 => to_unsigned(237, 10), 1521 => to_unsigned(83, 10), 1522 => to_unsigned(72, 10), 1523 => to_unsigned(79, 10), 1524 => to_unsigned(937, 10), 1525 => to_unsigned(892, 10), 1526 => to_unsigned(694, 10), 1527 => to_unsigned(680, 10), 1528 => to_unsigned(1003, 10), 1529 => to_unsigned(485, 10), 1530 => to_unsigned(320, 10), 1531 => to_unsigned(723, 10), 1532 => to_unsigned(215, 10), 1533 => to_unsigned(70, 10), 1534 => to_unsigned(84, 10), 1535 => to_unsigned(125, 10), 1536 => to_unsigned(902, 10), 1537 => to_unsigned(868, 10), 1538 => to_unsigned(495, 10), 1539 => to_unsigned(450, 10), 1540 => to_unsigned(274, 10), 1541 => to_unsigned(983, 10), 1542 => to_unsigned(799, 10), 1543 => to_unsigned(972, 10), 1544 => to_unsigned(51, 10), 1545 => to_unsigned(566, 10), 1546 => to_unsigned(793, 10), 1547 => to_unsigned(153, 10), 1548 => to_unsigned(1018, 10), 1549 => to_unsigned(516, 10), 1550 => to_unsigned(750, 10), 1551 => to_unsigned(22, 10), 1552 => to_unsigned(438, 10), 1553 => to_unsigned(881, 10), 1554 => to_unsigned(98, 10), 1555 => to_unsigned(985, 10), 1556 => to_unsigned(423, 10), 1557 => to_unsigned(426, 10), 1558 => to_unsigned(226, 10), 1559 => to_unsigned(824, 10), 1560 => to_unsigned(278, 10), 1561 => to_unsigned(325, 10), 1562 => to_unsigned(194, 10), 1563 => to_unsigned(1003, 10), 1564 => to_unsigned(242, 10), 1565 => to_unsigned(253, 10), 1566 => to_unsigned(987, 10), 1567 => to_unsigned(521, 10), 1568 => to_unsigned(82, 10), 1569 => to_unsigned(282, 10), 1570 => to_unsigned(103, 10), 1571 => to_unsigned(262, 10), 1572 => to_unsigned(269, 10), 1573 => to_unsigned(976, 10), 1574 => to_unsigned(352, 10), 1575 => to_unsigned(698, 10), 1576 => to_unsigned(857, 10), 1577 => to_unsigned(667, 10), 1578 => to_unsigned(280, 10), 1579 => to_unsigned(440, 10), 1580 => to_unsigned(214, 10), 1581 => to_unsigned(76, 10), 1582 => to_unsigned(668, 10), 1583 => to_unsigned(908, 10), 1584 => to_unsigned(580, 10), 1585 => to_unsigned(137, 10), 1586 => to_unsigned(72, 10), 1587 => to_unsigned(441, 10), 1588 => to_unsigned(486, 10), 1589 => to_unsigned(117, 10), 1590 => to_unsigned(802, 10), 1591 => to_unsigned(41, 10), 1592 => to_unsigned(64, 10), 1593 => to_unsigned(784, 10), 1594 => to_unsigned(345, 10), 1595 => to_unsigned(687, 10), 1596 => to_unsigned(851, 10), 1597 => to_unsigned(670, 10), 1598 => to_unsigned(546, 10), 1599 => to_unsigned(570, 10), 1600 => to_unsigned(743, 10), 1601 => to_unsigned(101, 10), 1602 => to_unsigned(661, 10), 1603 => to_unsigned(824, 10), 1604 => to_unsigned(584, 10), 1605 => to_unsigned(708, 10), 1606 => to_unsigned(970, 10), 1607 => to_unsigned(139, 10), 1608 => to_unsigned(763, 10), 1609 => to_unsigned(5, 10), 1610 => to_unsigned(944, 10), 1611 => to_unsigned(327, 10), 1612 => to_unsigned(891, 10), 1613 => to_unsigned(359, 10), 1614 => to_unsigned(192, 10), 1615 => to_unsigned(804, 10), 1616 => to_unsigned(286, 10), 1617 => to_unsigned(836, 10), 1618 => to_unsigned(385, 10), 1619 => to_unsigned(338, 10), 1620 => to_unsigned(62, 10), 1621 => to_unsigned(370, 10), 1622 => to_unsigned(668, 10), 1623 => to_unsigned(561, 10), 1624 => to_unsigned(963, 10), 1625 => to_unsigned(892, 10), 1626 => to_unsigned(286, 10), 1627 => to_unsigned(549, 10), 1628 => to_unsigned(790, 10), 1629 => to_unsigned(1015, 10), 1630 => to_unsigned(480, 10), 1631 => to_unsigned(125, 10), 1632 => to_unsigned(1002, 10), 1633 => to_unsigned(1004, 10), 1634 => to_unsigned(594, 10), 1635 => to_unsigned(508, 10), 1636 => to_unsigned(555, 10), 1637 => to_unsigned(116, 10), 1638 => to_unsigned(314, 10), 1639 => to_unsigned(907, 10), 1640 => to_unsigned(570, 10), 1641 => to_unsigned(244, 10), 1642 => to_unsigned(602, 10), 1643 => to_unsigned(517, 10), 1644 => to_unsigned(83, 10), 1645 => to_unsigned(470, 10), 1646 => to_unsigned(1006, 10), 1647 => to_unsigned(510, 10), 1648 => to_unsigned(696, 10), 1649 => to_unsigned(634, 10), 1650 => to_unsigned(836, 10), 1651 => to_unsigned(219, 10), 1652 => to_unsigned(813, 10), 1653 => to_unsigned(333, 10), 1654 => to_unsigned(197, 10), 1655 => to_unsigned(1006, 10), 1656 => to_unsigned(258, 10), 1657 => to_unsigned(169, 10), 1658 => to_unsigned(562, 10), 1659 => to_unsigned(829, 10), 1660 => to_unsigned(344, 10), 1661 => to_unsigned(173, 10), 1662 => to_unsigned(955, 10), 1663 => to_unsigned(429, 10), 1664 => to_unsigned(989, 10), 1665 => to_unsigned(668, 10), 1666 => to_unsigned(837, 10), 1667 => to_unsigned(737, 10), 1668 => to_unsigned(921, 10), 1669 => to_unsigned(736, 10), 1670 => to_unsigned(732, 10), 1671 => to_unsigned(605, 10), 1672 => to_unsigned(363, 10), 1673 => to_unsigned(201, 10), 1674 => to_unsigned(69, 10), 1675 => to_unsigned(1018, 10), 1676 => to_unsigned(916, 10), 1677 => to_unsigned(344, 10), 1678 => to_unsigned(766, 10), 1679 => to_unsigned(476, 10), 1680 => to_unsigned(536, 10), 1681 => to_unsigned(245, 10), 1682 => to_unsigned(785, 10), 1683 => to_unsigned(172, 10), 1684 => to_unsigned(322, 10), 1685 => to_unsigned(283, 10), 1686 => to_unsigned(25, 10), 1687 => to_unsigned(698, 10), 1688 => to_unsigned(144, 10), 1689 => to_unsigned(32, 10), 1690 => to_unsigned(614, 10), 1691 => to_unsigned(94, 10), 1692 => to_unsigned(47, 10), 1693 => to_unsigned(261, 10), 1694 => to_unsigned(40, 10), 1695 => to_unsigned(146, 10), 1696 => to_unsigned(794, 10), 1697 => to_unsigned(356, 10), 1698 => to_unsigned(175, 10), 1699 => to_unsigned(887, 10), 1700 => to_unsigned(498, 10), 1701 => to_unsigned(795, 10), 1702 => to_unsigned(814, 10), 1703 => to_unsigned(242, 10), 1704 => to_unsigned(675, 10), 1705 => to_unsigned(663, 10), 1706 => to_unsigned(312, 10), 1707 => to_unsigned(138, 10), 1708 => to_unsigned(948, 10), 1709 => to_unsigned(636, 10), 1710 => to_unsigned(639, 10), 1711 => to_unsigned(442, 10), 1712 => to_unsigned(394, 10), 1713 => to_unsigned(707, 10), 1714 => to_unsigned(11, 10), 1715 => to_unsigned(8, 10), 1716 => to_unsigned(1015, 10), 1717 => to_unsigned(145, 10), 1718 => to_unsigned(973, 10), 1719 => to_unsigned(853, 10), 1720 => to_unsigned(936, 10), 1721 => to_unsigned(9, 10), 1722 => to_unsigned(650, 10), 1723 => to_unsigned(662, 10), 1724 => to_unsigned(477, 10), 1725 => to_unsigned(470, 10), 1726 => to_unsigned(361, 10), 1727 => to_unsigned(733, 10), 1728 => to_unsigned(126, 10), 1729 => to_unsigned(609, 10), 1730 => to_unsigned(586, 10), 1731 => to_unsigned(199, 10), 1732 => to_unsigned(718, 10), 1733 => to_unsigned(106, 10), 1734 => to_unsigned(694, 10), 1735 => to_unsigned(99, 10), 1736 => to_unsigned(70, 10), 1737 => to_unsigned(408, 10), 1738 => to_unsigned(890, 10), 1739 => to_unsigned(875, 10), 1740 => to_unsigned(328, 10), 1741 => to_unsigned(435, 10), 1742 => to_unsigned(258, 10), 1743 => to_unsigned(167, 10), 1744 => to_unsigned(430, 10), 1745 => to_unsigned(809, 10), 1746 => to_unsigned(909, 10), 1747 => to_unsigned(788, 10), 1748 => to_unsigned(65, 10), 1749 => to_unsigned(850, 10), 1750 => to_unsigned(332, 10), 1751 => to_unsigned(385, 10), 1752 => to_unsigned(649, 10), 1753 => to_unsigned(598, 10), 1754 => to_unsigned(386, 10), 1755 => to_unsigned(572, 10), 1756 => to_unsigned(441, 10), 1757 => to_unsigned(204, 10), 1758 => to_unsigned(277, 10), 1759 => to_unsigned(218, 10), 1760 => to_unsigned(6, 10), 1761 => to_unsigned(164, 10), 1762 => to_unsigned(898, 10), 1763 => to_unsigned(316, 10), 1764 => to_unsigned(698, 10), 1765 => to_unsigned(357, 10), 1766 => to_unsigned(64, 10), 1767 => to_unsigned(908, 10), 1768 => to_unsigned(48, 10), 1769 => to_unsigned(941, 10), 1770 => to_unsigned(786, 10), 1771 => to_unsigned(292, 10), 1772 => to_unsigned(1018, 10), 1773 => to_unsigned(505, 10), 1774 => to_unsigned(112, 10), 1775 => to_unsigned(864, 10), 1776 => to_unsigned(881, 10), 1777 => to_unsigned(366, 10), 1778 => to_unsigned(777, 10), 1779 => to_unsigned(35, 10), 1780 => to_unsigned(124, 10), 1781 => to_unsigned(31, 10), 1782 => to_unsigned(251, 10), 1783 => to_unsigned(630, 10), 1784 => to_unsigned(922, 10), 1785 => to_unsigned(586, 10), 1786 => to_unsigned(402, 10), 1787 => to_unsigned(957, 10), 1788 => to_unsigned(767, 10), 1789 => to_unsigned(265, 10), 1790 => to_unsigned(786, 10), 1791 => to_unsigned(917, 10), 1792 => to_unsigned(176, 10), 1793 => to_unsigned(17, 10), 1794 => to_unsigned(1005, 10), 1795 => to_unsigned(724, 10), 1796 => to_unsigned(882, 10), 1797 => to_unsigned(589, 10), 1798 => to_unsigned(155, 10), 1799 => to_unsigned(243, 10), 1800 => to_unsigned(439, 10), 1801 => to_unsigned(103, 10), 1802 => to_unsigned(1014, 10), 1803 => to_unsigned(233, 10), 1804 => to_unsigned(95, 10), 1805 => to_unsigned(215, 10), 1806 => to_unsigned(725, 10), 1807 => to_unsigned(78, 10), 1808 => to_unsigned(98, 10), 1809 => to_unsigned(148, 10), 1810 => to_unsigned(286, 10), 1811 => to_unsigned(596, 10), 1812 => to_unsigned(454, 10), 1813 => to_unsigned(957, 10), 1814 => to_unsigned(739, 10), 1815 => to_unsigned(686, 10), 1816 => to_unsigned(949, 10), 1817 => to_unsigned(5, 10), 1818 => to_unsigned(406, 10), 1819 => to_unsigned(941, 10), 1820 => to_unsigned(820, 10), 1821 => to_unsigned(766, 10), 1822 => to_unsigned(340, 10), 1823 => to_unsigned(40, 10), 1824 => to_unsigned(830, 10), 1825 => to_unsigned(242, 10), 1826 => to_unsigned(175, 10), 1827 => to_unsigned(947, 10), 1828 => to_unsigned(531, 10), 1829 => to_unsigned(301, 10), 1830 => to_unsigned(917, 10), 1831 => to_unsigned(677, 10), 1832 => to_unsigned(724, 10), 1833 => to_unsigned(1011, 10), 1834 => to_unsigned(439, 10), 1835 => to_unsigned(151, 10), 1836 => to_unsigned(217, 10), 1837 => to_unsigned(409, 10), 1838 => to_unsigned(590, 10), 1839 => to_unsigned(120, 10), 1840 => to_unsigned(79, 10), 1841 => to_unsigned(311, 10), 1842 => to_unsigned(301, 10), 1843 => to_unsigned(656, 10), 1844 => to_unsigned(509, 10), 1845 => to_unsigned(254, 10), 1846 => to_unsigned(904, 10), 1847 => to_unsigned(970, 10), 1848 => to_unsigned(618, 10), 1849 => to_unsigned(405, 10), 1850 => to_unsigned(784, 10), 1851 => to_unsigned(350, 10), 1852 => to_unsigned(956, 10), 1853 => to_unsigned(406, 10), 1854 => to_unsigned(620, 10), 1855 => to_unsigned(601, 10), 1856 => to_unsigned(795, 10), 1857 => to_unsigned(937, 10), 1858 => to_unsigned(467, 10), 1859 => to_unsigned(30, 10), 1860 => to_unsigned(1019, 10), 1861 => to_unsigned(170, 10), 1862 => to_unsigned(570, 10), 1863 => to_unsigned(871, 10), 1864 => to_unsigned(417, 10), 1865 => to_unsigned(405, 10), 1866 => to_unsigned(970, 10), 1867 => to_unsigned(132, 10), 1868 => to_unsigned(616, 10), 1869 => to_unsigned(802, 10), 1870 => to_unsigned(116, 10), 1871 => to_unsigned(151, 10), 1872 => to_unsigned(576, 10), 1873 => to_unsigned(336, 10), 1874 => to_unsigned(1002, 10), 1875 => to_unsigned(846, 10), 1876 => to_unsigned(961, 10), 1877 => to_unsigned(201, 10), 1878 => to_unsigned(485, 10), 1879 => to_unsigned(19, 10), 1880 => to_unsigned(320, 10), 1881 => to_unsigned(131, 10), 1882 => to_unsigned(941, 10), 1883 => to_unsigned(425, 10), 1884 => to_unsigned(811, 10), 1885 => to_unsigned(631, 10), 1886 => to_unsigned(793, 10), 1887 => to_unsigned(705, 10), 1888 => to_unsigned(48, 10), 1889 => to_unsigned(280, 10), 1890 => to_unsigned(385, 10), 1891 => to_unsigned(907, 10), 1892 => to_unsigned(943, 10), 1893 => to_unsigned(335, 10), 1894 => to_unsigned(663, 10), 1895 => to_unsigned(734, 10), 1896 => to_unsigned(310, 10), 1897 => to_unsigned(660, 10), 1898 => to_unsigned(996, 10), 1899 => to_unsigned(514, 10), 1900 => to_unsigned(619, 10), 1901 => to_unsigned(312, 10), 1902 => to_unsigned(855, 10), 1903 => to_unsigned(489, 10), 1904 => to_unsigned(605, 10), 1905 => to_unsigned(433, 10), 1906 => to_unsigned(699, 10), 1907 => to_unsigned(802, 10), 1908 => to_unsigned(420, 10), 1909 => to_unsigned(349, 10), 1910 => to_unsigned(259, 10), 1911 => to_unsigned(571, 10), 1912 => to_unsigned(411, 10), 1913 => to_unsigned(723, 10), 1914 => to_unsigned(803, 10), 1915 => to_unsigned(772, 10), 1916 => to_unsigned(860, 10), 1917 => to_unsigned(819, 10), 1918 => to_unsigned(139, 10), 1919 => to_unsigned(878, 10), 1920 => to_unsigned(265, 10), 1921 => to_unsigned(204, 10), 1922 => to_unsigned(917, 10), 1923 => to_unsigned(285, 10), 1924 => to_unsigned(433, 10), 1925 => to_unsigned(241, 10), 1926 => to_unsigned(707, 10), 1927 => to_unsigned(710, 10), 1928 => to_unsigned(851, 10), 1929 => to_unsigned(24, 10), 1930 => to_unsigned(157, 10), 1931 => to_unsigned(410, 10), 1932 => to_unsigned(590, 10), 1933 => to_unsigned(953, 10), 1934 => to_unsigned(867, 10), 1935 => to_unsigned(741, 10), 1936 => to_unsigned(177, 10), 1937 => to_unsigned(365, 10), 1938 => to_unsigned(331, 10), 1939 => to_unsigned(897, 10), 1940 => to_unsigned(641, 10), 1941 => to_unsigned(546, 10), 1942 => to_unsigned(878, 10), 1943 => to_unsigned(1003, 10), 1944 => to_unsigned(82, 10), 1945 => to_unsigned(1014, 10), 1946 => to_unsigned(980, 10), 1947 => to_unsigned(297, 10), 1948 => to_unsigned(774, 10), 1949 => to_unsigned(808, 10), 1950 => to_unsigned(343, 10), 1951 => to_unsigned(228, 10), 1952 => to_unsigned(728, 10), 1953 => to_unsigned(24, 10), 1954 => to_unsigned(626, 10), 1955 => to_unsigned(622, 10), 1956 => to_unsigned(224, 10), 1957 => to_unsigned(726, 10), 1958 => to_unsigned(274, 10), 1959 => to_unsigned(655, 10), 1960 => to_unsigned(167, 10), 1961 => to_unsigned(602, 10), 1962 => to_unsigned(435, 10), 1963 => to_unsigned(615, 10), 1964 => to_unsigned(329, 10), 1965 => to_unsigned(900, 10), 1966 => to_unsigned(577, 10), 1967 => to_unsigned(26, 10), 1968 => to_unsigned(221, 10), 1969 => to_unsigned(927, 10), 1970 => to_unsigned(605, 10), 1971 => to_unsigned(549, 10), 1972 => to_unsigned(530, 10), 1973 => to_unsigned(347, 10), 1974 => to_unsigned(47, 10), 1975 => to_unsigned(800, 10), 1976 => to_unsigned(369, 10), 1977 => to_unsigned(567, 10), 1978 => to_unsigned(11, 10), 1979 => to_unsigned(699, 10), 1980 => to_unsigned(410, 10), 1981 => to_unsigned(188, 10), 1982 => to_unsigned(961, 10), 1983 => to_unsigned(229, 10), 1984 => to_unsigned(449, 10), 1985 => to_unsigned(167, 10), 1986 => to_unsigned(1015, 10), 1987 => to_unsigned(396, 10), 1988 => to_unsigned(348, 10), 1989 => to_unsigned(917, 10), 1990 => to_unsigned(987, 10), 1991 => to_unsigned(902, 10), 1992 => to_unsigned(624, 10), 1993 => to_unsigned(341, 10), 1994 => to_unsigned(150, 10), 1995 => to_unsigned(855, 10), 1996 => to_unsigned(544, 10), 1997 => to_unsigned(984, 10), 1998 => to_unsigned(98, 10), 1999 => to_unsigned(671, 10), 2000 => to_unsigned(288, 10), 2001 => to_unsigned(236, 10), 2002 => to_unsigned(157, 10), 2003 => to_unsigned(294, 10), 2004 => to_unsigned(382, 10), 2005 => to_unsigned(568, 10), 2006 => to_unsigned(80, 10), 2007 => to_unsigned(580, 10), 2008 => to_unsigned(962, 10), 2009 => to_unsigned(174, 10), 2010 => to_unsigned(414, 10), 2011 => to_unsigned(221, 10), 2012 => to_unsigned(39, 10), 2013 => to_unsigned(1002, 10), 2014 => to_unsigned(649, 10), 2015 => to_unsigned(567, 10), 2016 => to_unsigned(602, 10), 2017 => to_unsigned(198, 10), 2018 => to_unsigned(165, 10), 2019 => to_unsigned(217, 10), 2020 => to_unsigned(682, 10), 2021 => to_unsigned(564, 10), 2022 => to_unsigned(982, 10), 2023 => to_unsigned(890, 10), 2024 => to_unsigned(126, 10), 2025 => to_unsigned(450, 10), 2026 => to_unsigned(417, 10), 2027 => to_unsigned(435, 10), 2028 => to_unsigned(696, 10), 2029 => to_unsigned(778, 10), 2030 => to_unsigned(818, 10), 2031 => to_unsigned(355, 10), 2032 => to_unsigned(291, 10), 2033 => to_unsigned(769, 10), 2034 => to_unsigned(214, 10), 2035 => to_unsigned(590, 10), 2036 => to_unsigned(441, 10), 2037 => to_unsigned(289, 10), 2038 => to_unsigned(840, 10), 2039 => to_unsigned(918, 10), 2040 => to_unsigned(875, 10), 2041 => to_unsigned(575, 10), 2042 => to_unsigned(449, 10), 2043 => to_unsigned(179, 10), 2044 => to_unsigned(288, 10), 2045 => to_unsigned(490, 10), 2046 => to_unsigned(163, 10), 2047 => to_unsigned(832, 10)),
            5 => (0 => to_unsigned(84, 10), 1 => to_unsigned(957, 10), 2 => to_unsigned(537, 10), 3 => to_unsigned(83, 10), 4 => to_unsigned(1, 10), 5 => to_unsigned(54, 10), 6 => to_unsigned(859, 10), 7 => to_unsigned(100, 10), 8 => to_unsigned(704, 10), 9 => to_unsigned(586, 10), 10 => to_unsigned(560, 10), 11 => to_unsigned(962, 10), 12 => to_unsigned(268, 10), 13 => to_unsigned(958, 10), 14 => to_unsigned(437, 10), 15 => to_unsigned(588, 10), 16 => to_unsigned(208, 10), 17 => to_unsigned(503, 10), 18 => to_unsigned(323, 10), 19 => to_unsigned(634, 10), 20 => to_unsigned(809, 10), 21 => to_unsigned(718, 10), 22 => to_unsigned(1009, 10), 23 => to_unsigned(887, 10), 24 => to_unsigned(628, 10), 25 => to_unsigned(255, 10), 26 => to_unsigned(1001, 10), 27 => to_unsigned(725, 10), 28 => to_unsigned(972, 10), 29 => to_unsigned(241, 10), 30 => to_unsigned(861, 10), 31 => to_unsigned(376, 10), 32 => to_unsigned(908, 10), 33 => to_unsigned(58, 10), 34 => to_unsigned(201, 10), 35 => to_unsigned(475, 10), 36 => to_unsigned(225, 10), 37 => to_unsigned(293, 10), 38 => to_unsigned(46, 10), 39 => to_unsigned(699, 10), 40 => to_unsigned(335, 10), 41 => to_unsigned(722, 10), 42 => to_unsigned(123, 10), 43 => to_unsigned(485, 10), 44 => to_unsigned(617, 10), 45 => to_unsigned(370, 10), 46 => to_unsigned(1007, 10), 47 => to_unsigned(167, 10), 48 => to_unsigned(780, 10), 49 => to_unsigned(537, 10), 50 => to_unsigned(806, 10), 51 => to_unsigned(259, 10), 52 => to_unsigned(4, 10), 53 => to_unsigned(671, 10), 54 => to_unsigned(871, 10), 55 => to_unsigned(341, 10), 56 => to_unsigned(961, 10), 57 => to_unsigned(439, 10), 58 => to_unsigned(122, 10), 59 => to_unsigned(711, 10), 60 => to_unsigned(238, 10), 61 => to_unsigned(511, 10), 62 => to_unsigned(528, 10), 63 => to_unsigned(71, 10), 64 => to_unsigned(77, 10), 65 => to_unsigned(506, 10), 66 => to_unsigned(873, 10), 67 => to_unsigned(217, 10), 68 => to_unsigned(971, 10), 69 => to_unsigned(509, 10), 70 => to_unsigned(99, 10), 71 => to_unsigned(441, 10), 72 => to_unsigned(894, 10), 73 => to_unsigned(509, 10), 74 => to_unsigned(66, 10), 75 => to_unsigned(77, 10), 76 => to_unsigned(515, 10), 77 => to_unsigned(971, 10), 78 => to_unsigned(385, 10), 79 => to_unsigned(480, 10), 80 => to_unsigned(323, 10), 81 => to_unsigned(648, 10), 82 => to_unsigned(177, 10), 83 => to_unsigned(520, 10), 84 => to_unsigned(805, 10), 85 => to_unsigned(106, 10), 86 => to_unsigned(817, 10), 87 => to_unsigned(769, 10), 88 => to_unsigned(342, 10), 89 => to_unsigned(69, 10), 90 => to_unsigned(683, 10), 91 => to_unsigned(873, 10), 92 => to_unsigned(299, 10), 93 => to_unsigned(676, 10), 94 => to_unsigned(873, 10), 95 => to_unsigned(296, 10), 96 => to_unsigned(676, 10), 97 => to_unsigned(820, 10), 98 => to_unsigned(498, 10), 99 => to_unsigned(845, 10), 100 => to_unsigned(37, 10), 101 => to_unsigned(685, 10), 102 => to_unsigned(41, 10), 103 => to_unsigned(825, 10), 104 => to_unsigned(200, 10), 105 => to_unsigned(89, 10), 106 => to_unsigned(280, 10), 107 => to_unsigned(901, 10), 108 => to_unsigned(5, 10), 109 => to_unsigned(420, 10), 110 => to_unsigned(357, 10), 111 => to_unsigned(260, 10), 112 => to_unsigned(591, 10), 113 => to_unsigned(442, 10), 114 => to_unsigned(711, 10), 115 => to_unsigned(407, 10), 116 => to_unsigned(674, 10), 117 => to_unsigned(969, 10), 118 => to_unsigned(521, 10), 119 => to_unsigned(440, 10), 120 => to_unsigned(174, 10), 121 => to_unsigned(547, 10), 122 => to_unsigned(863, 10), 123 => to_unsigned(959, 10), 124 => to_unsigned(968, 10), 125 => to_unsigned(562, 10), 126 => to_unsigned(455, 10), 127 => to_unsigned(56, 10), 128 => to_unsigned(453, 10), 129 => to_unsigned(351, 10), 130 => to_unsigned(911, 10), 131 => to_unsigned(984, 10), 132 => to_unsigned(854, 10), 133 => to_unsigned(511, 10), 134 => to_unsigned(6, 10), 135 => to_unsigned(38, 10), 136 => to_unsigned(368, 10), 137 => to_unsigned(744, 10), 138 => to_unsigned(589, 10), 139 => to_unsigned(1017, 10), 140 => to_unsigned(274, 10), 141 => to_unsigned(452, 10), 142 => to_unsigned(388, 10), 143 => to_unsigned(510, 10), 144 => to_unsigned(1012, 10), 145 => to_unsigned(246, 10), 146 => to_unsigned(966, 10), 147 => to_unsigned(105, 10), 148 => to_unsigned(894, 10), 149 => to_unsigned(460, 10), 150 => to_unsigned(68, 10), 151 => to_unsigned(939, 10), 152 => to_unsigned(153, 10), 153 => to_unsigned(576, 10), 154 => to_unsigned(85, 10), 155 => to_unsigned(251, 10), 156 => to_unsigned(644, 10), 157 => to_unsigned(190, 10), 158 => to_unsigned(1020, 10), 159 => to_unsigned(804, 10), 160 => to_unsigned(292, 10), 161 => to_unsigned(626, 10), 162 => to_unsigned(188, 10), 163 => to_unsigned(26, 10), 164 => to_unsigned(830, 10), 165 => to_unsigned(190, 10), 166 => to_unsigned(669, 10), 167 => to_unsigned(872, 10), 168 => to_unsigned(414, 10), 169 => to_unsigned(207, 10), 170 => to_unsigned(195, 10), 171 => to_unsigned(340, 10), 172 => to_unsigned(1015, 10), 173 => to_unsigned(630, 10), 174 => to_unsigned(722, 10), 175 => to_unsigned(103, 10), 176 => to_unsigned(830, 10), 177 => to_unsigned(696, 10), 178 => to_unsigned(653, 10), 179 => to_unsigned(535, 10), 180 => to_unsigned(412, 10), 181 => to_unsigned(508, 10), 182 => to_unsigned(91, 10), 183 => to_unsigned(105, 10), 184 => to_unsigned(592, 10), 185 => to_unsigned(754, 10), 186 => to_unsigned(1023, 10), 187 => to_unsigned(261, 10), 188 => to_unsigned(450, 10), 189 => to_unsigned(57, 10), 190 => to_unsigned(780, 10), 191 => to_unsigned(644, 10), 192 => to_unsigned(21, 10), 193 => to_unsigned(193, 10), 194 => to_unsigned(507, 10), 195 => to_unsigned(757, 10), 196 => to_unsigned(923, 10), 197 => to_unsigned(158, 10), 198 => to_unsigned(101, 10), 199 => to_unsigned(1008, 10), 200 => to_unsigned(323, 10), 201 => to_unsigned(384, 10), 202 => to_unsigned(39, 10), 203 => to_unsigned(200, 10), 204 => to_unsigned(478, 10), 205 => to_unsigned(625, 10), 206 => to_unsigned(172, 10), 207 => to_unsigned(547, 10), 208 => to_unsigned(780, 10), 209 => to_unsigned(452, 10), 210 => to_unsigned(216, 10), 211 => to_unsigned(445, 10), 212 => to_unsigned(345, 10), 213 => to_unsigned(548, 10), 214 => to_unsigned(67, 10), 215 => to_unsigned(951, 10), 216 => to_unsigned(516, 10), 217 => to_unsigned(109, 10), 218 => to_unsigned(995, 10), 219 => to_unsigned(380, 10), 220 => to_unsigned(770, 10), 221 => to_unsigned(596, 10), 222 => to_unsigned(804, 10), 223 => to_unsigned(468, 10), 224 => to_unsigned(141, 10), 225 => to_unsigned(544, 10), 226 => to_unsigned(796, 10), 227 => to_unsigned(168, 10), 228 => to_unsigned(295, 10), 229 => to_unsigned(897, 10), 230 => to_unsigned(481, 10), 231 => to_unsigned(579, 10), 232 => to_unsigned(293, 10), 233 => to_unsigned(193, 10), 234 => to_unsigned(351, 10), 235 => to_unsigned(707, 10), 236 => to_unsigned(488, 10), 237 => to_unsigned(899, 10), 238 => to_unsigned(803, 10), 239 => to_unsigned(226, 10), 240 => to_unsigned(90, 10), 241 => to_unsigned(678, 10), 242 => to_unsigned(303, 10), 243 => to_unsigned(888, 10), 244 => to_unsigned(218, 10), 245 => to_unsigned(376, 10), 246 => to_unsigned(678, 10), 247 => to_unsigned(961, 10), 248 => to_unsigned(97, 10), 249 => to_unsigned(563, 10), 250 => to_unsigned(94, 10), 251 => to_unsigned(886, 10), 252 => to_unsigned(783, 10), 253 => to_unsigned(876, 10), 254 => to_unsigned(1014, 10), 255 => to_unsigned(869, 10), 256 => to_unsigned(190, 10), 257 => to_unsigned(427, 10), 258 => to_unsigned(357, 10), 259 => to_unsigned(614, 10), 260 => to_unsigned(378, 10), 261 => to_unsigned(666, 10), 262 => to_unsigned(948, 10), 263 => to_unsigned(175, 10), 264 => to_unsigned(448, 10), 265 => to_unsigned(1022, 10), 266 => to_unsigned(304, 10), 267 => to_unsigned(642, 10), 268 => to_unsigned(740, 10), 269 => to_unsigned(183, 10), 270 => to_unsigned(170, 10), 271 => to_unsigned(206, 10), 272 => to_unsigned(472, 10), 273 => to_unsigned(895, 10), 274 => to_unsigned(594, 10), 275 => to_unsigned(104, 10), 276 => to_unsigned(6, 10), 277 => to_unsigned(515, 10), 278 => to_unsigned(862, 10), 279 => to_unsigned(622, 10), 280 => to_unsigned(950, 10), 281 => to_unsigned(78, 10), 282 => to_unsigned(479, 10), 283 => to_unsigned(790, 10), 284 => to_unsigned(784, 10), 285 => to_unsigned(529, 10), 286 => to_unsigned(394, 10), 287 => to_unsigned(657, 10), 288 => to_unsigned(701, 10), 289 => to_unsigned(581, 10), 290 => to_unsigned(568, 10), 291 => to_unsigned(663, 10), 292 => to_unsigned(891, 10), 293 => to_unsigned(227, 10), 294 => to_unsigned(313, 10), 295 => to_unsigned(178, 10), 296 => to_unsigned(643, 10), 297 => to_unsigned(941, 10), 298 => to_unsigned(894, 10), 299 => to_unsigned(283, 10), 300 => to_unsigned(702, 10), 301 => to_unsigned(900, 10), 302 => to_unsigned(517, 10), 303 => to_unsigned(628, 10), 304 => to_unsigned(498, 10), 305 => to_unsigned(169, 10), 306 => to_unsigned(502, 10), 307 => to_unsigned(618, 10), 308 => to_unsigned(650, 10), 309 => to_unsigned(191, 10), 310 => to_unsigned(860, 10), 311 => to_unsigned(567, 10), 312 => to_unsigned(12, 10), 313 => to_unsigned(945, 10), 314 => to_unsigned(945, 10), 315 => to_unsigned(227, 10), 316 => to_unsigned(931, 10), 317 => to_unsigned(736, 10), 318 => to_unsigned(588, 10), 319 => to_unsigned(231, 10), 320 => to_unsigned(944, 10), 321 => to_unsigned(86, 10), 322 => to_unsigned(467, 10), 323 => to_unsigned(630, 10), 324 => to_unsigned(659, 10), 325 => to_unsigned(961, 10), 326 => to_unsigned(899, 10), 327 => to_unsigned(193, 10), 328 => to_unsigned(221, 10), 329 => to_unsigned(98, 10), 330 => to_unsigned(169, 10), 331 => to_unsigned(898, 10), 332 => to_unsigned(810, 10), 333 => to_unsigned(72, 10), 334 => to_unsigned(361, 10), 335 => to_unsigned(4, 10), 336 => to_unsigned(170, 10), 337 => to_unsigned(830, 10), 338 => to_unsigned(721, 10), 339 => to_unsigned(954, 10), 340 => to_unsigned(915, 10), 341 => to_unsigned(53, 10), 342 => to_unsigned(844, 10), 343 => to_unsigned(10, 10), 344 => to_unsigned(761, 10), 345 => to_unsigned(125, 10), 346 => to_unsigned(632, 10), 347 => to_unsigned(708, 10), 348 => to_unsigned(891, 10), 349 => to_unsigned(6, 10), 350 => to_unsigned(261, 10), 351 => to_unsigned(284, 10), 352 => to_unsigned(201, 10), 353 => to_unsigned(224, 10), 354 => to_unsigned(108, 10), 355 => to_unsigned(945, 10), 356 => to_unsigned(826, 10), 357 => to_unsigned(709, 10), 358 => to_unsigned(880, 10), 359 => to_unsigned(810, 10), 360 => to_unsigned(829, 10), 361 => to_unsigned(467, 10), 362 => to_unsigned(496, 10), 363 => to_unsigned(288, 10), 364 => to_unsigned(321, 10), 365 => to_unsigned(304, 10), 366 => to_unsigned(19, 10), 367 => to_unsigned(801, 10), 368 => to_unsigned(781, 10), 369 => to_unsigned(388, 10), 370 => to_unsigned(854, 10), 371 => to_unsigned(180, 10), 372 => to_unsigned(994, 10), 373 => to_unsigned(935, 10), 374 => to_unsigned(513, 10), 375 => to_unsigned(654, 10), 376 => to_unsigned(923, 10), 377 => to_unsigned(831, 10), 378 => to_unsigned(456, 10), 379 => to_unsigned(80, 10), 380 => to_unsigned(589, 10), 381 => to_unsigned(47, 10), 382 => to_unsigned(658, 10), 383 => to_unsigned(559, 10), 384 => to_unsigned(236, 10), 385 => to_unsigned(301, 10), 386 => to_unsigned(666, 10), 387 => to_unsigned(903, 10), 388 => to_unsigned(154, 10), 389 => to_unsigned(357, 10), 390 => to_unsigned(825, 10), 391 => to_unsigned(682, 10), 392 => to_unsigned(677, 10), 393 => to_unsigned(48, 10), 394 => to_unsigned(318, 10), 395 => to_unsigned(774, 10), 396 => to_unsigned(738, 10), 397 => to_unsigned(674, 10), 398 => to_unsigned(608, 10), 399 => to_unsigned(167, 10), 400 => to_unsigned(951, 10), 401 => to_unsigned(490, 10), 402 => to_unsigned(974, 10), 403 => to_unsigned(934, 10), 404 => to_unsigned(954, 10), 405 => to_unsigned(176, 10), 406 => to_unsigned(235, 10), 407 => to_unsigned(817, 10), 408 => to_unsigned(275, 10), 409 => to_unsigned(551, 10), 410 => to_unsigned(484, 10), 411 => to_unsigned(67, 10), 412 => to_unsigned(65, 10), 413 => to_unsigned(561, 10), 414 => to_unsigned(674, 10), 415 => to_unsigned(774, 10), 416 => to_unsigned(742, 10), 417 => to_unsigned(87, 10), 418 => to_unsigned(477, 10), 419 => to_unsigned(44, 10), 420 => to_unsigned(713, 10), 421 => to_unsigned(154, 10), 422 => to_unsigned(408, 10), 423 => to_unsigned(309, 10), 424 => to_unsigned(333, 10), 425 => to_unsigned(733, 10), 426 => to_unsigned(12, 10), 427 => to_unsigned(66, 10), 428 => to_unsigned(679, 10), 429 => to_unsigned(15, 10), 430 => to_unsigned(68, 10), 431 => to_unsigned(613, 10), 432 => to_unsigned(553, 10), 433 => to_unsigned(508, 10), 434 => to_unsigned(243, 10), 435 => to_unsigned(243, 10), 436 => to_unsigned(320, 10), 437 => to_unsigned(344, 10), 438 => to_unsigned(346, 10), 439 => to_unsigned(276, 10), 440 => to_unsigned(368, 10), 441 => to_unsigned(236, 10), 442 => to_unsigned(605, 10), 443 => to_unsigned(820, 10), 444 => to_unsigned(650, 10), 445 => to_unsigned(602, 10), 446 => to_unsigned(468, 10), 447 => to_unsigned(288, 10), 448 => to_unsigned(103, 10), 449 => to_unsigned(806, 10), 450 => to_unsigned(796, 10), 451 => to_unsigned(87, 10), 452 => to_unsigned(414, 10), 453 => to_unsigned(940, 10), 454 => to_unsigned(190, 10), 455 => to_unsigned(237, 10), 456 => to_unsigned(343, 10), 457 => to_unsigned(266, 10), 458 => to_unsigned(100, 10), 459 => to_unsigned(471, 10), 460 => to_unsigned(243, 10), 461 => to_unsigned(733, 10), 462 => to_unsigned(387, 10), 463 => to_unsigned(652, 10), 464 => to_unsigned(496, 10), 465 => to_unsigned(337, 10), 466 => to_unsigned(246, 10), 467 => to_unsigned(481, 10), 468 => to_unsigned(36, 10), 469 => to_unsigned(708, 10), 470 => to_unsigned(321, 10), 471 => to_unsigned(445, 10), 472 => to_unsigned(777, 10), 473 => to_unsigned(71, 10), 474 => to_unsigned(413, 10), 475 => to_unsigned(952, 10), 476 => to_unsigned(85, 10), 477 => to_unsigned(293, 10), 478 => to_unsigned(683, 10), 479 => to_unsigned(998, 10), 480 => to_unsigned(669, 10), 481 => to_unsigned(508, 10), 482 => to_unsigned(630, 10), 483 => to_unsigned(975, 10), 484 => to_unsigned(998, 10), 485 => to_unsigned(555, 10), 486 => to_unsigned(51, 10), 487 => to_unsigned(529, 10), 488 => to_unsigned(599, 10), 489 => to_unsigned(338, 10), 490 => to_unsigned(0, 10), 491 => to_unsigned(225, 10), 492 => to_unsigned(995, 10), 493 => to_unsigned(926, 10), 494 => to_unsigned(890, 10), 495 => to_unsigned(802, 10), 496 => to_unsigned(298, 10), 497 => to_unsigned(565, 10), 498 => to_unsigned(443, 10), 499 => to_unsigned(710, 10), 500 => to_unsigned(537, 10), 501 => to_unsigned(805, 10), 502 => to_unsigned(949, 10), 503 => to_unsigned(292, 10), 504 => to_unsigned(723, 10), 505 => to_unsigned(578, 10), 506 => to_unsigned(711, 10), 507 => to_unsigned(906, 10), 508 => to_unsigned(146, 10), 509 => to_unsigned(636, 10), 510 => to_unsigned(151, 10), 511 => to_unsigned(55, 10), 512 => to_unsigned(812, 10), 513 => to_unsigned(917, 10), 514 => to_unsigned(251, 10), 515 => to_unsigned(76, 10), 516 => to_unsigned(411, 10), 517 => to_unsigned(38, 10), 518 => to_unsigned(403, 10), 519 => to_unsigned(869, 10), 520 => to_unsigned(317, 10), 521 => to_unsigned(623, 10), 522 => to_unsigned(529, 10), 523 => to_unsigned(288, 10), 524 => to_unsigned(635, 10), 525 => to_unsigned(37, 10), 526 => to_unsigned(709, 10), 527 => to_unsigned(684, 10), 528 => to_unsigned(852, 10), 529 => to_unsigned(840, 10), 530 => to_unsigned(243, 10), 531 => to_unsigned(1, 10), 532 => to_unsigned(800, 10), 533 => to_unsigned(414, 10), 534 => to_unsigned(577, 10), 535 => to_unsigned(419, 10), 536 => to_unsigned(121, 10), 537 => to_unsigned(972, 10), 538 => to_unsigned(161, 10), 539 => to_unsigned(37, 10), 540 => to_unsigned(907, 10), 541 => to_unsigned(733, 10), 542 => to_unsigned(92, 10), 543 => to_unsigned(803, 10), 544 => to_unsigned(846, 10), 545 => to_unsigned(991, 10), 546 => to_unsigned(881, 10), 547 => to_unsigned(944, 10), 548 => to_unsigned(1004, 10), 549 => to_unsigned(98, 10), 550 => to_unsigned(639, 10), 551 => to_unsigned(523, 10), 552 => to_unsigned(134, 10), 553 => to_unsigned(322, 10), 554 => to_unsigned(726, 10), 555 => to_unsigned(158, 10), 556 => to_unsigned(216, 10), 557 => to_unsigned(622, 10), 558 => to_unsigned(656, 10), 559 => to_unsigned(82, 10), 560 => to_unsigned(654, 10), 561 => to_unsigned(291, 10), 562 => to_unsigned(994, 10), 563 => to_unsigned(130, 10), 564 => to_unsigned(387, 10), 565 => to_unsigned(558, 10), 566 => to_unsigned(967, 10), 567 => to_unsigned(257, 10), 568 => to_unsigned(83, 10), 569 => to_unsigned(67, 10), 570 => to_unsigned(343, 10), 571 => to_unsigned(3, 10), 572 => to_unsigned(730, 10), 573 => to_unsigned(355, 10), 574 => to_unsigned(74, 10), 575 => to_unsigned(579, 10), 576 => to_unsigned(534, 10), 577 => to_unsigned(918, 10), 578 => to_unsigned(193, 10), 579 => to_unsigned(397, 10), 580 => to_unsigned(446, 10), 581 => to_unsigned(80, 10), 582 => to_unsigned(141, 10), 583 => to_unsigned(784, 10), 584 => to_unsigned(162, 10), 585 => to_unsigned(796, 10), 586 => to_unsigned(601, 10), 587 => to_unsigned(17, 10), 588 => to_unsigned(723, 10), 589 => to_unsigned(558, 10), 590 => to_unsigned(444, 10), 591 => to_unsigned(781, 10), 592 => to_unsigned(77, 10), 593 => to_unsigned(416, 10), 594 => to_unsigned(498, 10), 595 => to_unsigned(390, 10), 596 => to_unsigned(187, 10), 597 => to_unsigned(787, 10), 598 => to_unsigned(662, 10), 599 => to_unsigned(692, 10), 600 => to_unsigned(515, 10), 601 => to_unsigned(680, 10), 602 => to_unsigned(279, 10), 603 => to_unsigned(892, 10), 604 => to_unsigned(352, 10), 605 => to_unsigned(974, 10), 606 => to_unsigned(131, 10), 607 => to_unsigned(938, 10), 608 => to_unsigned(914, 10), 609 => to_unsigned(867, 10), 610 => to_unsigned(908, 10), 611 => to_unsigned(849, 10), 612 => to_unsigned(363, 10), 613 => to_unsigned(966, 10), 614 => to_unsigned(238, 10), 615 => to_unsigned(206, 10), 616 => to_unsigned(385, 10), 617 => to_unsigned(158, 10), 618 => to_unsigned(327, 10), 619 => to_unsigned(504, 10), 620 => to_unsigned(473, 10), 621 => to_unsigned(189, 10), 622 => to_unsigned(98, 10), 623 => to_unsigned(608, 10), 624 => to_unsigned(16, 10), 625 => to_unsigned(633, 10), 626 => to_unsigned(899, 10), 627 => to_unsigned(178, 10), 628 => to_unsigned(389, 10), 629 => to_unsigned(820, 10), 630 => to_unsigned(422, 10), 631 => to_unsigned(53, 10), 632 => to_unsigned(111, 10), 633 => to_unsigned(427, 10), 634 => to_unsigned(216, 10), 635 => to_unsigned(614, 10), 636 => to_unsigned(367, 10), 637 => to_unsigned(597, 10), 638 => to_unsigned(612, 10), 639 => to_unsigned(1001, 10), 640 => to_unsigned(855, 10), 641 => to_unsigned(946, 10), 642 => to_unsigned(254, 10), 643 => to_unsigned(592, 10), 644 => to_unsigned(832, 10), 645 => to_unsigned(904, 10), 646 => to_unsigned(658, 10), 647 => to_unsigned(996, 10), 648 => to_unsigned(564, 10), 649 => to_unsigned(420, 10), 650 => to_unsigned(934, 10), 651 => to_unsigned(725, 10), 652 => to_unsigned(668, 10), 653 => to_unsigned(144, 10), 654 => to_unsigned(156, 10), 655 => to_unsigned(903, 10), 656 => to_unsigned(127, 10), 657 => to_unsigned(863, 10), 658 => to_unsigned(190, 10), 659 => to_unsigned(89, 10), 660 => to_unsigned(5, 10), 661 => to_unsigned(942, 10), 662 => to_unsigned(54, 10), 663 => to_unsigned(910, 10), 664 => to_unsigned(474, 10), 665 => to_unsigned(46, 10), 666 => to_unsigned(135, 10), 667 => to_unsigned(980, 10), 668 => to_unsigned(465, 10), 669 => to_unsigned(780, 10), 670 => to_unsigned(764, 10), 671 => to_unsigned(782, 10), 672 => to_unsigned(549, 10), 673 => to_unsigned(557, 10), 674 => to_unsigned(394, 10), 675 => to_unsigned(741, 10), 676 => to_unsigned(890, 10), 677 => to_unsigned(304, 10), 678 => to_unsigned(278, 10), 679 => to_unsigned(301, 10), 680 => to_unsigned(361, 10), 681 => to_unsigned(1001, 10), 682 => to_unsigned(290, 10), 683 => to_unsigned(804, 10), 684 => to_unsigned(491, 10), 685 => to_unsigned(375, 10), 686 => to_unsigned(767, 10), 687 => to_unsigned(982, 10), 688 => to_unsigned(725, 10), 689 => to_unsigned(625, 10), 690 => to_unsigned(362, 10), 691 => to_unsigned(844, 10), 692 => to_unsigned(452, 10), 693 => to_unsigned(940, 10), 694 => to_unsigned(629, 10), 695 => to_unsigned(390, 10), 696 => to_unsigned(799, 10), 697 => to_unsigned(504, 10), 698 => to_unsigned(290, 10), 699 => to_unsigned(419, 10), 700 => to_unsigned(381, 10), 701 => to_unsigned(0, 10), 702 => to_unsigned(898, 10), 703 => to_unsigned(870, 10), 704 => to_unsigned(362, 10), 705 => to_unsigned(719, 10), 706 => to_unsigned(922, 10), 707 => to_unsigned(905, 10), 708 => to_unsigned(963, 10), 709 => to_unsigned(627, 10), 710 => to_unsigned(901, 10), 711 => to_unsigned(355, 10), 712 => to_unsigned(554, 10), 713 => to_unsigned(246, 10), 714 => to_unsigned(564, 10), 715 => to_unsigned(535, 10), 716 => to_unsigned(435, 10), 717 => to_unsigned(920, 10), 718 => to_unsigned(638, 10), 719 => to_unsigned(806, 10), 720 => to_unsigned(973, 10), 721 => to_unsigned(1003, 10), 722 => to_unsigned(160, 10), 723 => to_unsigned(407, 10), 724 => to_unsigned(932, 10), 725 => to_unsigned(108, 10), 726 => to_unsigned(80, 10), 727 => to_unsigned(611, 10), 728 => to_unsigned(245, 10), 729 => to_unsigned(233, 10), 730 => to_unsigned(9, 10), 731 => to_unsigned(758, 10), 732 => to_unsigned(890, 10), 733 => to_unsigned(935, 10), 734 => to_unsigned(248, 10), 735 => to_unsigned(829, 10), 736 => to_unsigned(617, 10), 737 => to_unsigned(190, 10), 738 => to_unsigned(157, 10), 739 => to_unsigned(57, 10), 740 => to_unsigned(151, 10), 741 => to_unsigned(917, 10), 742 => to_unsigned(383, 10), 743 => to_unsigned(894, 10), 744 => to_unsigned(922, 10), 745 => to_unsigned(108, 10), 746 => to_unsigned(32, 10), 747 => to_unsigned(609, 10), 748 => to_unsigned(754, 10), 749 => to_unsigned(287, 10), 750 => to_unsigned(230, 10), 751 => to_unsigned(411, 10), 752 => to_unsigned(257, 10), 753 => to_unsigned(479, 10), 754 => to_unsigned(218, 10), 755 => to_unsigned(447, 10), 756 => to_unsigned(434, 10), 757 => to_unsigned(375, 10), 758 => to_unsigned(165, 10), 759 => to_unsigned(439, 10), 760 => to_unsigned(423, 10), 761 => to_unsigned(645, 10), 762 => to_unsigned(988, 10), 763 => to_unsigned(775, 10), 764 => to_unsigned(229, 10), 765 => to_unsigned(599, 10), 766 => to_unsigned(512, 10), 767 => to_unsigned(424, 10), 768 => to_unsigned(388, 10), 769 => to_unsigned(424, 10), 770 => to_unsigned(57, 10), 771 => to_unsigned(291, 10), 772 => to_unsigned(573, 10), 773 => to_unsigned(685, 10), 774 => to_unsigned(572, 10), 775 => to_unsigned(559, 10), 776 => to_unsigned(589, 10), 777 => to_unsigned(443, 10), 778 => to_unsigned(261, 10), 779 => to_unsigned(818, 10), 780 => to_unsigned(200, 10), 781 => to_unsigned(629, 10), 782 => to_unsigned(876, 10), 783 => to_unsigned(414, 10), 784 => to_unsigned(940, 10), 785 => to_unsigned(300, 10), 786 => to_unsigned(749, 10), 787 => to_unsigned(176, 10), 788 => to_unsigned(342, 10), 789 => to_unsigned(372, 10), 790 => to_unsigned(976, 10), 791 => to_unsigned(377, 10), 792 => to_unsigned(974, 10), 793 => to_unsigned(517, 10), 794 => to_unsigned(10, 10), 795 => to_unsigned(867, 10), 796 => to_unsigned(852, 10), 797 => to_unsigned(924, 10), 798 => to_unsigned(390, 10), 799 => to_unsigned(948, 10), 800 => to_unsigned(828, 10), 801 => to_unsigned(500, 10), 802 => to_unsigned(291, 10), 803 => to_unsigned(84, 10), 804 => to_unsigned(605, 10), 805 => to_unsigned(340, 10), 806 => to_unsigned(999, 10), 807 => to_unsigned(27, 10), 808 => to_unsigned(215, 10), 809 => to_unsigned(110, 10), 810 => to_unsigned(336, 10), 811 => to_unsigned(542, 10), 812 => to_unsigned(354, 10), 813 => to_unsigned(472, 10), 814 => to_unsigned(556, 10), 815 => to_unsigned(190, 10), 816 => to_unsigned(100, 10), 817 => to_unsigned(174, 10), 818 => to_unsigned(965, 10), 819 => to_unsigned(267, 10), 820 => to_unsigned(449, 10), 821 => to_unsigned(763, 10), 822 => to_unsigned(26, 10), 823 => to_unsigned(510, 10), 824 => to_unsigned(51, 10), 825 => to_unsigned(116, 10), 826 => to_unsigned(364, 10), 827 => to_unsigned(275, 10), 828 => to_unsigned(856, 10), 829 => to_unsigned(931, 10), 830 => to_unsigned(436, 10), 831 => to_unsigned(588, 10), 832 => to_unsigned(351, 10), 833 => to_unsigned(433, 10), 834 => to_unsigned(450, 10), 835 => to_unsigned(28, 10), 836 => to_unsigned(500, 10), 837 => to_unsigned(24, 10), 838 => to_unsigned(553, 10), 839 => to_unsigned(168, 10), 840 => to_unsigned(401, 10), 841 => to_unsigned(150, 10), 842 => to_unsigned(876, 10), 843 => to_unsigned(582, 10), 844 => to_unsigned(501, 10), 845 => to_unsigned(762, 10), 846 => to_unsigned(339, 10), 847 => to_unsigned(717, 10), 848 => to_unsigned(257, 10), 849 => to_unsigned(803, 10), 850 => to_unsigned(219, 10), 851 => to_unsigned(67, 10), 852 => to_unsigned(1008, 10), 853 => to_unsigned(443, 10), 854 => to_unsigned(522, 10), 855 => to_unsigned(788, 10), 856 => to_unsigned(743, 10), 857 => to_unsigned(0, 10), 858 => to_unsigned(145, 10), 859 => to_unsigned(191, 10), 860 => to_unsigned(137, 10), 861 => to_unsigned(731, 10), 862 => to_unsigned(172, 10), 863 => to_unsigned(96, 10), 864 => to_unsigned(240, 10), 865 => to_unsigned(525, 10), 866 => to_unsigned(322, 10), 867 => to_unsigned(239, 10), 868 => to_unsigned(365, 10), 869 => to_unsigned(172, 10), 870 => to_unsigned(134, 10), 871 => to_unsigned(281, 10), 872 => to_unsigned(35, 10), 873 => to_unsigned(759, 10), 874 => to_unsigned(649, 10), 875 => to_unsigned(800, 10), 876 => to_unsigned(79, 10), 877 => to_unsigned(249, 10), 878 => to_unsigned(618, 10), 879 => to_unsigned(822, 10), 880 => to_unsigned(921, 10), 881 => to_unsigned(203, 10), 882 => to_unsigned(292, 10), 883 => to_unsigned(192, 10), 884 => to_unsigned(223, 10), 885 => to_unsigned(761, 10), 886 => to_unsigned(237, 10), 887 => to_unsigned(621, 10), 888 => to_unsigned(759, 10), 889 => to_unsigned(739, 10), 890 => to_unsigned(958, 10), 891 => to_unsigned(657, 10), 892 => to_unsigned(330, 10), 893 => to_unsigned(422, 10), 894 => to_unsigned(714, 10), 895 => to_unsigned(246, 10), 896 => to_unsigned(263, 10), 897 => to_unsigned(573, 10), 898 => to_unsigned(874, 10), 899 => to_unsigned(298, 10), 900 => to_unsigned(383, 10), 901 => to_unsigned(742, 10), 902 => to_unsigned(26, 10), 903 => to_unsigned(513, 10), 904 => to_unsigned(657, 10), 905 => to_unsigned(369, 10), 906 => to_unsigned(460, 10), 907 => to_unsigned(90, 10), 908 => to_unsigned(254, 10), 909 => to_unsigned(479, 10), 910 => to_unsigned(380, 10), 911 => to_unsigned(811, 10), 912 => to_unsigned(606, 10), 913 => to_unsigned(798, 10), 914 => to_unsigned(502, 10), 915 => to_unsigned(889, 10), 916 => to_unsigned(205, 10), 917 => to_unsigned(920, 10), 918 => to_unsigned(988, 10), 919 => to_unsigned(710, 10), 920 => to_unsigned(63, 10), 921 => to_unsigned(212, 10), 922 => to_unsigned(1001, 10), 923 => to_unsigned(996, 10), 924 => to_unsigned(266, 10), 925 => to_unsigned(231, 10), 926 => to_unsigned(643, 10), 927 => to_unsigned(964, 10), 928 => to_unsigned(342, 10), 929 => to_unsigned(539, 10), 930 => to_unsigned(592, 10), 931 => to_unsigned(540, 10), 932 => to_unsigned(487, 10), 933 => to_unsigned(998, 10), 934 => to_unsigned(850, 10), 935 => to_unsigned(563, 10), 936 => to_unsigned(652, 10), 937 => to_unsigned(216, 10), 938 => to_unsigned(638, 10), 939 => to_unsigned(933, 10), 940 => to_unsigned(391, 10), 941 => to_unsigned(51, 10), 942 => to_unsigned(76, 10), 943 => to_unsigned(833, 10), 944 => to_unsigned(73, 10), 945 => to_unsigned(561, 10), 946 => to_unsigned(283, 10), 947 => to_unsigned(236, 10), 948 => to_unsigned(99, 10), 949 => to_unsigned(104, 10), 950 => to_unsigned(72, 10), 951 => to_unsigned(690, 10), 952 => to_unsigned(433, 10), 953 => to_unsigned(967, 10), 954 => to_unsigned(195, 10), 955 => to_unsigned(122, 10), 956 => to_unsigned(970, 10), 957 => to_unsigned(470, 10), 958 => to_unsigned(997, 10), 959 => to_unsigned(751, 10), 960 => to_unsigned(654, 10), 961 => to_unsigned(867, 10), 962 => to_unsigned(978, 10), 963 => to_unsigned(51, 10), 964 => to_unsigned(501, 10), 965 => to_unsigned(717, 10), 966 => to_unsigned(386, 10), 967 => to_unsigned(338, 10), 968 => to_unsigned(838, 10), 969 => to_unsigned(488, 10), 970 => to_unsigned(903, 10), 971 => to_unsigned(854, 10), 972 => to_unsigned(808, 10), 973 => to_unsigned(655, 10), 974 => to_unsigned(1003, 10), 975 => to_unsigned(539, 10), 976 => to_unsigned(757, 10), 977 => to_unsigned(1001, 10), 978 => to_unsigned(902, 10), 979 => to_unsigned(760, 10), 980 => to_unsigned(488, 10), 981 => to_unsigned(707, 10), 982 => to_unsigned(508, 10), 983 => to_unsigned(101, 10), 984 => to_unsigned(846, 10), 985 => to_unsigned(93, 10), 986 => to_unsigned(288, 10), 987 => to_unsigned(791, 10), 988 => to_unsigned(528, 10), 989 => to_unsigned(304, 10), 990 => to_unsigned(857, 10), 991 => to_unsigned(453, 10), 992 => to_unsigned(680, 10), 993 => to_unsigned(167, 10), 994 => to_unsigned(382, 10), 995 => to_unsigned(802, 10), 996 => to_unsigned(845, 10), 997 => to_unsigned(295, 10), 998 => to_unsigned(467, 10), 999 => to_unsigned(855, 10), 1000 => to_unsigned(45, 10), 1001 => to_unsigned(506, 10), 1002 => to_unsigned(564, 10), 1003 => to_unsigned(399, 10), 1004 => to_unsigned(196, 10), 1005 => to_unsigned(159, 10), 1006 => to_unsigned(891, 10), 1007 => to_unsigned(578, 10), 1008 => to_unsigned(34, 10), 1009 => to_unsigned(520, 10), 1010 => to_unsigned(214, 10), 1011 => to_unsigned(942, 10), 1012 => to_unsigned(993, 10), 1013 => to_unsigned(879, 10), 1014 => to_unsigned(755, 10), 1015 => to_unsigned(328, 10), 1016 => to_unsigned(241, 10), 1017 => to_unsigned(181, 10), 1018 => to_unsigned(595, 10), 1019 => to_unsigned(377, 10), 1020 => to_unsigned(925, 10), 1021 => to_unsigned(255, 10), 1022 => to_unsigned(264, 10), 1023 => to_unsigned(910, 10), 1024 => to_unsigned(485, 10), 1025 => to_unsigned(213, 10), 1026 => to_unsigned(918, 10), 1027 => to_unsigned(483, 10), 1028 => to_unsigned(484, 10), 1029 => to_unsigned(470, 10), 1030 => to_unsigned(197, 10), 1031 => to_unsigned(557, 10), 1032 => to_unsigned(538, 10), 1033 => to_unsigned(675, 10), 1034 => to_unsigned(235, 10), 1035 => to_unsigned(32, 10), 1036 => to_unsigned(84, 10), 1037 => to_unsigned(583, 10), 1038 => to_unsigned(985, 10), 1039 => to_unsigned(325, 10), 1040 => to_unsigned(559, 10), 1041 => to_unsigned(502, 10), 1042 => to_unsigned(729, 10), 1043 => to_unsigned(500, 10), 1044 => to_unsigned(652, 10), 1045 => to_unsigned(553, 10), 1046 => to_unsigned(520, 10), 1047 => to_unsigned(496, 10), 1048 => to_unsigned(72, 10), 1049 => to_unsigned(346, 10), 1050 => to_unsigned(46, 10), 1051 => to_unsigned(734, 10), 1052 => to_unsigned(278, 10), 1053 => to_unsigned(982, 10), 1054 => to_unsigned(513, 10), 1055 => to_unsigned(628, 10), 1056 => to_unsigned(1012, 10), 1057 => to_unsigned(714, 10), 1058 => to_unsigned(178, 10), 1059 => to_unsigned(840, 10), 1060 => to_unsigned(497, 10), 1061 => to_unsigned(971, 10), 1062 => to_unsigned(597, 10), 1063 => to_unsigned(259, 10), 1064 => to_unsigned(488, 10), 1065 => to_unsigned(573, 10), 1066 => to_unsigned(683, 10), 1067 => to_unsigned(803, 10), 1068 => to_unsigned(352, 10), 1069 => to_unsigned(231, 10), 1070 => to_unsigned(387, 10), 1071 => to_unsigned(747, 10), 1072 => to_unsigned(655, 10), 1073 => to_unsigned(617, 10), 1074 => to_unsigned(260, 10), 1075 => to_unsigned(389, 10), 1076 => to_unsigned(814, 10), 1077 => to_unsigned(13, 10), 1078 => to_unsigned(217, 10), 1079 => to_unsigned(634, 10), 1080 => to_unsigned(978, 10), 1081 => to_unsigned(551, 10), 1082 => to_unsigned(197, 10), 1083 => to_unsigned(526, 10), 1084 => to_unsigned(715, 10), 1085 => to_unsigned(826, 10), 1086 => to_unsigned(940, 10), 1087 => to_unsigned(586, 10), 1088 => to_unsigned(555, 10), 1089 => to_unsigned(335, 10), 1090 => to_unsigned(655, 10), 1091 => to_unsigned(23, 10), 1092 => to_unsigned(228, 10), 1093 => to_unsigned(447, 10), 1094 => to_unsigned(528, 10), 1095 => to_unsigned(62, 10), 1096 => to_unsigned(849, 10), 1097 => to_unsigned(424, 10), 1098 => to_unsigned(865, 10), 1099 => to_unsigned(949, 10), 1100 => to_unsigned(761, 10), 1101 => to_unsigned(176, 10), 1102 => to_unsigned(506, 10), 1103 => to_unsigned(621, 10), 1104 => to_unsigned(623, 10), 1105 => to_unsigned(180, 10), 1106 => to_unsigned(15, 10), 1107 => to_unsigned(894, 10), 1108 => to_unsigned(23, 10), 1109 => to_unsigned(974, 10), 1110 => to_unsigned(305, 10), 1111 => to_unsigned(520, 10), 1112 => to_unsigned(288, 10), 1113 => to_unsigned(929, 10), 1114 => to_unsigned(379, 10), 1115 => to_unsigned(657, 10), 1116 => to_unsigned(899, 10), 1117 => to_unsigned(405, 10), 1118 => to_unsigned(56, 10), 1119 => to_unsigned(75, 10), 1120 => to_unsigned(988, 10), 1121 => to_unsigned(502, 10), 1122 => to_unsigned(1000, 10), 1123 => to_unsigned(672, 10), 1124 => to_unsigned(281, 10), 1125 => to_unsigned(858, 10), 1126 => to_unsigned(989, 10), 1127 => to_unsigned(308, 10), 1128 => to_unsigned(774, 10), 1129 => to_unsigned(223, 10), 1130 => to_unsigned(847, 10), 1131 => to_unsigned(521, 10), 1132 => to_unsigned(857, 10), 1133 => to_unsigned(737, 10), 1134 => to_unsigned(847, 10), 1135 => to_unsigned(219, 10), 1136 => to_unsigned(747, 10), 1137 => to_unsigned(246, 10), 1138 => to_unsigned(670, 10), 1139 => to_unsigned(760, 10), 1140 => to_unsigned(894, 10), 1141 => to_unsigned(738, 10), 1142 => to_unsigned(872, 10), 1143 => to_unsigned(883, 10), 1144 => to_unsigned(706, 10), 1145 => to_unsigned(270, 10), 1146 => to_unsigned(480, 10), 1147 => to_unsigned(107, 10), 1148 => to_unsigned(912, 10), 1149 => to_unsigned(399, 10), 1150 => to_unsigned(207, 10), 1151 => to_unsigned(430, 10), 1152 => to_unsigned(526, 10), 1153 => to_unsigned(126, 10), 1154 => to_unsigned(487, 10), 1155 => to_unsigned(989, 10), 1156 => to_unsigned(436, 10), 1157 => to_unsigned(405, 10), 1158 => to_unsigned(359, 10), 1159 => to_unsigned(25, 10), 1160 => to_unsigned(588, 10), 1161 => to_unsigned(459, 10), 1162 => to_unsigned(545, 10), 1163 => to_unsigned(576, 10), 1164 => to_unsigned(231, 10), 1165 => to_unsigned(430, 10), 1166 => to_unsigned(299, 10), 1167 => to_unsigned(611, 10), 1168 => to_unsigned(20, 10), 1169 => to_unsigned(40, 10), 1170 => to_unsigned(540, 10), 1171 => to_unsigned(661, 10), 1172 => to_unsigned(14, 10), 1173 => to_unsigned(850, 10), 1174 => to_unsigned(795, 10), 1175 => to_unsigned(394, 10), 1176 => to_unsigned(144, 10), 1177 => to_unsigned(1003, 10), 1178 => to_unsigned(268, 10), 1179 => to_unsigned(687, 10), 1180 => to_unsigned(180, 10), 1181 => to_unsigned(556, 10), 1182 => to_unsigned(433, 10), 1183 => to_unsigned(790, 10), 1184 => to_unsigned(627, 10), 1185 => to_unsigned(320, 10), 1186 => to_unsigned(778, 10), 1187 => to_unsigned(921, 10), 1188 => to_unsigned(139, 10), 1189 => to_unsigned(383, 10), 1190 => to_unsigned(975, 10), 1191 => to_unsigned(671, 10), 1192 => to_unsigned(195, 10), 1193 => to_unsigned(994, 10), 1194 => to_unsigned(998, 10), 1195 => to_unsigned(334, 10), 1196 => to_unsigned(1009, 10), 1197 => to_unsigned(862, 10), 1198 => to_unsigned(836, 10), 1199 => to_unsigned(936, 10), 1200 => to_unsigned(281, 10), 1201 => to_unsigned(415, 10), 1202 => to_unsigned(934, 10), 1203 => to_unsigned(134, 10), 1204 => to_unsigned(793, 10), 1205 => to_unsigned(555, 10), 1206 => to_unsigned(787, 10), 1207 => to_unsigned(290, 10), 1208 => to_unsigned(55, 10), 1209 => to_unsigned(277, 10), 1210 => to_unsigned(487, 10), 1211 => to_unsigned(78, 10), 1212 => to_unsigned(751, 10), 1213 => to_unsigned(310, 10), 1214 => to_unsigned(273, 10), 1215 => to_unsigned(756, 10), 1216 => to_unsigned(793, 10), 1217 => to_unsigned(670, 10), 1218 => to_unsigned(793, 10), 1219 => to_unsigned(1007, 10), 1220 => to_unsigned(693, 10), 1221 => to_unsigned(245, 10), 1222 => to_unsigned(191, 10), 1223 => to_unsigned(346, 10), 1224 => to_unsigned(888, 10), 1225 => to_unsigned(518, 10), 1226 => to_unsigned(1, 10), 1227 => to_unsigned(362, 10), 1228 => to_unsigned(612, 10), 1229 => to_unsigned(453, 10), 1230 => to_unsigned(375, 10), 1231 => to_unsigned(429, 10), 1232 => to_unsigned(51, 10), 1233 => to_unsigned(598, 10), 1234 => to_unsigned(322, 10), 1235 => to_unsigned(17, 10), 1236 => to_unsigned(438, 10), 1237 => to_unsigned(409, 10), 1238 => to_unsigned(206, 10), 1239 => to_unsigned(942, 10), 1240 => to_unsigned(123, 10), 1241 => to_unsigned(307, 10), 1242 => to_unsigned(95, 10), 1243 => to_unsigned(483, 10), 1244 => to_unsigned(496, 10), 1245 => to_unsigned(1012, 10), 1246 => to_unsigned(558, 10), 1247 => to_unsigned(928, 10), 1248 => to_unsigned(355, 10), 1249 => to_unsigned(580, 10), 1250 => to_unsigned(457, 10), 1251 => to_unsigned(591, 10), 1252 => to_unsigned(862, 10), 1253 => to_unsigned(862, 10), 1254 => to_unsigned(1011, 10), 1255 => to_unsigned(927, 10), 1256 => to_unsigned(430, 10), 1257 => to_unsigned(197, 10), 1258 => to_unsigned(877, 10), 1259 => to_unsigned(808, 10), 1260 => to_unsigned(839, 10), 1261 => to_unsigned(222, 10), 1262 => to_unsigned(67, 10), 1263 => to_unsigned(336, 10), 1264 => to_unsigned(155, 10), 1265 => to_unsigned(552, 10), 1266 => to_unsigned(97, 10), 1267 => to_unsigned(253, 10), 1268 => to_unsigned(753, 10), 1269 => to_unsigned(883, 10), 1270 => to_unsigned(550, 10), 1271 => to_unsigned(143, 10), 1272 => to_unsigned(545, 10), 1273 => to_unsigned(461, 10), 1274 => to_unsigned(165, 10), 1275 => to_unsigned(819, 10), 1276 => to_unsigned(711, 10), 1277 => to_unsigned(945, 10), 1278 => to_unsigned(600, 10), 1279 => to_unsigned(132, 10), 1280 => to_unsigned(192, 10), 1281 => to_unsigned(844, 10), 1282 => to_unsigned(247, 10), 1283 => to_unsigned(651, 10), 1284 => to_unsigned(1007, 10), 1285 => to_unsigned(392, 10), 1286 => to_unsigned(351, 10), 1287 => to_unsigned(363, 10), 1288 => to_unsigned(879, 10), 1289 => to_unsigned(359, 10), 1290 => to_unsigned(608, 10), 1291 => to_unsigned(552, 10), 1292 => to_unsigned(37, 10), 1293 => to_unsigned(1003, 10), 1294 => to_unsigned(252, 10), 1295 => to_unsigned(613, 10), 1296 => to_unsigned(397, 10), 1297 => to_unsigned(15, 10), 1298 => to_unsigned(249, 10), 1299 => to_unsigned(238, 10), 1300 => to_unsigned(627, 10), 1301 => to_unsigned(442, 10), 1302 => to_unsigned(347, 10), 1303 => to_unsigned(246, 10), 1304 => to_unsigned(39, 10), 1305 => to_unsigned(785, 10), 1306 => to_unsigned(598, 10), 1307 => to_unsigned(754, 10), 1308 => to_unsigned(139, 10), 1309 => to_unsigned(367, 10), 1310 => to_unsigned(474, 10), 1311 => to_unsigned(955, 10), 1312 => to_unsigned(19, 10), 1313 => to_unsigned(428, 10), 1314 => to_unsigned(19, 10), 1315 => to_unsigned(437, 10), 1316 => to_unsigned(460, 10), 1317 => to_unsigned(118, 10), 1318 => to_unsigned(851, 10), 1319 => to_unsigned(103, 10), 1320 => to_unsigned(886, 10), 1321 => to_unsigned(169, 10), 1322 => to_unsigned(50, 10), 1323 => to_unsigned(876, 10), 1324 => to_unsigned(50, 10), 1325 => to_unsigned(676, 10), 1326 => to_unsigned(939, 10), 1327 => to_unsigned(994, 10), 1328 => to_unsigned(170, 10), 1329 => to_unsigned(105, 10), 1330 => to_unsigned(948, 10), 1331 => to_unsigned(130, 10), 1332 => to_unsigned(253, 10), 1333 => to_unsigned(516, 10), 1334 => to_unsigned(791, 10), 1335 => to_unsigned(549, 10), 1336 => to_unsigned(878, 10), 1337 => to_unsigned(887, 10), 1338 => to_unsigned(205, 10), 1339 => to_unsigned(118, 10), 1340 => to_unsigned(669, 10), 1341 => to_unsigned(659, 10), 1342 => to_unsigned(37, 10), 1343 => to_unsigned(606, 10), 1344 => to_unsigned(430, 10), 1345 => to_unsigned(39, 10), 1346 => to_unsigned(496, 10), 1347 => to_unsigned(534, 10), 1348 => to_unsigned(570, 10), 1349 => to_unsigned(96, 10), 1350 => to_unsigned(272, 10), 1351 => to_unsigned(86, 10), 1352 => to_unsigned(470, 10), 1353 => to_unsigned(361, 10), 1354 => to_unsigned(395, 10), 1355 => to_unsigned(435, 10), 1356 => to_unsigned(304, 10), 1357 => to_unsigned(755, 10), 1358 => to_unsigned(806, 10), 1359 => to_unsigned(920, 10), 1360 => to_unsigned(746, 10), 1361 => to_unsigned(492, 10), 1362 => to_unsigned(11, 10), 1363 => to_unsigned(888, 10), 1364 => to_unsigned(816, 10), 1365 => to_unsigned(511, 10), 1366 => to_unsigned(436, 10), 1367 => to_unsigned(510, 10), 1368 => to_unsigned(371, 10), 1369 => to_unsigned(300, 10), 1370 => to_unsigned(549, 10), 1371 => to_unsigned(976, 10), 1372 => to_unsigned(792, 10), 1373 => to_unsigned(1010, 10), 1374 => to_unsigned(704, 10), 1375 => to_unsigned(646, 10), 1376 => to_unsigned(718, 10), 1377 => to_unsigned(998, 10), 1378 => to_unsigned(1001, 10), 1379 => to_unsigned(172, 10), 1380 => to_unsigned(476, 10), 1381 => to_unsigned(553, 10), 1382 => to_unsigned(88, 10), 1383 => to_unsigned(185, 10), 1384 => to_unsigned(866, 10), 1385 => to_unsigned(52, 10), 1386 => to_unsigned(719, 10), 1387 => to_unsigned(412, 10), 1388 => to_unsigned(134, 10), 1389 => to_unsigned(792, 10), 1390 => to_unsigned(790, 10), 1391 => to_unsigned(386, 10), 1392 => to_unsigned(392, 10), 1393 => to_unsigned(683, 10), 1394 => to_unsigned(164, 10), 1395 => to_unsigned(236, 10), 1396 => to_unsigned(692, 10), 1397 => to_unsigned(391, 10), 1398 => to_unsigned(868, 10), 1399 => to_unsigned(303, 10), 1400 => to_unsigned(195, 10), 1401 => to_unsigned(34, 10), 1402 => to_unsigned(584, 10), 1403 => to_unsigned(708, 10), 1404 => to_unsigned(244, 10), 1405 => to_unsigned(664, 10), 1406 => to_unsigned(69, 10), 1407 => to_unsigned(717, 10), 1408 => to_unsigned(805, 10), 1409 => to_unsigned(36, 10), 1410 => to_unsigned(374, 10), 1411 => to_unsigned(890, 10), 1412 => to_unsigned(585, 10), 1413 => to_unsigned(710, 10), 1414 => to_unsigned(117, 10), 1415 => to_unsigned(851, 10), 1416 => to_unsigned(566, 10), 1417 => to_unsigned(804, 10), 1418 => to_unsigned(864, 10), 1419 => to_unsigned(186, 10), 1420 => to_unsigned(414, 10), 1421 => to_unsigned(238, 10), 1422 => to_unsigned(775, 10), 1423 => to_unsigned(455, 10), 1424 => to_unsigned(749, 10), 1425 => to_unsigned(242, 10), 1426 => to_unsigned(144, 10), 1427 => to_unsigned(136, 10), 1428 => to_unsigned(495, 10), 1429 => to_unsigned(837, 10), 1430 => to_unsigned(699, 10), 1431 => to_unsigned(885, 10), 1432 => to_unsigned(895, 10), 1433 => to_unsigned(695, 10), 1434 => to_unsigned(758, 10), 1435 => to_unsigned(340, 10), 1436 => to_unsigned(996, 10), 1437 => to_unsigned(654, 10), 1438 => to_unsigned(754, 10), 1439 => to_unsigned(643, 10), 1440 => to_unsigned(405, 10), 1441 => to_unsigned(391, 10), 1442 => to_unsigned(623, 10), 1443 => to_unsigned(688, 10), 1444 => to_unsigned(258, 10), 1445 => to_unsigned(745, 10), 1446 => to_unsigned(165, 10), 1447 => to_unsigned(244, 10), 1448 => to_unsigned(734, 10), 1449 => to_unsigned(533, 10), 1450 => to_unsigned(628, 10), 1451 => to_unsigned(195, 10), 1452 => to_unsigned(356, 10), 1453 => to_unsigned(591, 10), 1454 => to_unsigned(445, 10), 1455 => to_unsigned(923, 10), 1456 => to_unsigned(1006, 10), 1457 => to_unsigned(696, 10), 1458 => to_unsigned(263, 10), 1459 => to_unsigned(101, 10), 1460 => to_unsigned(695, 10), 1461 => to_unsigned(204, 10), 1462 => to_unsigned(294, 10), 1463 => to_unsigned(977, 10), 1464 => to_unsigned(772, 10), 1465 => to_unsigned(590, 10), 1466 => to_unsigned(302, 10), 1467 => to_unsigned(775, 10), 1468 => to_unsigned(201, 10), 1469 => to_unsigned(513, 10), 1470 => to_unsigned(276, 10), 1471 => to_unsigned(630, 10), 1472 => to_unsigned(388, 10), 1473 => to_unsigned(997, 10), 1474 => to_unsigned(320, 10), 1475 => to_unsigned(988, 10), 1476 => to_unsigned(94, 10), 1477 => to_unsigned(679, 10), 1478 => to_unsigned(670, 10), 1479 => to_unsigned(695, 10), 1480 => to_unsigned(940, 10), 1481 => to_unsigned(617, 10), 1482 => to_unsigned(562, 10), 1483 => to_unsigned(618, 10), 1484 => to_unsigned(228, 10), 1485 => to_unsigned(24, 10), 1486 => to_unsigned(341, 10), 1487 => to_unsigned(273, 10), 1488 => to_unsigned(71, 10), 1489 => to_unsigned(154, 10), 1490 => to_unsigned(162, 10), 1491 => to_unsigned(1019, 10), 1492 => to_unsigned(741, 10), 1493 => to_unsigned(360, 10), 1494 => to_unsigned(315, 10), 1495 => to_unsigned(999, 10), 1496 => to_unsigned(948, 10), 1497 => to_unsigned(707, 10), 1498 => to_unsigned(752, 10), 1499 => to_unsigned(23, 10), 1500 => to_unsigned(505, 10), 1501 => to_unsigned(73, 10), 1502 => to_unsigned(356, 10), 1503 => to_unsigned(238, 10), 1504 => to_unsigned(1005, 10), 1505 => to_unsigned(101, 10), 1506 => to_unsigned(734, 10), 1507 => to_unsigned(405, 10), 1508 => to_unsigned(419, 10), 1509 => to_unsigned(772, 10), 1510 => to_unsigned(83, 10), 1511 => to_unsigned(326, 10), 1512 => to_unsigned(54, 10), 1513 => to_unsigned(890, 10), 1514 => to_unsigned(792, 10), 1515 => to_unsigned(228, 10), 1516 => to_unsigned(457, 10), 1517 => to_unsigned(359, 10), 1518 => to_unsigned(613, 10), 1519 => to_unsigned(63, 10), 1520 => to_unsigned(776, 10), 1521 => to_unsigned(224, 10), 1522 => to_unsigned(627, 10), 1523 => to_unsigned(978, 10), 1524 => to_unsigned(215, 10), 1525 => to_unsigned(14, 10), 1526 => to_unsigned(905, 10), 1527 => to_unsigned(959, 10), 1528 => to_unsigned(168, 10), 1529 => to_unsigned(121, 10), 1530 => to_unsigned(877, 10), 1531 => to_unsigned(482, 10), 1532 => to_unsigned(771, 10), 1533 => to_unsigned(872, 10), 1534 => to_unsigned(4, 10), 1535 => to_unsigned(760, 10), 1536 => to_unsigned(592, 10), 1537 => to_unsigned(204, 10), 1538 => to_unsigned(900, 10), 1539 => to_unsigned(761, 10), 1540 => to_unsigned(95, 10), 1541 => to_unsigned(32, 10), 1542 => to_unsigned(207, 10), 1543 => to_unsigned(284, 10), 1544 => to_unsigned(213, 10), 1545 => to_unsigned(949, 10), 1546 => to_unsigned(372, 10), 1547 => to_unsigned(717, 10), 1548 => to_unsigned(552, 10), 1549 => to_unsigned(819, 10), 1550 => to_unsigned(1011, 10), 1551 => to_unsigned(220, 10), 1552 => to_unsigned(960, 10), 1553 => to_unsigned(713, 10), 1554 => to_unsigned(13, 10), 1555 => to_unsigned(602, 10), 1556 => to_unsigned(587, 10), 1557 => to_unsigned(428, 10), 1558 => to_unsigned(777, 10), 1559 => to_unsigned(634, 10), 1560 => to_unsigned(150, 10), 1561 => to_unsigned(281, 10), 1562 => to_unsigned(320, 10), 1563 => to_unsigned(438, 10), 1564 => to_unsigned(152, 10), 1565 => to_unsigned(708, 10), 1566 => to_unsigned(175, 10), 1567 => to_unsigned(1009, 10), 1568 => to_unsigned(617, 10), 1569 => to_unsigned(916, 10), 1570 => to_unsigned(140, 10), 1571 => to_unsigned(884, 10), 1572 => to_unsigned(276, 10), 1573 => to_unsigned(861, 10), 1574 => to_unsigned(202, 10), 1575 => to_unsigned(971, 10), 1576 => to_unsigned(981, 10), 1577 => to_unsigned(793, 10), 1578 => to_unsigned(606, 10), 1579 => to_unsigned(423, 10), 1580 => to_unsigned(280, 10), 1581 => to_unsigned(981, 10), 1582 => to_unsigned(329, 10), 1583 => to_unsigned(550, 10), 1584 => to_unsigned(36, 10), 1585 => to_unsigned(989, 10), 1586 => to_unsigned(1016, 10), 1587 => to_unsigned(657, 10), 1588 => to_unsigned(753, 10), 1589 => to_unsigned(959, 10), 1590 => to_unsigned(425, 10), 1591 => to_unsigned(486, 10), 1592 => to_unsigned(866, 10), 1593 => to_unsigned(326, 10), 1594 => to_unsigned(956, 10), 1595 => to_unsigned(972, 10), 1596 => to_unsigned(345, 10), 1597 => to_unsigned(206, 10), 1598 => to_unsigned(12, 10), 1599 => to_unsigned(275, 10), 1600 => to_unsigned(326, 10), 1601 => to_unsigned(565, 10), 1602 => to_unsigned(777, 10), 1603 => to_unsigned(885, 10), 1604 => to_unsigned(809, 10), 1605 => to_unsigned(479, 10), 1606 => to_unsigned(948, 10), 1607 => to_unsigned(467, 10), 1608 => to_unsigned(573, 10), 1609 => to_unsigned(115, 10), 1610 => to_unsigned(1003, 10), 1611 => to_unsigned(141, 10), 1612 => to_unsigned(36, 10), 1613 => to_unsigned(830, 10), 1614 => to_unsigned(662, 10), 1615 => to_unsigned(652, 10), 1616 => to_unsigned(579, 10), 1617 => to_unsigned(975, 10), 1618 => to_unsigned(747, 10), 1619 => to_unsigned(387, 10), 1620 => to_unsigned(443, 10), 1621 => to_unsigned(930, 10), 1622 => to_unsigned(102, 10), 1623 => to_unsigned(291, 10), 1624 => to_unsigned(902, 10), 1625 => to_unsigned(651, 10), 1626 => to_unsigned(829, 10), 1627 => to_unsigned(962, 10), 1628 => to_unsigned(347, 10), 1629 => to_unsigned(75, 10), 1630 => to_unsigned(954, 10), 1631 => to_unsigned(198, 10), 1632 => to_unsigned(568, 10), 1633 => to_unsigned(479, 10), 1634 => to_unsigned(846, 10), 1635 => to_unsigned(408, 10), 1636 => to_unsigned(28, 10), 1637 => to_unsigned(874, 10), 1638 => to_unsigned(937, 10), 1639 => to_unsigned(526, 10), 1640 => to_unsigned(292, 10), 1641 => to_unsigned(851, 10), 1642 => to_unsigned(689, 10), 1643 => to_unsigned(297, 10), 1644 => to_unsigned(914, 10), 1645 => to_unsigned(440, 10), 1646 => to_unsigned(567, 10), 1647 => to_unsigned(242, 10), 1648 => to_unsigned(494, 10), 1649 => to_unsigned(692, 10), 1650 => to_unsigned(747, 10), 1651 => to_unsigned(433, 10), 1652 => to_unsigned(794, 10), 1653 => to_unsigned(547, 10), 1654 => to_unsigned(881, 10), 1655 => to_unsigned(627, 10), 1656 => to_unsigned(629, 10), 1657 => to_unsigned(209, 10), 1658 => to_unsigned(1016, 10), 1659 => to_unsigned(902, 10), 1660 => to_unsigned(836, 10), 1661 => to_unsigned(756, 10), 1662 => to_unsigned(250, 10), 1663 => to_unsigned(570, 10), 1664 => to_unsigned(741, 10), 1665 => to_unsigned(721, 10), 1666 => to_unsigned(38, 10), 1667 => to_unsigned(542, 10), 1668 => to_unsigned(695, 10), 1669 => to_unsigned(675, 10), 1670 => to_unsigned(976, 10), 1671 => to_unsigned(472, 10), 1672 => to_unsigned(429, 10), 1673 => to_unsigned(5, 10), 1674 => to_unsigned(978, 10), 1675 => to_unsigned(994, 10), 1676 => to_unsigned(815, 10), 1677 => to_unsigned(622, 10), 1678 => to_unsigned(1005, 10), 1679 => to_unsigned(444, 10), 1680 => to_unsigned(599, 10), 1681 => to_unsigned(987, 10), 1682 => to_unsigned(704, 10), 1683 => to_unsigned(1012, 10), 1684 => to_unsigned(840, 10), 1685 => to_unsigned(549, 10), 1686 => to_unsigned(974, 10), 1687 => to_unsigned(28, 10), 1688 => to_unsigned(658, 10), 1689 => to_unsigned(838, 10), 1690 => to_unsigned(264, 10), 1691 => to_unsigned(612, 10), 1692 => to_unsigned(358, 10), 1693 => to_unsigned(66, 10), 1694 => to_unsigned(483, 10), 1695 => to_unsigned(462, 10), 1696 => to_unsigned(55, 10), 1697 => to_unsigned(769, 10), 1698 => to_unsigned(189, 10), 1699 => to_unsigned(659, 10), 1700 => to_unsigned(183, 10), 1701 => to_unsigned(754, 10), 1702 => to_unsigned(369, 10), 1703 => to_unsigned(698, 10), 1704 => to_unsigned(231, 10), 1705 => to_unsigned(864, 10), 1706 => to_unsigned(458, 10), 1707 => to_unsigned(527, 10), 1708 => to_unsigned(16, 10), 1709 => to_unsigned(413, 10), 1710 => to_unsigned(157, 10), 1711 => to_unsigned(43, 10), 1712 => to_unsigned(788, 10), 1713 => to_unsigned(441, 10), 1714 => to_unsigned(861, 10), 1715 => to_unsigned(215, 10), 1716 => to_unsigned(54, 10), 1717 => to_unsigned(173, 10), 1718 => to_unsigned(38, 10), 1719 => to_unsigned(115, 10), 1720 => to_unsigned(294, 10), 1721 => to_unsigned(862, 10), 1722 => to_unsigned(44, 10), 1723 => to_unsigned(278, 10), 1724 => to_unsigned(454, 10), 1725 => to_unsigned(1011, 10), 1726 => to_unsigned(782, 10), 1727 => to_unsigned(85, 10), 1728 => to_unsigned(69, 10), 1729 => to_unsigned(350, 10), 1730 => to_unsigned(344, 10), 1731 => to_unsigned(498, 10), 1732 => to_unsigned(199, 10), 1733 => to_unsigned(192, 10), 1734 => to_unsigned(124, 10), 1735 => to_unsigned(761, 10), 1736 => to_unsigned(816, 10), 1737 => to_unsigned(571, 10), 1738 => to_unsigned(63, 10), 1739 => to_unsigned(1004, 10), 1740 => to_unsigned(789, 10), 1741 => to_unsigned(174, 10), 1742 => to_unsigned(506, 10), 1743 => to_unsigned(337, 10), 1744 => to_unsigned(467, 10), 1745 => to_unsigned(783, 10), 1746 => to_unsigned(517, 10), 1747 => to_unsigned(680, 10), 1748 => to_unsigned(286, 10), 1749 => to_unsigned(177, 10), 1750 => to_unsigned(358, 10), 1751 => to_unsigned(557, 10), 1752 => to_unsigned(162, 10), 1753 => to_unsigned(709, 10), 1754 => to_unsigned(728, 10), 1755 => to_unsigned(981, 10), 1756 => to_unsigned(322, 10), 1757 => to_unsigned(296, 10), 1758 => to_unsigned(332, 10), 1759 => to_unsigned(229, 10), 1760 => to_unsigned(243, 10), 1761 => to_unsigned(672, 10), 1762 => to_unsigned(10, 10), 1763 => to_unsigned(847, 10), 1764 => to_unsigned(216, 10), 1765 => to_unsigned(379, 10), 1766 => to_unsigned(552, 10), 1767 => to_unsigned(1003, 10), 1768 => to_unsigned(23, 10), 1769 => to_unsigned(763, 10), 1770 => to_unsigned(665, 10), 1771 => to_unsigned(830, 10), 1772 => to_unsigned(774, 10), 1773 => to_unsigned(287, 10), 1774 => to_unsigned(619, 10), 1775 => to_unsigned(504, 10), 1776 => to_unsigned(607, 10), 1777 => to_unsigned(840, 10), 1778 => to_unsigned(135, 10), 1779 => to_unsigned(936, 10), 1780 => to_unsigned(676, 10), 1781 => to_unsigned(691, 10), 1782 => to_unsigned(529, 10), 1783 => to_unsigned(713, 10), 1784 => to_unsigned(830, 10), 1785 => to_unsigned(855, 10), 1786 => to_unsigned(366, 10), 1787 => to_unsigned(696, 10), 1788 => to_unsigned(1005, 10), 1789 => to_unsigned(25, 10), 1790 => to_unsigned(816, 10), 1791 => to_unsigned(283, 10), 1792 => to_unsigned(923, 10), 1793 => to_unsigned(13, 10), 1794 => to_unsigned(809, 10), 1795 => to_unsigned(489, 10), 1796 => to_unsigned(200, 10), 1797 => to_unsigned(669, 10), 1798 => to_unsigned(695, 10), 1799 => to_unsigned(809, 10), 1800 => to_unsigned(174, 10), 1801 => to_unsigned(315, 10), 1802 => to_unsigned(418, 10), 1803 => to_unsigned(30, 10), 1804 => to_unsigned(286, 10), 1805 => to_unsigned(788, 10), 1806 => to_unsigned(794, 10), 1807 => to_unsigned(235, 10), 1808 => to_unsigned(425, 10), 1809 => to_unsigned(268, 10), 1810 => to_unsigned(399, 10), 1811 => to_unsigned(119, 10), 1812 => to_unsigned(544, 10), 1813 => to_unsigned(344, 10), 1814 => to_unsigned(867, 10), 1815 => to_unsigned(835, 10), 1816 => to_unsigned(42, 10), 1817 => to_unsigned(772, 10), 1818 => to_unsigned(943, 10), 1819 => to_unsigned(615, 10), 1820 => to_unsigned(573, 10), 1821 => to_unsigned(149, 10), 1822 => to_unsigned(945, 10), 1823 => to_unsigned(555, 10), 1824 => to_unsigned(100, 10), 1825 => to_unsigned(607, 10), 1826 => to_unsigned(708, 10), 1827 => to_unsigned(338, 10), 1828 => to_unsigned(414, 10), 1829 => to_unsigned(664, 10), 1830 => to_unsigned(397, 10), 1831 => to_unsigned(925, 10), 1832 => to_unsigned(122, 10), 1833 => to_unsigned(798, 10), 1834 => to_unsigned(484, 10), 1835 => to_unsigned(665, 10), 1836 => to_unsigned(446, 10), 1837 => to_unsigned(690, 10), 1838 => to_unsigned(991, 10), 1839 => to_unsigned(833, 10), 1840 => to_unsigned(853, 10), 1841 => to_unsigned(134, 10), 1842 => to_unsigned(865, 10), 1843 => to_unsigned(37, 10), 1844 => to_unsigned(914, 10), 1845 => to_unsigned(281, 10), 1846 => to_unsigned(394, 10), 1847 => to_unsigned(71, 10), 1848 => to_unsigned(205, 10), 1849 => to_unsigned(229, 10), 1850 => to_unsigned(638, 10), 1851 => to_unsigned(721, 10), 1852 => to_unsigned(256, 10), 1853 => to_unsigned(401, 10), 1854 => to_unsigned(735, 10), 1855 => to_unsigned(175, 10), 1856 => to_unsigned(217, 10), 1857 => to_unsigned(327, 10), 1858 => to_unsigned(45, 10), 1859 => to_unsigned(51, 10), 1860 => to_unsigned(683, 10), 1861 => to_unsigned(912, 10), 1862 => to_unsigned(599, 10), 1863 => to_unsigned(871, 10), 1864 => to_unsigned(484, 10), 1865 => to_unsigned(902, 10), 1866 => to_unsigned(1021, 10), 1867 => to_unsigned(22, 10), 1868 => to_unsigned(587, 10), 1869 => to_unsigned(119, 10), 1870 => to_unsigned(338, 10), 1871 => to_unsigned(949, 10), 1872 => to_unsigned(618, 10), 1873 => to_unsigned(885, 10), 1874 => to_unsigned(831, 10), 1875 => to_unsigned(226, 10), 1876 => to_unsigned(438, 10), 1877 => to_unsigned(156, 10), 1878 => to_unsigned(285, 10), 1879 => to_unsigned(763, 10), 1880 => to_unsigned(733, 10), 1881 => to_unsigned(459, 10), 1882 => to_unsigned(44, 10), 1883 => to_unsigned(465, 10), 1884 => to_unsigned(437, 10), 1885 => to_unsigned(918, 10), 1886 => to_unsigned(162, 10), 1887 => to_unsigned(649, 10), 1888 => to_unsigned(513, 10), 1889 => to_unsigned(811, 10), 1890 => to_unsigned(92, 10), 1891 => to_unsigned(645, 10), 1892 => to_unsigned(264, 10), 1893 => to_unsigned(26, 10), 1894 => to_unsigned(6, 10), 1895 => to_unsigned(948, 10), 1896 => to_unsigned(73, 10), 1897 => to_unsigned(63, 10), 1898 => to_unsigned(477, 10), 1899 => to_unsigned(739, 10), 1900 => to_unsigned(748, 10), 1901 => to_unsigned(766, 10), 1902 => to_unsigned(285, 10), 1903 => to_unsigned(154, 10), 1904 => to_unsigned(449, 10), 1905 => to_unsigned(1015, 10), 1906 => to_unsigned(101, 10), 1907 => to_unsigned(402, 10), 1908 => to_unsigned(922, 10), 1909 => to_unsigned(483, 10), 1910 => to_unsigned(227, 10), 1911 => to_unsigned(855, 10), 1912 => to_unsigned(812, 10), 1913 => to_unsigned(667, 10), 1914 => to_unsigned(575, 10), 1915 => to_unsigned(683, 10), 1916 => to_unsigned(708, 10), 1917 => to_unsigned(66, 10), 1918 => to_unsigned(799, 10), 1919 => to_unsigned(953, 10), 1920 => to_unsigned(840, 10), 1921 => to_unsigned(521, 10), 1922 => to_unsigned(938, 10), 1923 => to_unsigned(916, 10), 1924 => to_unsigned(311, 10), 1925 => to_unsigned(160, 10), 1926 => to_unsigned(72, 10), 1927 => to_unsigned(892, 10), 1928 => to_unsigned(934, 10), 1929 => to_unsigned(760, 10), 1930 => to_unsigned(492, 10), 1931 => to_unsigned(985, 10), 1932 => to_unsigned(404, 10), 1933 => to_unsigned(402, 10), 1934 => to_unsigned(468, 10), 1935 => to_unsigned(174, 10), 1936 => to_unsigned(435, 10), 1937 => to_unsigned(923, 10), 1938 => to_unsigned(498, 10), 1939 => to_unsigned(305, 10), 1940 => to_unsigned(593, 10), 1941 => to_unsigned(153, 10), 1942 => to_unsigned(561, 10), 1943 => to_unsigned(902, 10), 1944 => to_unsigned(89, 10), 1945 => to_unsigned(549, 10), 1946 => to_unsigned(425, 10), 1947 => to_unsigned(582, 10), 1948 => to_unsigned(1003, 10), 1949 => to_unsigned(281, 10), 1950 => to_unsigned(1020, 10), 1951 => to_unsigned(464, 10), 1952 => to_unsigned(914, 10), 1953 => to_unsigned(314, 10), 1954 => to_unsigned(111, 10), 1955 => to_unsigned(618, 10), 1956 => to_unsigned(575, 10), 1957 => to_unsigned(334, 10), 1958 => to_unsigned(144, 10), 1959 => to_unsigned(275, 10), 1960 => to_unsigned(932, 10), 1961 => to_unsigned(453, 10), 1962 => to_unsigned(531, 10), 1963 => to_unsigned(682, 10), 1964 => to_unsigned(980, 10), 1965 => to_unsigned(845, 10), 1966 => to_unsigned(799, 10), 1967 => to_unsigned(525, 10), 1968 => to_unsigned(14, 10), 1969 => to_unsigned(908, 10), 1970 => to_unsigned(949, 10), 1971 => to_unsigned(54, 10), 1972 => to_unsigned(686, 10), 1973 => to_unsigned(79, 10), 1974 => to_unsigned(199, 10), 1975 => to_unsigned(23, 10), 1976 => to_unsigned(111, 10), 1977 => to_unsigned(242, 10), 1978 => to_unsigned(358, 10), 1979 => to_unsigned(329, 10), 1980 => to_unsigned(132, 10), 1981 => to_unsigned(614, 10), 1982 => to_unsigned(275, 10), 1983 => to_unsigned(231, 10), 1984 => to_unsigned(153, 10), 1985 => to_unsigned(528, 10), 1986 => to_unsigned(936, 10), 1987 => to_unsigned(684, 10), 1988 => to_unsigned(1017, 10), 1989 => to_unsigned(486, 10), 1990 => to_unsigned(456, 10), 1991 => to_unsigned(21, 10), 1992 => to_unsigned(879, 10), 1993 => to_unsigned(197, 10), 1994 => to_unsigned(427, 10), 1995 => to_unsigned(797, 10), 1996 => to_unsigned(875, 10), 1997 => to_unsigned(528, 10), 1998 => to_unsigned(796, 10), 1999 => to_unsigned(561, 10), 2000 => to_unsigned(924, 10), 2001 => to_unsigned(869, 10), 2002 => to_unsigned(263, 10), 2003 => to_unsigned(68, 10), 2004 => to_unsigned(811, 10), 2005 => to_unsigned(461, 10), 2006 => to_unsigned(379, 10), 2007 => to_unsigned(633, 10), 2008 => to_unsigned(42, 10), 2009 => to_unsigned(510, 10), 2010 => to_unsigned(920, 10), 2011 => to_unsigned(765, 10), 2012 => to_unsigned(189, 10), 2013 => to_unsigned(955, 10), 2014 => to_unsigned(129, 10), 2015 => to_unsigned(632, 10), 2016 => to_unsigned(96, 10), 2017 => to_unsigned(870, 10), 2018 => to_unsigned(379, 10), 2019 => to_unsigned(445, 10), 2020 => to_unsigned(432, 10), 2021 => to_unsigned(235, 10), 2022 => to_unsigned(910, 10), 2023 => to_unsigned(482, 10), 2024 => to_unsigned(479, 10), 2025 => to_unsigned(772, 10), 2026 => to_unsigned(473, 10), 2027 => to_unsigned(921, 10), 2028 => to_unsigned(167, 10), 2029 => to_unsigned(892, 10), 2030 => to_unsigned(6, 10), 2031 => to_unsigned(891, 10), 2032 => to_unsigned(57, 10), 2033 => to_unsigned(758, 10), 2034 => to_unsigned(234, 10), 2035 => to_unsigned(306, 10), 2036 => to_unsigned(735, 10), 2037 => to_unsigned(193, 10), 2038 => to_unsigned(514, 10), 2039 => to_unsigned(856, 10), 2040 => to_unsigned(951, 10), 2041 => to_unsigned(553, 10), 2042 => to_unsigned(879, 10), 2043 => to_unsigned(518, 10), 2044 => to_unsigned(237, 10), 2045 => to_unsigned(562, 10), 2046 => to_unsigned(571, 10), 2047 => to_unsigned(934, 10)),
            6 => (0 => to_unsigned(584, 10), 1 => to_unsigned(716, 10), 2 => to_unsigned(67, 10), 3 => to_unsigned(322, 10), 4 => to_unsigned(412, 10), 5 => to_unsigned(880, 10), 6 => to_unsigned(459, 10), 7 => to_unsigned(6, 10), 8 => to_unsigned(682, 10), 9 => to_unsigned(536, 10), 10 => to_unsigned(436, 10), 11 => to_unsigned(528, 10), 12 => to_unsigned(601, 10), 13 => to_unsigned(197, 10), 14 => to_unsigned(436, 10), 15 => to_unsigned(782, 10), 16 => to_unsigned(379, 10), 17 => to_unsigned(221, 10), 18 => to_unsigned(291, 10), 19 => to_unsigned(43, 10), 20 => to_unsigned(283, 10), 21 => to_unsigned(1021, 10), 22 => to_unsigned(620, 10), 23 => to_unsigned(311, 10), 24 => to_unsigned(637, 10), 25 => to_unsigned(496, 10), 26 => to_unsigned(326, 10), 27 => to_unsigned(441, 10), 28 => to_unsigned(936, 10), 29 => to_unsigned(701, 10), 30 => to_unsigned(167, 10), 31 => to_unsigned(816, 10), 32 => to_unsigned(387, 10), 33 => to_unsigned(182, 10), 34 => to_unsigned(907, 10), 35 => to_unsigned(34, 10), 36 => to_unsigned(710, 10), 37 => to_unsigned(486, 10), 38 => to_unsigned(704, 10), 39 => to_unsigned(482, 10), 40 => to_unsigned(613, 10), 41 => to_unsigned(798, 10), 42 => to_unsigned(17, 10), 43 => to_unsigned(75, 10), 44 => to_unsigned(74, 10), 45 => to_unsigned(1004, 10), 46 => to_unsigned(212, 10), 47 => to_unsigned(318, 10), 48 => to_unsigned(676, 10), 49 => to_unsigned(582, 10), 50 => to_unsigned(765, 10), 51 => to_unsigned(572, 10), 52 => to_unsigned(391, 10), 53 => to_unsigned(512, 10), 54 => to_unsigned(833, 10), 55 => to_unsigned(145, 10), 56 => to_unsigned(44, 10), 57 => to_unsigned(655, 10), 58 => to_unsigned(443, 10), 59 => to_unsigned(302, 10), 60 => to_unsigned(638, 10), 61 => to_unsigned(620, 10), 62 => to_unsigned(623, 10), 63 => to_unsigned(616, 10), 64 => to_unsigned(630, 10), 65 => to_unsigned(469, 10), 66 => to_unsigned(184, 10), 67 => to_unsigned(786, 10), 68 => to_unsigned(1014, 10), 69 => to_unsigned(166, 10), 70 => to_unsigned(710, 10), 71 => to_unsigned(662, 10), 72 => to_unsigned(22, 10), 73 => to_unsigned(50, 10), 74 => to_unsigned(196, 10), 75 => to_unsigned(215, 10), 76 => to_unsigned(848, 10), 77 => to_unsigned(84, 10), 78 => to_unsigned(319, 10), 79 => to_unsigned(898, 10), 80 => to_unsigned(326, 10), 81 => to_unsigned(438, 10), 82 => to_unsigned(33, 10), 83 => to_unsigned(898, 10), 84 => to_unsigned(981, 10), 85 => to_unsigned(383, 10), 86 => to_unsigned(842, 10), 87 => to_unsigned(363, 10), 88 => to_unsigned(445, 10), 89 => to_unsigned(553, 10), 90 => to_unsigned(294, 10), 91 => to_unsigned(244, 10), 92 => to_unsigned(991, 10), 93 => to_unsigned(741, 10), 94 => to_unsigned(114, 10), 95 => to_unsigned(66, 10), 96 => to_unsigned(107, 10), 97 => to_unsigned(938, 10), 98 => to_unsigned(953, 10), 99 => to_unsigned(548, 10), 100 => to_unsigned(965, 10), 101 => to_unsigned(452, 10), 102 => to_unsigned(189, 10), 103 => to_unsigned(237, 10), 104 => to_unsigned(953, 10), 105 => to_unsigned(894, 10), 106 => to_unsigned(1, 10), 107 => to_unsigned(14, 10), 108 => to_unsigned(31, 10), 109 => to_unsigned(125, 10), 110 => to_unsigned(825, 10), 111 => to_unsigned(194, 10), 112 => to_unsigned(561, 10), 113 => to_unsigned(952, 10), 114 => to_unsigned(379, 10), 115 => to_unsigned(821, 10), 116 => to_unsigned(269, 10), 117 => to_unsigned(793, 10), 118 => to_unsigned(4, 10), 119 => to_unsigned(823, 10), 120 => to_unsigned(666, 10), 121 => to_unsigned(40, 10), 122 => to_unsigned(782, 10), 123 => to_unsigned(774, 10), 124 => to_unsigned(814, 10), 125 => to_unsigned(741, 10), 126 => to_unsigned(611, 10), 127 => to_unsigned(475, 10), 128 => to_unsigned(252, 10), 129 => to_unsigned(827, 10), 130 => to_unsigned(887, 10), 131 => to_unsigned(374, 10), 132 => to_unsigned(614, 10), 133 => to_unsigned(897, 10), 134 => to_unsigned(91, 10), 135 => to_unsigned(809, 10), 136 => to_unsigned(507, 10), 137 => to_unsigned(727, 10), 138 => to_unsigned(953, 10), 139 => to_unsigned(227, 10), 140 => to_unsigned(253, 10), 141 => to_unsigned(798, 10), 142 => to_unsigned(564, 10), 143 => to_unsigned(352, 10), 144 => to_unsigned(117, 10), 145 => to_unsigned(673, 10), 146 => to_unsigned(160, 10), 147 => to_unsigned(590, 10), 148 => to_unsigned(196, 10), 149 => to_unsigned(798, 10), 150 => to_unsigned(53, 10), 151 => to_unsigned(28, 10), 152 => to_unsigned(818, 10), 153 => to_unsigned(885, 10), 154 => to_unsigned(28, 10), 155 => to_unsigned(526, 10), 156 => to_unsigned(901, 10), 157 => to_unsigned(289, 10), 158 => to_unsigned(332, 10), 159 => to_unsigned(174, 10), 160 => to_unsigned(862, 10), 161 => to_unsigned(245, 10), 162 => to_unsigned(447, 10), 163 => to_unsigned(913, 10), 164 => to_unsigned(806, 10), 165 => to_unsigned(77, 10), 166 => to_unsigned(99, 10), 167 => to_unsigned(27, 10), 168 => to_unsigned(931, 10), 169 => to_unsigned(654, 10), 170 => to_unsigned(98, 10), 171 => to_unsigned(285, 10), 172 => to_unsigned(258, 10), 173 => to_unsigned(278, 10), 174 => to_unsigned(773, 10), 175 => to_unsigned(849, 10), 176 => to_unsigned(684, 10), 177 => to_unsigned(335, 10), 178 => to_unsigned(185, 10), 179 => to_unsigned(341, 10), 180 => to_unsigned(784, 10), 181 => to_unsigned(847, 10), 182 => to_unsigned(859, 10), 183 => to_unsigned(973, 10), 184 => to_unsigned(582, 10), 185 => to_unsigned(67, 10), 186 => to_unsigned(9, 10), 187 => to_unsigned(819, 10), 188 => to_unsigned(571, 10), 189 => to_unsigned(860, 10), 190 => to_unsigned(589, 10), 191 => to_unsigned(996, 10), 192 => to_unsigned(266, 10), 193 => to_unsigned(863, 10), 194 => to_unsigned(701, 10), 195 => to_unsigned(884, 10), 196 => to_unsigned(908, 10), 197 => to_unsigned(423, 10), 198 => to_unsigned(116, 10), 199 => to_unsigned(702, 10), 200 => to_unsigned(642, 10), 201 => to_unsigned(28, 10), 202 => to_unsigned(217, 10), 203 => to_unsigned(404, 10), 204 => to_unsigned(176, 10), 205 => to_unsigned(560, 10), 206 => to_unsigned(559, 10), 207 => to_unsigned(202, 10), 208 => to_unsigned(780, 10), 209 => to_unsigned(863, 10), 210 => to_unsigned(71, 10), 211 => to_unsigned(74, 10), 212 => to_unsigned(833, 10), 213 => to_unsigned(341, 10), 214 => to_unsigned(988, 10), 215 => to_unsigned(510, 10), 216 => to_unsigned(832, 10), 217 => to_unsigned(459, 10), 218 => to_unsigned(483, 10), 219 => to_unsigned(54, 10), 220 => to_unsigned(901, 10), 221 => to_unsigned(230, 10), 222 => to_unsigned(770, 10), 223 => to_unsigned(1002, 10), 224 => to_unsigned(64, 10), 225 => to_unsigned(570, 10), 226 => to_unsigned(779, 10), 227 => to_unsigned(830, 10), 228 => to_unsigned(143, 10), 229 => to_unsigned(161, 10), 230 => to_unsigned(789, 10), 231 => to_unsigned(867, 10), 232 => to_unsigned(346, 10), 233 => to_unsigned(363, 10), 234 => to_unsigned(851, 10), 235 => to_unsigned(1023, 10), 236 => to_unsigned(574, 10), 237 => to_unsigned(453, 10), 238 => to_unsigned(882, 10), 239 => to_unsigned(901, 10), 240 => to_unsigned(661, 10), 241 => to_unsigned(995, 10), 242 => to_unsigned(856, 10), 243 => to_unsigned(595, 10), 244 => to_unsigned(813, 10), 245 => to_unsigned(540, 10), 246 => to_unsigned(563, 10), 247 => to_unsigned(959, 10), 248 => to_unsigned(96, 10), 249 => to_unsigned(728, 10), 250 => to_unsigned(128, 10), 251 => to_unsigned(730, 10), 252 => to_unsigned(765, 10), 253 => to_unsigned(108, 10), 254 => to_unsigned(954, 10), 255 => to_unsigned(413, 10), 256 => to_unsigned(522, 10), 257 => to_unsigned(827, 10), 258 => to_unsigned(654, 10), 259 => to_unsigned(415, 10), 260 => to_unsigned(638, 10), 261 => to_unsigned(279, 10), 262 => to_unsigned(711, 10), 263 => to_unsigned(284, 10), 264 => to_unsigned(638, 10), 265 => to_unsigned(948, 10), 266 => to_unsigned(620, 10), 267 => to_unsigned(709, 10), 268 => to_unsigned(84, 10), 269 => to_unsigned(855, 10), 270 => to_unsigned(758, 10), 271 => to_unsigned(986, 10), 272 => to_unsigned(24, 10), 273 => to_unsigned(416, 10), 274 => to_unsigned(522, 10), 275 => to_unsigned(129, 10), 276 => to_unsigned(325, 10), 277 => to_unsigned(818, 10), 278 => to_unsigned(125, 10), 279 => to_unsigned(471, 10), 280 => to_unsigned(467, 10), 281 => to_unsigned(465, 10), 282 => to_unsigned(108, 10), 283 => to_unsigned(421, 10), 284 => to_unsigned(703, 10), 285 => to_unsigned(404, 10), 286 => to_unsigned(32, 10), 287 => to_unsigned(869, 10), 288 => to_unsigned(622, 10), 289 => to_unsigned(931, 10), 290 => to_unsigned(321, 10), 291 => to_unsigned(641, 10), 292 => to_unsigned(1020, 10), 293 => to_unsigned(854, 10), 294 => to_unsigned(17, 10), 295 => to_unsigned(519, 10), 296 => to_unsigned(522, 10), 297 => to_unsigned(252, 10), 298 => to_unsigned(899, 10), 299 => to_unsigned(61, 10), 300 => to_unsigned(743, 10), 301 => to_unsigned(32, 10), 302 => to_unsigned(65, 10), 303 => to_unsigned(779, 10), 304 => to_unsigned(663, 10), 305 => to_unsigned(632, 10), 306 => to_unsigned(427, 10), 307 => to_unsigned(429, 10), 308 => to_unsigned(303, 10), 309 => to_unsigned(944, 10), 310 => to_unsigned(71, 10), 311 => to_unsigned(323, 10), 312 => to_unsigned(716, 10), 313 => to_unsigned(82, 10), 314 => to_unsigned(825, 10), 315 => to_unsigned(914, 10), 316 => to_unsigned(96, 10), 317 => to_unsigned(512, 10), 318 => to_unsigned(964, 10), 319 => to_unsigned(596, 10), 320 => to_unsigned(876, 10), 321 => to_unsigned(312, 10), 322 => to_unsigned(630, 10), 323 => to_unsigned(841, 10), 324 => to_unsigned(100, 10), 325 => to_unsigned(279, 10), 326 => to_unsigned(285, 10), 327 => to_unsigned(429, 10), 328 => to_unsigned(860, 10), 329 => to_unsigned(232, 10), 330 => to_unsigned(314, 10), 331 => to_unsigned(940, 10), 332 => to_unsigned(284, 10), 333 => to_unsigned(513, 10), 334 => to_unsigned(205, 10), 335 => to_unsigned(101, 10), 336 => to_unsigned(852, 10), 337 => to_unsigned(902, 10), 338 => to_unsigned(939, 10), 339 => to_unsigned(555, 10), 340 => to_unsigned(303, 10), 341 => to_unsigned(932, 10), 342 => to_unsigned(235, 10), 343 => to_unsigned(463, 10), 344 => to_unsigned(664, 10), 345 => to_unsigned(860, 10), 346 => to_unsigned(571, 10), 347 => to_unsigned(732, 10), 348 => to_unsigned(695, 10), 349 => to_unsigned(423, 10), 350 => to_unsigned(966, 10), 351 => to_unsigned(720, 10), 352 => to_unsigned(313, 10), 353 => to_unsigned(87, 10), 354 => to_unsigned(441, 10), 355 => to_unsigned(222, 10), 356 => to_unsigned(128, 10), 357 => to_unsigned(234, 10), 358 => to_unsigned(816, 10), 359 => to_unsigned(970, 10), 360 => to_unsigned(161, 10), 361 => to_unsigned(85, 10), 362 => to_unsigned(910, 10), 363 => to_unsigned(439, 10), 364 => to_unsigned(552, 10), 365 => to_unsigned(821, 10), 366 => to_unsigned(593, 10), 367 => to_unsigned(1004, 10), 368 => to_unsigned(694, 10), 369 => to_unsigned(1010, 10), 370 => to_unsigned(43, 10), 371 => to_unsigned(115, 10), 372 => to_unsigned(660, 10), 373 => to_unsigned(916, 10), 374 => to_unsigned(857, 10), 375 => to_unsigned(407, 10), 376 => to_unsigned(915, 10), 377 => to_unsigned(497, 10), 378 => to_unsigned(328, 10), 379 => to_unsigned(457, 10), 380 => to_unsigned(602, 10), 381 => to_unsigned(345, 10), 382 => to_unsigned(904, 10), 383 => to_unsigned(387, 10), 384 => to_unsigned(989, 10), 385 => to_unsigned(978, 10), 386 => to_unsigned(98, 10), 387 => to_unsigned(928, 10), 388 => to_unsigned(146, 10), 389 => to_unsigned(149, 10), 390 => to_unsigned(657, 10), 391 => to_unsigned(109, 10), 392 => to_unsigned(213, 10), 393 => to_unsigned(715, 10), 394 => to_unsigned(935, 10), 395 => to_unsigned(1002, 10), 396 => to_unsigned(277, 10), 397 => to_unsigned(70, 10), 398 => to_unsigned(1020, 10), 399 => to_unsigned(415, 10), 400 => to_unsigned(755, 10), 401 => to_unsigned(191, 10), 402 => to_unsigned(676, 10), 403 => to_unsigned(998, 10), 404 => to_unsigned(247, 10), 405 => to_unsigned(316, 10), 406 => to_unsigned(362, 10), 407 => to_unsigned(684, 10), 408 => to_unsigned(899, 10), 409 => to_unsigned(161, 10), 410 => to_unsigned(137, 10), 411 => to_unsigned(931, 10), 412 => to_unsigned(789, 10), 413 => to_unsigned(82, 10), 414 => to_unsigned(249, 10), 415 => to_unsigned(423, 10), 416 => to_unsigned(289, 10), 417 => to_unsigned(651, 10), 418 => to_unsigned(148, 10), 419 => to_unsigned(653, 10), 420 => to_unsigned(405, 10), 421 => to_unsigned(571, 10), 422 => to_unsigned(778, 10), 423 => to_unsigned(947, 10), 424 => to_unsigned(375, 10), 425 => to_unsigned(193, 10), 426 => to_unsigned(334, 10), 427 => to_unsigned(279, 10), 428 => to_unsigned(755, 10), 429 => to_unsigned(733, 10), 430 => to_unsigned(575, 10), 431 => to_unsigned(572, 10), 432 => to_unsigned(336, 10), 433 => to_unsigned(643, 10), 434 => to_unsigned(176, 10), 435 => to_unsigned(492, 10), 436 => to_unsigned(412, 10), 437 => to_unsigned(185, 10), 438 => to_unsigned(393, 10), 439 => to_unsigned(272, 10), 440 => to_unsigned(505, 10), 441 => to_unsigned(353, 10), 442 => to_unsigned(914, 10), 443 => to_unsigned(926, 10), 444 => to_unsigned(379, 10), 445 => to_unsigned(666, 10), 446 => to_unsigned(671, 10), 447 => to_unsigned(569, 10), 448 => to_unsigned(910, 10), 449 => to_unsigned(187, 10), 450 => to_unsigned(66, 10), 451 => to_unsigned(987, 10), 452 => to_unsigned(698, 10), 453 => to_unsigned(804, 10), 454 => to_unsigned(510, 10), 455 => to_unsigned(318, 10), 456 => to_unsigned(550, 10), 457 => to_unsigned(838, 10), 458 => to_unsigned(335, 10), 459 => to_unsigned(707, 10), 460 => to_unsigned(1012, 10), 461 => to_unsigned(481, 10), 462 => to_unsigned(673, 10), 463 => to_unsigned(499, 10), 464 => to_unsigned(611, 10), 465 => to_unsigned(219, 10), 466 => to_unsigned(161, 10), 467 => to_unsigned(175, 10), 468 => to_unsigned(319, 10), 469 => to_unsigned(227, 10), 470 => to_unsigned(530, 10), 471 => to_unsigned(785, 10), 472 => to_unsigned(225, 10), 473 => to_unsigned(241, 10), 474 => to_unsigned(808, 10), 475 => to_unsigned(145, 10), 476 => to_unsigned(708, 10), 477 => to_unsigned(873, 10), 478 => to_unsigned(539, 10), 479 => to_unsigned(212, 10), 480 => to_unsigned(77, 10), 481 => to_unsigned(142, 10), 482 => to_unsigned(415, 10), 483 => to_unsigned(314, 10), 484 => to_unsigned(843, 10), 485 => to_unsigned(892, 10), 486 => to_unsigned(880, 10), 487 => to_unsigned(466, 10), 488 => to_unsigned(405, 10), 489 => to_unsigned(87, 10), 490 => to_unsigned(276, 10), 491 => to_unsigned(976, 10), 492 => to_unsigned(875, 10), 493 => to_unsigned(307, 10), 494 => to_unsigned(452, 10), 495 => to_unsigned(837, 10), 496 => to_unsigned(771, 10), 497 => to_unsigned(313, 10), 498 => to_unsigned(636, 10), 499 => to_unsigned(456, 10), 500 => to_unsigned(285, 10), 501 => to_unsigned(881, 10), 502 => to_unsigned(609, 10), 503 => to_unsigned(949, 10), 504 => to_unsigned(830, 10), 505 => to_unsigned(412, 10), 506 => to_unsigned(659, 10), 507 => to_unsigned(64, 10), 508 => to_unsigned(428, 10), 509 => to_unsigned(850, 10), 510 => to_unsigned(885, 10), 511 => to_unsigned(924, 10), 512 => to_unsigned(98, 10), 513 => to_unsigned(807, 10), 514 => to_unsigned(234, 10), 515 => to_unsigned(89, 10), 516 => to_unsigned(518, 10), 517 => to_unsigned(637, 10), 518 => to_unsigned(971, 10), 519 => to_unsigned(772, 10), 520 => to_unsigned(500, 10), 521 => to_unsigned(711, 10), 522 => to_unsigned(442, 10), 523 => to_unsigned(96, 10), 524 => to_unsigned(708, 10), 525 => to_unsigned(109, 10), 526 => to_unsigned(458, 10), 527 => to_unsigned(460, 10), 528 => to_unsigned(502, 10), 529 => to_unsigned(156, 10), 530 => to_unsigned(273, 10), 531 => to_unsigned(820, 10), 532 => to_unsigned(109, 10), 533 => to_unsigned(266, 10), 534 => to_unsigned(557, 10), 535 => to_unsigned(493, 10), 536 => to_unsigned(981, 10), 537 => to_unsigned(450, 10), 538 => to_unsigned(255, 10), 539 => to_unsigned(355, 10), 540 => to_unsigned(544, 10), 541 => to_unsigned(239, 10), 542 => to_unsigned(307, 10), 543 => to_unsigned(449, 10), 544 => to_unsigned(245, 10), 545 => to_unsigned(491, 10), 546 => to_unsigned(747, 10), 547 => to_unsigned(262, 10), 548 => to_unsigned(987, 10), 549 => to_unsigned(471, 10), 550 => to_unsigned(695, 10), 551 => to_unsigned(987, 10), 552 => to_unsigned(888, 10), 553 => to_unsigned(272, 10), 554 => to_unsigned(824, 10), 555 => to_unsigned(637, 10), 556 => to_unsigned(278, 10), 557 => to_unsigned(538, 10), 558 => to_unsigned(172, 10), 559 => to_unsigned(759, 10), 560 => to_unsigned(436, 10), 561 => to_unsigned(590, 10), 562 => to_unsigned(466, 10), 563 => to_unsigned(144, 10), 564 => to_unsigned(712, 10), 565 => to_unsigned(401, 10), 566 => to_unsigned(156, 10), 567 => to_unsigned(547, 10), 568 => to_unsigned(410, 10), 569 => to_unsigned(812, 10), 570 => to_unsigned(72, 10), 571 => to_unsigned(994, 10), 572 => to_unsigned(381, 10), 573 => to_unsigned(814, 10), 574 => to_unsigned(226, 10), 575 => to_unsigned(98, 10), 576 => to_unsigned(672, 10), 577 => to_unsigned(851, 10), 578 => to_unsigned(703, 10), 579 => to_unsigned(617, 10), 580 => to_unsigned(108, 10), 581 => to_unsigned(689, 10), 582 => to_unsigned(44, 10), 583 => to_unsigned(536, 10), 584 => to_unsigned(577, 10), 585 => to_unsigned(500, 10), 586 => to_unsigned(994, 10), 587 => to_unsigned(671, 10), 588 => to_unsigned(419, 10), 589 => to_unsigned(721, 10), 590 => to_unsigned(198, 10), 591 => to_unsigned(190, 10), 592 => to_unsigned(423, 10), 593 => to_unsigned(257, 10), 594 => to_unsigned(969, 10), 595 => to_unsigned(399, 10), 596 => to_unsigned(994, 10), 597 => to_unsigned(431, 10), 598 => to_unsigned(850, 10), 599 => to_unsigned(800, 10), 600 => to_unsigned(630, 10), 601 => to_unsigned(98, 10), 602 => to_unsigned(503, 10), 603 => to_unsigned(633, 10), 604 => to_unsigned(797, 10), 605 => to_unsigned(224, 10), 606 => to_unsigned(284, 10), 607 => to_unsigned(522, 10), 608 => to_unsigned(215, 10), 609 => to_unsigned(953, 10), 610 => to_unsigned(127, 10), 611 => to_unsigned(287, 10), 612 => to_unsigned(711, 10), 613 => to_unsigned(559, 10), 614 => to_unsigned(855, 10), 615 => to_unsigned(416, 10), 616 => to_unsigned(280, 10), 617 => to_unsigned(121, 10), 618 => to_unsigned(420, 10), 619 => to_unsigned(297, 10), 620 => to_unsigned(749, 10), 621 => to_unsigned(823, 10), 622 => to_unsigned(823, 10), 623 => to_unsigned(453, 10), 624 => to_unsigned(733, 10), 625 => to_unsigned(1011, 10), 626 => to_unsigned(362, 10), 627 => to_unsigned(764, 10), 628 => to_unsigned(339, 10), 629 => to_unsigned(22, 10), 630 => to_unsigned(25, 10), 631 => to_unsigned(894, 10), 632 => to_unsigned(651, 10), 633 => to_unsigned(826, 10), 634 => to_unsigned(962, 10), 635 => to_unsigned(719, 10), 636 => to_unsigned(416, 10), 637 => to_unsigned(911, 10), 638 => to_unsigned(948, 10), 639 => to_unsigned(878, 10), 640 => to_unsigned(1023, 10), 641 => to_unsigned(627, 10), 642 => to_unsigned(992, 10), 643 => to_unsigned(66, 10), 644 => to_unsigned(911, 10), 645 => to_unsigned(982, 10), 646 => to_unsigned(527, 10), 647 => to_unsigned(492, 10), 648 => to_unsigned(742, 10), 649 => to_unsigned(254, 10), 650 => to_unsigned(998, 10), 651 => to_unsigned(596, 10), 652 => to_unsigned(284, 10), 653 => to_unsigned(364, 10), 654 => to_unsigned(263, 10), 655 => to_unsigned(578, 10), 656 => to_unsigned(143, 10), 657 => to_unsigned(550, 10), 658 => to_unsigned(69, 10), 659 => to_unsigned(678, 10), 660 => to_unsigned(370, 10), 661 => to_unsigned(855, 10), 662 => to_unsigned(553, 10), 663 => to_unsigned(405, 10), 664 => to_unsigned(138, 10), 665 => to_unsigned(370, 10), 666 => to_unsigned(150, 10), 667 => to_unsigned(327, 10), 668 => to_unsigned(409, 10), 669 => to_unsigned(762, 10), 670 => to_unsigned(103, 10), 671 => to_unsigned(318, 10), 672 => to_unsigned(504, 10), 673 => to_unsigned(649, 10), 674 => to_unsigned(996, 10), 675 => to_unsigned(433, 10), 676 => to_unsigned(744, 10), 677 => to_unsigned(808, 10), 678 => to_unsigned(553, 10), 679 => to_unsigned(917, 10), 680 => to_unsigned(184, 10), 681 => to_unsigned(697, 10), 682 => to_unsigned(821, 10), 683 => to_unsigned(529, 10), 684 => to_unsigned(761, 10), 685 => to_unsigned(651, 10), 686 => to_unsigned(1015, 10), 687 => to_unsigned(221, 10), 688 => to_unsigned(506, 10), 689 => to_unsigned(233, 10), 690 => to_unsigned(762, 10), 691 => to_unsigned(289, 10), 692 => to_unsigned(149, 10), 693 => to_unsigned(415, 10), 694 => to_unsigned(909, 10), 695 => to_unsigned(115, 10), 696 => to_unsigned(701, 10), 697 => to_unsigned(451, 10), 698 => to_unsigned(505, 10), 699 => to_unsigned(366, 10), 700 => to_unsigned(850, 10), 701 => to_unsigned(701, 10), 702 => to_unsigned(674, 10), 703 => to_unsigned(189, 10), 704 => to_unsigned(593, 10), 705 => to_unsigned(95, 10), 706 => to_unsigned(419, 10), 707 => to_unsigned(14, 10), 708 => to_unsigned(408, 10), 709 => to_unsigned(354, 10), 710 => to_unsigned(378, 10), 711 => to_unsigned(172, 10), 712 => to_unsigned(74, 10), 713 => to_unsigned(726, 10), 714 => to_unsigned(209, 10), 715 => to_unsigned(58, 10), 716 => to_unsigned(697, 10), 717 => to_unsigned(247, 10), 718 => to_unsigned(307, 10), 719 => to_unsigned(1014, 10), 720 => to_unsigned(426, 10), 721 => to_unsigned(109, 10), 722 => to_unsigned(793, 10), 723 => to_unsigned(524, 10), 724 => to_unsigned(857, 10), 725 => to_unsigned(409, 10), 726 => to_unsigned(701, 10), 727 => to_unsigned(480, 10), 728 => to_unsigned(500, 10), 729 => to_unsigned(630, 10), 730 => to_unsigned(903, 10), 731 => to_unsigned(284, 10), 732 => to_unsigned(716, 10), 733 => to_unsigned(320, 10), 734 => to_unsigned(811, 10), 735 => to_unsigned(986, 10), 736 => to_unsigned(243, 10), 737 => to_unsigned(347, 10), 738 => to_unsigned(118, 10), 739 => to_unsigned(405, 10), 740 => to_unsigned(179, 10), 741 => to_unsigned(239, 10), 742 => to_unsigned(744, 10), 743 => to_unsigned(333, 10), 744 => to_unsigned(841, 10), 745 => to_unsigned(77, 10), 746 => to_unsigned(1023, 10), 747 => to_unsigned(315, 10), 748 => to_unsigned(691, 10), 749 => to_unsigned(976, 10), 750 => to_unsigned(235, 10), 751 => to_unsigned(121, 10), 752 => to_unsigned(680, 10), 753 => to_unsigned(423, 10), 754 => to_unsigned(372, 10), 755 => to_unsigned(125, 10), 756 => to_unsigned(127, 10), 757 => to_unsigned(277, 10), 758 => to_unsigned(513, 10), 759 => to_unsigned(82, 10), 760 => to_unsigned(937, 10), 761 => to_unsigned(505, 10), 762 => to_unsigned(452, 10), 763 => to_unsigned(303, 10), 764 => to_unsigned(902, 10), 765 => to_unsigned(561, 10), 766 => to_unsigned(742, 10), 767 => to_unsigned(866, 10), 768 => to_unsigned(229, 10), 769 => to_unsigned(229, 10), 770 => to_unsigned(435, 10), 771 => to_unsigned(65, 10), 772 => to_unsigned(383, 10), 773 => to_unsigned(700, 10), 774 => to_unsigned(996, 10), 775 => to_unsigned(61, 10), 776 => to_unsigned(953, 10), 777 => to_unsigned(220, 10), 778 => to_unsigned(375, 10), 779 => to_unsigned(706, 10), 780 => to_unsigned(995, 10), 781 => to_unsigned(330, 10), 782 => to_unsigned(317, 10), 783 => to_unsigned(541, 10), 784 => to_unsigned(47, 10), 785 => to_unsigned(8, 10), 786 => to_unsigned(637, 10), 787 => to_unsigned(54, 10), 788 => to_unsigned(483, 10), 789 => to_unsigned(190, 10), 790 => to_unsigned(491, 10), 791 => to_unsigned(319, 10), 792 => to_unsigned(824, 10), 793 => to_unsigned(990, 10), 794 => to_unsigned(504, 10), 795 => to_unsigned(136, 10), 796 => to_unsigned(455, 10), 797 => to_unsigned(964, 10), 798 => to_unsigned(564, 10), 799 => to_unsigned(783, 10), 800 => to_unsigned(215, 10), 801 => to_unsigned(390, 10), 802 => to_unsigned(778, 10), 803 => to_unsigned(98, 10), 804 => to_unsigned(269, 10), 805 => to_unsigned(234, 10), 806 => to_unsigned(690, 10), 807 => to_unsigned(846, 10), 808 => to_unsigned(649, 10), 809 => to_unsigned(991, 10), 810 => to_unsigned(200, 10), 811 => to_unsigned(62, 10), 812 => to_unsigned(357, 10), 813 => to_unsigned(15, 10), 814 => to_unsigned(635, 10), 815 => to_unsigned(375, 10), 816 => to_unsigned(696, 10), 817 => to_unsigned(1013, 10), 818 => to_unsigned(994, 10), 819 => to_unsigned(508, 10), 820 => to_unsigned(124, 10), 821 => to_unsigned(280, 10), 822 => to_unsigned(690, 10), 823 => to_unsigned(813, 10), 824 => to_unsigned(906, 10), 825 => to_unsigned(658, 10), 826 => to_unsigned(989, 10), 827 => to_unsigned(255, 10), 828 => to_unsigned(560, 10), 829 => to_unsigned(1003, 10), 830 => to_unsigned(235, 10), 831 => to_unsigned(904, 10), 832 => to_unsigned(758, 10), 833 => to_unsigned(344, 10), 834 => to_unsigned(364, 10), 835 => to_unsigned(110, 10), 836 => to_unsigned(218, 10), 837 => to_unsigned(772, 10), 838 => to_unsigned(898, 10), 839 => to_unsigned(223, 10), 840 => to_unsigned(635, 10), 841 => to_unsigned(757, 10), 842 => to_unsigned(608, 10), 843 => to_unsigned(429, 10), 844 => to_unsigned(110, 10), 845 => to_unsigned(262, 10), 846 => to_unsigned(646, 10), 847 => to_unsigned(399, 10), 848 => to_unsigned(773, 10), 849 => to_unsigned(839, 10), 850 => to_unsigned(702, 10), 851 => to_unsigned(500, 10), 852 => to_unsigned(83, 10), 853 => to_unsigned(339, 10), 854 => to_unsigned(524, 10), 855 => to_unsigned(305, 10), 856 => to_unsigned(238, 10), 857 => to_unsigned(478, 10), 858 => to_unsigned(642, 10), 859 => to_unsigned(372, 10), 860 => to_unsigned(580, 10), 861 => to_unsigned(776, 10), 862 => to_unsigned(211, 10), 863 => to_unsigned(528, 10), 864 => to_unsigned(226, 10), 865 => to_unsigned(697, 10), 866 => to_unsigned(345, 10), 867 => to_unsigned(492, 10), 868 => to_unsigned(406, 10), 869 => to_unsigned(79, 10), 870 => to_unsigned(924, 10), 871 => to_unsigned(428, 10), 872 => to_unsigned(49, 10), 873 => to_unsigned(219, 10), 874 => to_unsigned(776, 10), 875 => to_unsigned(417, 10), 876 => to_unsigned(897, 10), 877 => to_unsigned(574, 10), 878 => to_unsigned(382, 10), 879 => to_unsigned(540, 10), 880 => to_unsigned(406, 10), 881 => to_unsigned(91, 10), 882 => to_unsigned(959, 10), 883 => to_unsigned(90, 10), 884 => to_unsigned(959, 10), 885 => to_unsigned(293, 10), 886 => to_unsigned(725, 10), 887 => to_unsigned(761, 10), 888 => to_unsigned(571, 10), 889 => to_unsigned(914, 10), 890 => to_unsigned(580, 10), 891 => to_unsigned(326, 10), 892 => to_unsigned(400, 10), 893 => to_unsigned(305, 10), 894 => to_unsigned(451, 10), 895 => to_unsigned(394, 10), 896 => to_unsigned(591, 10), 897 => to_unsigned(761, 10), 898 => to_unsigned(295, 10), 899 => to_unsigned(310, 10), 900 => to_unsigned(542, 10), 901 => to_unsigned(248, 10), 902 => to_unsigned(204, 10), 903 => to_unsigned(937, 10), 904 => to_unsigned(189, 10), 905 => to_unsigned(354, 10), 906 => to_unsigned(420, 10), 907 => to_unsigned(846, 10), 908 => to_unsigned(485, 10), 909 => to_unsigned(885, 10), 910 => to_unsigned(671, 10), 911 => to_unsigned(712, 10), 912 => to_unsigned(112, 10), 913 => to_unsigned(843, 10), 914 => to_unsigned(163, 10), 915 => to_unsigned(847, 10), 916 => to_unsigned(528, 10), 917 => to_unsigned(904, 10), 918 => to_unsigned(911, 10), 919 => to_unsigned(599, 10), 920 => to_unsigned(695, 10), 921 => to_unsigned(52, 10), 922 => to_unsigned(315, 10), 923 => to_unsigned(880, 10), 924 => to_unsigned(409, 10), 925 => to_unsigned(684, 10), 926 => to_unsigned(595, 10), 927 => to_unsigned(466, 10), 928 => to_unsigned(663, 10), 929 => to_unsigned(541, 10), 930 => to_unsigned(443, 10), 931 => to_unsigned(760, 10), 932 => to_unsigned(71, 10), 933 => to_unsigned(275, 10), 934 => to_unsigned(69, 10), 935 => to_unsigned(5, 10), 936 => to_unsigned(810, 10), 937 => to_unsigned(556, 10), 938 => to_unsigned(2, 10), 939 => to_unsigned(683, 10), 940 => to_unsigned(623, 10), 941 => to_unsigned(399, 10), 942 => to_unsigned(101, 10), 943 => to_unsigned(565, 10), 944 => to_unsigned(637, 10), 945 => to_unsigned(392, 10), 946 => to_unsigned(696, 10), 947 => to_unsigned(724, 10), 948 => to_unsigned(332, 10), 949 => to_unsigned(704, 10), 950 => to_unsigned(469, 10), 951 => to_unsigned(371, 10), 952 => to_unsigned(96, 10), 953 => to_unsigned(502, 10), 954 => to_unsigned(130, 10), 955 => to_unsigned(901, 10), 956 => to_unsigned(629, 10), 957 => to_unsigned(159, 10), 958 => to_unsigned(754, 10), 959 => to_unsigned(204, 10), 960 => to_unsigned(599, 10), 961 => to_unsigned(525, 10), 962 => to_unsigned(472, 10), 963 => to_unsigned(457, 10), 964 => to_unsigned(181, 10), 965 => to_unsigned(687, 10), 966 => to_unsigned(395, 10), 967 => to_unsigned(56, 10), 968 => to_unsigned(761, 10), 969 => to_unsigned(86, 10), 970 => to_unsigned(414, 10), 971 => to_unsigned(586, 10), 972 => to_unsigned(547, 10), 973 => to_unsigned(342, 10), 974 => to_unsigned(236, 10), 975 => to_unsigned(362, 10), 976 => to_unsigned(788, 10), 977 => to_unsigned(307, 10), 978 => to_unsigned(191, 10), 979 => to_unsigned(894, 10), 980 => to_unsigned(416, 10), 981 => to_unsigned(700, 10), 982 => to_unsigned(986, 10), 983 => to_unsigned(410, 10), 984 => to_unsigned(173, 10), 985 => to_unsigned(328, 10), 986 => to_unsigned(636, 10), 987 => to_unsigned(720, 10), 988 => to_unsigned(142, 10), 989 => to_unsigned(709, 10), 990 => to_unsigned(941, 10), 991 => to_unsigned(841, 10), 992 => to_unsigned(14, 10), 993 => to_unsigned(475, 10), 994 => to_unsigned(979, 10), 995 => to_unsigned(814, 10), 996 => to_unsigned(818, 10), 997 => to_unsigned(606, 10), 998 => to_unsigned(73, 10), 999 => to_unsigned(291, 10), 1000 => to_unsigned(137, 10), 1001 => to_unsigned(843, 10), 1002 => to_unsigned(614, 10), 1003 => to_unsigned(1009, 10), 1004 => to_unsigned(975, 10), 1005 => to_unsigned(825, 10), 1006 => to_unsigned(428, 10), 1007 => to_unsigned(298, 10), 1008 => to_unsigned(974, 10), 1009 => to_unsigned(525, 10), 1010 => to_unsigned(123, 10), 1011 => to_unsigned(703, 10), 1012 => to_unsigned(473, 10), 1013 => to_unsigned(470, 10), 1014 => to_unsigned(596, 10), 1015 => to_unsigned(986, 10), 1016 => to_unsigned(734, 10), 1017 => to_unsigned(799, 10), 1018 => to_unsigned(949, 10), 1019 => to_unsigned(815, 10), 1020 => to_unsigned(992, 10), 1021 => to_unsigned(882, 10), 1022 => to_unsigned(7, 10), 1023 => to_unsigned(555, 10), 1024 => to_unsigned(859, 10), 1025 => to_unsigned(418, 10), 1026 => to_unsigned(585, 10), 1027 => to_unsigned(989, 10), 1028 => to_unsigned(403, 10), 1029 => to_unsigned(830, 10), 1030 => to_unsigned(281, 10), 1031 => to_unsigned(285, 10), 1032 => to_unsigned(948, 10), 1033 => to_unsigned(428, 10), 1034 => to_unsigned(565, 10), 1035 => to_unsigned(811, 10), 1036 => to_unsigned(18, 10), 1037 => to_unsigned(25, 10), 1038 => to_unsigned(1021, 10), 1039 => to_unsigned(735, 10), 1040 => to_unsigned(359, 10), 1041 => to_unsigned(661, 10), 1042 => to_unsigned(706, 10), 1043 => to_unsigned(665, 10), 1044 => to_unsigned(193, 10), 1045 => to_unsigned(610, 10), 1046 => to_unsigned(212, 10), 1047 => to_unsigned(747, 10), 1048 => to_unsigned(877, 10), 1049 => to_unsigned(838, 10), 1050 => to_unsigned(338, 10), 1051 => to_unsigned(254, 10), 1052 => to_unsigned(271, 10), 1053 => to_unsigned(88, 10), 1054 => to_unsigned(633, 10), 1055 => to_unsigned(442, 10), 1056 => to_unsigned(314, 10), 1057 => to_unsigned(180, 10), 1058 => to_unsigned(1019, 10), 1059 => to_unsigned(478, 10), 1060 => to_unsigned(897, 10), 1061 => to_unsigned(586, 10), 1062 => to_unsigned(615, 10), 1063 => to_unsigned(255, 10), 1064 => to_unsigned(525, 10), 1065 => to_unsigned(669, 10), 1066 => to_unsigned(44, 10), 1067 => to_unsigned(919, 10), 1068 => to_unsigned(116, 10), 1069 => to_unsigned(709, 10), 1070 => to_unsigned(578, 10), 1071 => to_unsigned(978, 10), 1072 => to_unsigned(608, 10), 1073 => to_unsigned(345, 10), 1074 => to_unsigned(581, 10), 1075 => to_unsigned(655, 10), 1076 => to_unsigned(102, 10), 1077 => to_unsigned(806, 10), 1078 => to_unsigned(819, 10), 1079 => to_unsigned(144, 10), 1080 => to_unsigned(457, 10), 1081 => to_unsigned(287, 10), 1082 => to_unsigned(1002, 10), 1083 => to_unsigned(877, 10), 1084 => to_unsigned(215, 10), 1085 => to_unsigned(328, 10), 1086 => to_unsigned(867, 10), 1087 => to_unsigned(920, 10), 1088 => to_unsigned(959, 10), 1089 => to_unsigned(861, 10), 1090 => to_unsigned(265, 10), 1091 => to_unsigned(643, 10), 1092 => to_unsigned(266, 10), 1093 => to_unsigned(882, 10), 1094 => to_unsigned(587, 10), 1095 => to_unsigned(330, 10), 1096 => to_unsigned(165, 10), 1097 => to_unsigned(113, 10), 1098 => to_unsigned(401, 10), 1099 => to_unsigned(734, 10), 1100 => to_unsigned(991, 10), 1101 => to_unsigned(737, 10), 1102 => to_unsigned(358, 10), 1103 => to_unsigned(222, 10), 1104 => to_unsigned(490, 10), 1105 => to_unsigned(600, 10), 1106 => to_unsigned(322, 10), 1107 => to_unsigned(708, 10), 1108 => to_unsigned(726, 10), 1109 => to_unsigned(744, 10), 1110 => to_unsigned(894, 10), 1111 => to_unsigned(850, 10), 1112 => to_unsigned(547, 10), 1113 => to_unsigned(157, 10), 1114 => to_unsigned(569, 10), 1115 => to_unsigned(674, 10), 1116 => to_unsigned(212, 10), 1117 => to_unsigned(1007, 10), 1118 => to_unsigned(994, 10), 1119 => to_unsigned(893, 10), 1120 => to_unsigned(982, 10), 1121 => to_unsigned(912, 10), 1122 => to_unsigned(743, 10), 1123 => to_unsigned(185, 10), 1124 => to_unsigned(434, 10), 1125 => to_unsigned(294, 10), 1126 => to_unsigned(738, 10), 1127 => to_unsigned(951, 10), 1128 => to_unsigned(410, 10), 1129 => to_unsigned(226, 10), 1130 => to_unsigned(992, 10), 1131 => to_unsigned(119, 10), 1132 => to_unsigned(665, 10), 1133 => to_unsigned(288, 10), 1134 => to_unsigned(240, 10), 1135 => to_unsigned(300, 10), 1136 => to_unsigned(1004, 10), 1137 => to_unsigned(128, 10), 1138 => to_unsigned(217, 10), 1139 => to_unsigned(342, 10), 1140 => to_unsigned(48, 10), 1141 => to_unsigned(797, 10), 1142 => to_unsigned(420, 10), 1143 => to_unsigned(475, 10), 1144 => to_unsigned(924, 10), 1145 => to_unsigned(656, 10), 1146 => to_unsigned(8, 10), 1147 => to_unsigned(848, 10), 1148 => to_unsigned(546, 10), 1149 => to_unsigned(996, 10), 1150 => to_unsigned(686, 10), 1151 => to_unsigned(160, 10), 1152 => to_unsigned(316, 10), 1153 => to_unsigned(982, 10), 1154 => to_unsigned(277, 10), 1155 => to_unsigned(171, 10), 1156 => to_unsigned(224, 10), 1157 => to_unsigned(426, 10), 1158 => to_unsigned(479, 10), 1159 => to_unsigned(119, 10), 1160 => to_unsigned(998, 10), 1161 => to_unsigned(365, 10), 1162 => to_unsigned(193, 10), 1163 => to_unsigned(46, 10), 1164 => to_unsigned(962, 10), 1165 => to_unsigned(795, 10), 1166 => to_unsigned(329, 10), 1167 => to_unsigned(433, 10), 1168 => to_unsigned(732, 10), 1169 => to_unsigned(21, 10), 1170 => to_unsigned(635, 10), 1171 => to_unsigned(356, 10), 1172 => to_unsigned(786, 10), 1173 => to_unsigned(870, 10), 1174 => to_unsigned(870, 10), 1175 => to_unsigned(972, 10), 1176 => to_unsigned(209, 10), 1177 => to_unsigned(546, 10), 1178 => to_unsigned(484, 10), 1179 => to_unsigned(99, 10), 1180 => to_unsigned(178, 10), 1181 => to_unsigned(758, 10), 1182 => to_unsigned(408, 10), 1183 => to_unsigned(1008, 10), 1184 => to_unsigned(540, 10), 1185 => to_unsigned(488, 10), 1186 => to_unsigned(792, 10), 1187 => to_unsigned(866, 10), 1188 => to_unsigned(871, 10), 1189 => to_unsigned(540, 10), 1190 => to_unsigned(478, 10), 1191 => to_unsigned(151, 10), 1192 => to_unsigned(624, 10), 1193 => to_unsigned(453, 10), 1194 => to_unsigned(325, 10), 1195 => to_unsigned(673, 10), 1196 => to_unsigned(674, 10), 1197 => to_unsigned(739, 10), 1198 => to_unsigned(945, 10), 1199 => to_unsigned(118, 10), 1200 => to_unsigned(948, 10), 1201 => to_unsigned(820, 10), 1202 => to_unsigned(63, 10), 1203 => to_unsigned(979, 10), 1204 => to_unsigned(1012, 10), 1205 => to_unsigned(429, 10), 1206 => to_unsigned(124, 10), 1207 => to_unsigned(276, 10), 1208 => to_unsigned(728, 10), 1209 => to_unsigned(636, 10), 1210 => to_unsigned(811, 10), 1211 => to_unsigned(947, 10), 1212 => to_unsigned(91, 10), 1213 => to_unsigned(103, 10), 1214 => to_unsigned(333, 10), 1215 => to_unsigned(404, 10), 1216 => to_unsigned(436, 10), 1217 => to_unsigned(180, 10), 1218 => to_unsigned(1006, 10), 1219 => to_unsigned(678, 10), 1220 => to_unsigned(1002, 10), 1221 => to_unsigned(618, 10), 1222 => to_unsigned(134, 10), 1223 => to_unsigned(442, 10), 1224 => to_unsigned(344, 10), 1225 => to_unsigned(144, 10), 1226 => to_unsigned(839, 10), 1227 => to_unsigned(786, 10), 1228 => to_unsigned(755, 10), 1229 => to_unsigned(370, 10), 1230 => to_unsigned(253, 10), 1231 => to_unsigned(279, 10), 1232 => to_unsigned(786, 10), 1233 => to_unsigned(254, 10), 1234 => to_unsigned(60, 10), 1235 => to_unsigned(38, 10), 1236 => to_unsigned(309, 10), 1237 => to_unsigned(304, 10), 1238 => to_unsigned(178, 10), 1239 => to_unsigned(797, 10), 1240 => to_unsigned(300, 10), 1241 => to_unsigned(753, 10), 1242 => to_unsigned(604, 10), 1243 => to_unsigned(790, 10), 1244 => to_unsigned(641, 10), 1245 => to_unsigned(185, 10), 1246 => to_unsigned(534, 10), 1247 => to_unsigned(594, 10), 1248 => to_unsigned(205, 10), 1249 => to_unsigned(126, 10), 1250 => to_unsigned(830, 10), 1251 => to_unsigned(1021, 10), 1252 => to_unsigned(303, 10), 1253 => to_unsigned(347, 10), 1254 => to_unsigned(232, 10), 1255 => to_unsigned(496, 10), 1256 => to_unsigned(85, 10), 1257 => to_unsigned(834, 10), 1258 => to_unsigned(595, 10), 1259 => to_unsigned(553, 10), 1260 => to_unsigned(435, 10), 1261 => to_unsigned(244, 10), 1262 => to_unsigned(553, 10), 1263 => to_unsigned(775, 10), 1264 => to_unsigned(580, 10), 1265 => to_unsigned(66, 10), 1266 => to_unsigned(995, 10), 1267 => to_unsigned(319, 10), 1268 => to_unsigned(397, 10), 1269 => to_unsigned(632, 10), 1270 => to_unsigned(748, 10), 1271 => to_unsigned(113, 10), 1272 => to_unsigned(412, 10), 1273 => to_unsigned(38, 10), 1274 => to_unsigned(260, 10), 1275 => to_unsigned(422, 10), 1276 => to_unsigned(445, 10), 1277 => to_unsigned(779, 10), 1278 => to_unsigned(902, 10), 1279 => to_unsigned(335, 10), 1280 => to_unsigned(832, 10), 1281 => to_unsigned(731, 10), 1282 => to_unsigned(674, 10), 1283 => to_unsigned(111, 10), 1284 => to_unsigned(354, 10), 1285 => to_unsigned(321, 10), 1286 => to_unsigned(789, 10), 1287 => to_unsigned(665, 10), 1288 => to_unsigned(69, 10), 1289 => to_unsigned(616, 10), 1290 => to_unsigned(791, 10), 1291 => to_unsigned(594, 10), 1292 => to_unsigned(155, 10), 1293 => to_unsigned(38, 10), 1294 => to_unsigned(307, 10), 1295 => to_unsigned(524, 10), 1296 => to_unsigned(917, 10), 1297 => to_unsigned(353, 10), 1298 => to_unsigned(685, 10), 1299 => to_unsigned(648, 10), 1300 => to_unsigned(641, 10), 1301 => to_unsigned(412, 10), 1302 => to_unsigned(947, 10), 1303 => to_unsigned(430, 10), 1304 => to_unsigned(351, 10), 1305 => to_unsigned(261, 10), 1306 => to_unsigned(607, 10), 1307 => to_unsigned(358, 10), 1308 => to_unsigned(785, 10), 1309 => to_unsigned(631, 10), 1310 => to_unsigned(941, 10), 1311 => to_unsigned(290, 10), 1312 => to_unsigned(445, 10), 1313 => to_unsigned(859, 10), 1314 => to_unsigned(396, 10), 1315 => to_unsigned(484, 10), 1316 => to_unsigned(214, 10), 1317 => to_unsigned(864, 10), 1318 => to_unsigned(342, 10), 1319 => to_unsigned(692, 10), 1320 => to_unsigned(266, 10), 1321 => to_unsigned(556, 10), 1322 => to_unsigned(880, 10), 1323 => to_unsigned(81, 10), 1324 => to_unsigned(902, 10), 1325 => to_unsigned(874, 10), 1326 => to_unsigned(231, 10), 1327 => to_unsigned(170, 10), 1328 => to_unsigned(601, 10), 1329 => to_unsigned(548, 10), 1330 => to_unsigned(609, 10), 1331 => to_unsigned(816, 10), 1332 => to_unsigned(410, 10), 1333 => to_unsigned(916, 10), 1334 => to_unsigned(147, 10), 1335 => to_unsigned(640, 10), 1336 => to_unsigned(868, 10), 1337 => to_unsigned(93, 10), 1338 => to_unsigned(204, 10), 1339 => to_unsigned(697, 10), 1340 => to_unsigned(231, 10), 1341 => to_unsigned(229, 10), 1342 => to_unsigned(852, 10), 1343 => to_unsigned(563, 10), 1344 => to_unsigned(748, 10), 1345 => to_unsigned(869, 10), 1346 => to_unsigned(753, 10), 1347 => to_unsigned(383, 10), 1348 => to_unsigned(292, 10), 1349 => to_unsigned(247, 10), 1350 => to_unsigned(746, 10), 1351 => to_unsigned(73, 10), 1352 => to_unsigned(944, 10), 1353 => to_unsigned(530, 10), 1354 => to_unsigned(455, 10), 1355 => to_unsigned(843, 10), 1356 => to_unsigned(677, 10), 1357 => to_unsigned(657, 10), 1358 => to_unsigned(845, 10), 1359 => to_unsigned(138, 10), 1360 => to_unsigned(346, 10), 1361 => to_unsigned(238, 10), 1362 => to_unsigned(177, 10), 1363 => to_unsigned(891, 10), 1364 => to_unsigned(39, 10), 1365 => to_unsigned(109, 10), 1366 => to_unsigned(24, 10), 1367 => to_unsigned(448, 10), 1368 => to_unsigned(185, 10), 1369 => to_unsigned(364, 10), 1370 => to_unsigned(546, 10), 1371 => to_unsigned(949, 10), 1372 => to_unsigned(939, 10), 1373 => to_unsigned(218, 10), 1374 => to_unsigned(117, 10), 1375 => to_unsigned(252, 10), 1376 => to_unsigned(707, 10), 1377 => to_unsigned(327, 10), 1378 => to_unsigned(286, 10), 1379 => to_unsigned(162, 10), 1380 => to_unsigned(529, 10), 1381 => to_unsigned(780, 10), 1382 => to_unsigned(846, 10), 1383 => to_unsigned(562, 10), 1384 => to_unsigned(186, 10), 1385 => to_unsigned(265, 10), 1386 => to_unsigned(580, 10), 1387 => to_unsigned(377, 10), 1388 => to_unsigned(575, 10), 1389 => to_unsigned(505, 10), 1390 => to_unsigned(872, 10), 1391 => to_unsigned(125, 10), 1392 => to_unsigned(729, 10), 1393 => to_unsigned(790, 10), 1394 => to_unsigned(27, 10), 1395 => to_unsigned(545, 10), 1396 => to_unsigned(23, 10), 1397 => to_unsigned(695, 10), 1398 => to_unsigned(118, 10), 1399 => to_unsigned(676, 10), 1400 => to_unsigned(498, 10), 1401 => to_unsigned(283, 10), 1402 => to_unsigned(944, 10), 1403 => to_unsigned(154, 10), 1404 => to_unsigned(873, 10), 1405 => to_unsigned(994, 10), 1406 => to_unsigned(831, 10), 1407 => to_unsigned(44, 10), 1408 => to_unsigned(489, 10), 1409 => to_unsigned(834, 10), 1410 => to_unsigned(405, 10), 1411 => to_unsigned(257, 10), 1412 => to_unsigned(516, 10), 1413 => to_unsigned(485, 10), 1414 => to_unsigned(332, 10), 1415 => to_unsigned(571, 10), 1416 => to_unsigned(409, 10), 1417 => to_unsigned(826, 10), 1418 => to_unsigned(708, 10), 1419 => to_unsigned(747, 10), 1420 => to_unsigned(927, 10), 1421 => to_unsigned(0, 10), 1422 => to_unsigned(69, 10), 1423 => to_unsigned(570, 10), 1424 => to_unsigned(89, 10), 1425 => to_unsigned(160, 10), 1426 => to_unsigned(396, 10), 1427 => to_unsigned(1011, 10), 1428 => to_unsigned(444, 10), 1429 => to_unsigned(100, 10), 1430 => to_unsigned(52, 10), 1431 => to_unsigned(447, 10), 1432 => to_unsigned(539, 10), 1433 => to_unsigned(733, 10), 1434 => to_unsigned(558, 10), 1435 => to_unsigned(172, 10), 1436 => to_unsigned(399, 10), 1437 => to_unsigned(843, 10), 1438 => to_unsigned(365, 10), 1439 => to_unsigned(102, 10), 1440 => to_unsigned(487, 10), 1441 => to_unsigned(932, 10), 1442 => to_unsigned(58, 10), 1443 => to_unsigned(400, 10), 1444 => to_unsigned(130, 10), 1445 => to_unsigned(383, 10), 1446 => to_unsigned(62, 10), 1447 => to_unsigned(328, 10), 1448 => to_unsigned(330, 10), 1449 => to_unsigned(591, 10), 1450 => to_unsigned(812, 10), 1451 => to_unsigned(607, 10), 1452 => to_unsigned(436, 10), 1453 => to_unsigned(1013, 10), 1454 => to_unsigned(611, 10), 1455 => to_unsigned(708, 10), 1456 => to_unsigned(248, 10), 1457 => to_unsigned(534, 10), 1458 => to_unsigned(114, 10), 1459 => to_unsigned(696, 10), 1460 => to_unsigned(616, 10), 1461 => to_unsigned(246, 10), 1462 => to_unsigned(25, 10), 1463 => to_unsigned(592, 10), 1464 => to_unsigned(451, 10), 1465 => to_unsigned(732, 10), 1466 => to_unsigned(923, 10), 1467 => to_unsigned(415, 10), 1468 => to_unsigned(145, 10), 1469 => to_unsigned(513, 10), 1470 => to_unsigned(726, 10), 1471 => to_unsigned(735, 10), 1472 => to_unsigned(809, 10), 1473 => to_unsigned(173, 10), 1474 => to_unsigned(1004, 10), 1475 => to_unsigned(167, 10), 1476 => to_unsigned(991, 10), 1477 => to_unsigned(951, 10), 1478 => to_unsigned(985, 10), 1479 => to_unsigned(344, 10), 1480 => to_unsigned(413, 10), 1481 => to_unsigned(141, 10), 1482 => to_unsigned(242, 10), 1483 => to_unsigned(374, 10), 1484 => to_unsigned(560, 10), 1485 => to_unsigned(706, 10), 1486 => to_unsigned(532, 10), 1487 => to_unsigned(929, 10), 1488 => to_unsigned(176, 10), 1489 => to_unsigned(683, 10), 1490 => to_unsigned(774, 10), 1491 => to_unsigned(684, 10), 1492 => to_unsigned(844, 10), 1493 => to_unsigned(128, 10), 1494 => to_unsigned(410, 10), 1495 => to_unsigned(664, 10), 1496 => to_unsigned(868, 10), 1497 => to_unsigned(452, 10), 1498 => to_unsigned(181, 10), 1499 => to_unsigned(651, 10), 1500 => to_unsigned(641, 10), 1501 => to_unsigned(642, 10), 1502 => to_unsigned(707, 10), 1503 => to_unsigned(642, 10), 1504 => to_unsigned(421, 10), 1505 => to_unsigned(593, 10), 1506 => to_unsigned(284, 10), 1507 => to_unsigned(158, 10), 1508 => to_unsigned(152, 10), 1509 => to_unsigned(833, 10), 1510 => to_unsigned(195, 10), 1511 => to_unsigned(614, 10), 1512 => to_unsigned(978, 10), 1513 => to_unsigned(230, 10), 1514 => to_unsigned(289, 10), 1515 => to_unsigned(719, 10), 1516 => to_unsigned(90, 10), 1517 => to_unsigned(904, 10), 1518 => to_unsigned(65, 10), 1519 => to_unsigned(792, 10), 1520 => to_unsigned(199, 10), 1521 => to_unsigned(630, 10), 1522 => to_unsigned(846, 10), 1523 => to_unsigned(422, 10), 1524 => to_unsigned(491, 10), 1525 => to_unsigned(938, 10), 1526 => to_unsigned(255, 10), 1527 => to_unsigned(694, 10), 1528 => to_unsigned(499, 10), 1529 => to_unsigned(135, 10), 1530 => to_unsigned(457, 10), 1531 => to_unsigned(369, 10), 1532 => to_unsigned(7, 10), 1533 => to_unsigned(450, 10), 1534 => to_unsigned(1012, 10), 1535 => to_unsigned(579, 10), 1536 => to_unsigned(133, 10), 1537 => to_unsigned(7, 10), 1538 => to_unsigned(70, 10), 1539 => to_unsigned(911, 10), 1540 => to_unsigned(934, 10), 1541 => to_unsigned(46, 10), 1542 => to_unsigned(192, 10), 1543 => to_unsigned(663, 10), 1544 => to_unsigned(593, 10), 1545 => to_unsigned(363, 10), 1546 => to_unsigned(912, 10), 1547 => to_unsigned(231, 10), 1548 => to_unsigned(1015, 10), 1549 => to_unsigned(890, 10), 1550 => to_unsigned(1017, 10), 1551 => to_unsigned(508, 10), 1552 => to_unsigned(232, 10), 1553 => to_unsigned(605, 10), 1554 => to_unsigned(78, 10), 1555 => to_unsigned(1003, 10), 1556 => to_unsigned(194, 10), 1557 => to_unsigned(831, 10), 1558 => to_unsigned(263, 10), 1559 => to_unsigned(503, 10), 1560 => to_unsigned(528, 10), 1561 => to_unsigned(1008, 10), 1562 => to_unsigned(132, 10), 1563 => to_unsigned(525, 10), 1564 => to_unsigned(169, 10), 1565 => to_unsigned(502, 10), 1566 => to_unsigned(601, 10), 1567 => to_unsigned(776, 10), 1568 => to_unsigned(474, 10), 1569 => to_unsigned(591, 10), 1570 => to_unsigned(173, 10), 1571 => to_unsigned(47, 10), 1572 => to_unsigned(491, 10), 1573 => to_unsigned(1005, 10), 1574 => to_unsigned(1007, 10), 1575 => to_unsigned(236, 10), 1576 => to_unsigned(713, 10), 1577 => to_unsigned(372, 10), 1578 => to_unsigned(509, 10), 1579 => to_unsigned(188, 10), 1580 => to_unsigned(977, 10), 1581 => to_unsigned(495, 10), 1582 => to_unsigned(994, 10), 1583 => to_unsigned(188, 10), 1584 => to_unsigned(177, 10), 1585 => to_unsigned(997, 10), 1586 => to_unsigned(335, 10), 1587 => to_unsigned(258, 10), 1588 => to_unsigned(751, 10), 1589 => to_unsigned(764, 10), 1590 => to_unsigned(774, 10), 1591 => to_unsigned(523, 10), 1592 => to_unsigned(799, 10), 1593 => to_unsigned(991, 10), 1594 => to_unsigned(597, 10), 1595 => to_unsigned(538, 10), 1596 => to_unsigned(1020, 10), 1597 => to_unsigned(454, 10), 1598 => to_unsigned(580, 10), 1599 => to_unsigned(690, 10), 1600 => to_unsigned(575, 10), 1601 => to_unsigned(338, 10), 1602 => to_unsigned(487, 10), 1603 => to_unsigned(1011, 10), 1604 => to_unsigned(724, 10), 1605 => to_unsigned(823, 10), 1606 => to_unsigned(991, 10), 1607 => to_unsigned(210, 10), 1608 => to_unsigned(426, 10), 1609 => to_unsigned(872, 10), 1610 => to_unsigned(695, 10), 1611 => to_unsigned(276, 10), 1612 => to_unsigned(724, 10), 1613 => to_unsigned(904, 10), 1614 => to_unsigned(934, 10), 1615 => to_unsigned(459, 10), 1616 => to_unsigned(851, 10), 1617 => to_unsigned(665, 10), 1618 => to_unsigned(288, 10), 1619 => to_unsigned(137, 10), 1620 => to_unsigned(1019, 10), 1621 => to_unsigned(168, 10), 1622 => to_unsigned(284, 10), 1623 => to_unsigned(395, 10), 1624 => to_unsigned(482, 10), 1625 => to_unsigned(153, 10), 1626 => to_unsigned(530, 10), 1627 => to_unsigned(756, 10), 1628 => to_unsigned(249, 10), 1629 => to_unsigned(289, 10), 1630 => to_unsigned(753, 10), 1631 => to_unsigned(795, 10), 1632 => to_unsigned(688, 10), 1633 => to_unsigned(258, 10), 1634 => to_unsigned(55, 10), 1635 => to_unsigned(563, 10), 1636 => to_unsigned(101, 10), 1637 => to_unsigned(90, 10), 1638 => to_unsigned(671, 10), 1639 => to_unsigned(719, 10), 1640 => to_unsigned(854, 10), 1641 => to_unsigned(200, 10), 1642 => to_unsigned(142, 10), 1643 => to_unsigned(487, 10), 1644 => to_unsigned(273, 10), 1645 => to_unsigned(306, 10), 1646 => to_unsigned(538, 10), 1647 => to_unsigned(283, 10), 1648 => to_unsigned(961, 10), 1649 => to_unsigned(39, 10), 1650 => to_unsigned(549, 10), 1651 => to_unsigned(979, 10), 1652 => to_unsigned(623, 10), 1653 => to_unsigned(969, 10), 1654 => to_unsigned(245, 10), 1655 => to_unsigned(525, 10), 1656 => to_unsigned(183, 10), 1657 => to_unsigned(228, 10), 1658 => to_unsigned(824, 10), 1659 => to_unsigned(645, 10), 1660 => to_unsigned(459, 10), 1661 => to_unsigned(583, 10), 1662 => to_unsigned(813, 10), 1663 => to_unsigned(957, 10), 1664 => to_unsigned(324, 10), 1665 => to_unsigned(151, 10), 1666 => to_unsigned(494, 10), 1667 => to_unsigned(117, 10), 1668 => to_unsigned(142, 10), 1669 => to_unsigned(546, 10), 1670 => to_unsigned(716, 10), 1671 => to_unsigned(597, 10), 1672 => to_unsigned(981, 10), 1673 => to_unsigned(400, 10), 1674 => to_unsigned(871, 10), 1675 => to_unsigned(225, 10), 1676 => to_unsigned(621, 10), 1677 => to_unsigned(972, 10), 1678 => to_unsigned(60, 10), 1679 => to_unsigned(953, 10), 1680 => to_unsigned(697, 10), 1681 => to_unsigned(820, 10), 1682 => to_unsigned(985, 10), 1683 => to_unsigned(546, 10), 1684 => to_unsigned(248, 10), 1685 => to_unsigned(103, 10), 1686 => to_unsigned(9, 10), 1687 => to_unsigned(730, 10), 1688 => to_unsigned(985, 10), 1689 => to_unsigned(428, 10), 1690 => to_unsigned(357, 10), 1691 => to_unsigned(952, 10), 1692 => to_unsigned(685, 10), 1693 => to_unsigned(523, 10), 1694 => to_unsigned(303, 10), 1695 => to_unsigned(328, 10), 1696 => to_unsigned(144, 10), 1697 => to_unsigned(445, 10), 1698 => to_unsigned(267, 10), 1699 => to_unsigned(406, 10), 1700 => to_unsigned(866, 10), 1701 => to_unsigned(966, 10), 1702 => to_unsigned(45, 10), 1703 => to_unsigned(274, 10), 1704 => to_unsigned(506, 10), 1705 => to_unsigned(664, 10), 1706 => to_unsigned(554, 10), 1707 => to_unsigned(563, 10), 1708 => to_unsigned(154, 10), 1709 => to_unsigned(858, 10), 1710 => to_unsigned(189, 10), 1711 => to_unsigned(109, 10), 1712 => to_unsigned(604, 10), 1713 => to_unsigned(178, 10), 1714 => to_unsigned(619, 10), 1715 => to_unsigned(12, 10), 1716 => to_unsigned(676, 10), 1717 => to_unsigned(420, 10), 1718 => to_unsigned(647, 10), 1719 => to_unsigned(439, 10), 1720 => to_unsigned(157, 10), 1721 => to_unsigned(731, 10), 1722 => to_unsigned(48, 10), 1723 => to_unsigned(638, 10), 1724 => to_unsigned(59, 10), 1725 => to_unsigned(566, 10), 1726 => to_unsigned(813, 10), 1727 => to_unsigned(980, 10), 1728 => to_unsigned(624, 10), 1729 => to_unsigned(209, 10), 1730 => to_unsigned(215, 10), 1731 => to_unsigned(553, 10), 1732 => to_unsigned(467, 10), 1733 => to_unsigned(49, 10), 1734 => to_unsigned(335, 10), 1735 => to_unsigned(934, 10), 1736 => to_unsigned(794, 10), 1737 => to_unsigned(610, 10), 1738 => to_unsigned(473, 10), 1739 => to_unsigned(397, 10), 1740 => to_unsigned(376, 10), 1741 => to_unsigned(366, 10), 1742 => to_unsigned(710, 10), 1743 => to_unsigned(959, 10), 1744 => to_unsigned(24, 10), 1745 => to_unsigned(802, 10), 1746 => to_unsigned(575, 10), 1747 => to_unsigned(398, 10), 1748 => to_unsigned(170, 10), 1749 => to_unsigned(336, 10), 1750 => to_unsigned(985, 10), 1751 => to_unsigned(221, 10), 1752 => to_unsigned(163, 10), 1753 => to_unsigned(418, 10), 1754 => to_unsigned(397, 10), 1755 => to_unsigned(233, 10), 1756 => to_unsigned(225, 10), 1757 => to_unsigned(947, 10), 1758 => to_unsigned(8, 10), 1759 => to_unsigned(92, 10), 1760 => to_unsigned(275, 10), 1761 => to_unsigned(30, 10), 1762 => to_unsigned(450, 10), 1763 => to_unsigned(739, 10), 1764 => to_unsigned(898, 10), 1765 => to_unsigned(938, 10), 1766 => to_unsigned(53, 10), 1767 => to_unsigned(882, 10), 1768 => to_unsigned(461, 10), 1769 => to_unsigned(793, 10), 1770 => to_unsigned(903, 10), 1771 => to_unsigned(742, 10), 1772 => to_unsigned(952, 10), 1773 => to_unsigned(756, 10), 1774 => to_unsigned(861, 10), 1775 => to_unsigned(272, 10), 1776 => to_unsigned(833, 10), 1777 => to_unsigned(439, 10), 1778 => to_unsigned(721, 10), 1779 => to_unsigned(385, 10), 1780 => to_unsigned(737, 10), 1781 => to_unsigned(286, 10), 1782 => to_unsigned(773, 10), 1783 => to_unsigned(565, 10), 1784 => to_unsigned(272, 10), 1785 => to_unsigned(899, 10), 1786 => to_unsigned(467, 10), 1787 => to_unsigned(879, 10), 1788 => to_unsigned(242, 10), 1789 => to_unsigned(500, 10), 1790 => to_unsigned(892, 10), 1791 => to_unsigned(1011, 10), 1792 => to_unsigned(587, 10), 1793 => to_unsigned(749, 10), 1794 => to_unsigned(74, 10), 1795 => to_unsigned(966, 10), 1796 => to_unsigned(747, 10), 1797 => to_unsigned(411, 10), 1798 => to_unsigned(389, 10), 1799 => to_unsigned(195, 10), 1800 => to_unsigned(437, 10), 1801 => to_unsigned(19, 10), 1802 => to_unsigned(548, 10), 1803 => to_unsigned(516, 10), 1804 => to_unsigned(755, 10), 1805 => to_unsigned(411, 10), 1806 => to_unsigned(198, 10), 1807 => to_unsigned(758, 10), 1808 => to_unsigned(231, 10), 1809 => to_unsigned(383, 10), 1810 => to_unsigned(757, 10), 1811 => to_unsigned(715, 10), 1812 => to_unsigned(451, 10), 1813 => to_unsigned(978, 10), 1814 => to_unsigned(666, 10), 1815 => to_unsigned(267, 10), 1816 => to_unsigned(398, 10), 1817 => to_unsigned(85, 10), 1818 => to_unsigned(487, 10), 1819 => to_unsigned(771, 10), 1820 => to_unsigned(861, 10), 1821 => to_unsigned(133, 10), 1822 => to_unsigned(149, 10), 1823 => to_unsigned(864, 10), 1824 => to_unsigned(792, 10), 1825 => to_unsigned(651, 10), 1826 => to_unsigned(31, 10), 1827 => to_unsigned(399, 10), 1828 => to_unsigned(122, 10), 1829 => to_unsigned(712, 10), 1830 => to_unsigned(690, 10), 1831 => to_unsigned(363, 10), 1832 => to_unsigned(773, 10), 1833 => to_unsigned(398, 10), 1834 => to_unsigned(26, 10), 1835 => to_unsigned(472, 10), 1836 => to_unsigned(677, 10), 1837 => to_unsigned(370, 10), 1838 => to_unsigned(762, 10), 1839 => to_unsigned(920, 10), 1840 => to_unsigned(413, 10), 1841 => to_unsigned(823, 10), 1842 => to_unsigned(147, 10), 1843 => to_unsigned(161, 10), 1844 => to_unsigned(710, 10), 1845 => to_unsigned(841, 10), 1846 => to_unsigned(93, 10), 1847 => to_unsigned(106, 10), 1848 => to_unsigned(165, 10), 1849 => to_unsigned(187, 10), 1850 => to_unsigned(789, 10), 1851 => to_unsigned(943, 10), 1852 => to_unsigned(908, 10), 1853 => to_unsigned(444, 10), 1854 => to_unsigned(757, 10), 1855 => to_unsigned(349, 10), 1856 => to_unsigned(532, 10), 1857 => to_unsigned(586, 10), 1858 => to_unsigned(1012, 10), 1859 => to_unsigned(717, 10), 1860 => to_unsigned(639, 10), 1861 => to_unsigned(452, 10), 1862 => to_unsigned(747, 10), 1863 => to_unsigned(674, 10), 1864 => to_unsigned(1006, 10), 1865 => to_unsigned(50, 10), 1866 => to_unsigned(783, 10), 1867 => to_unsigned(956, 10), 1868 => to_unsigned(805, 10), 1869 => to_unsigned(692, 10), 1870 => to_unsigned(892, 10), 1871 => to_unsigned(901, 10), 1872 => to_unsigned(389, 10), 1873 => to_unsigned(975, 10), 1874 => to_unsigned(345, 10), 1875 => to_unsigned(434, 10), 1876 => to_unsigned(573, 10), 1877 => to_unsigned(856, 10), 1878 => to_unsigned(449, 10), 1879 => to_unsigned(195, 10), 1880 => to_unsigned(209, 10), 1881 => to_unsigned(608, 10), 1882 => to_unsigned(310, 10), 1883 => to_unsigned(925, 10), 1884 => to_unsigned(781, 10), 1885 => to_unsigned(679, 10), 1886 => to_unsigned(407, 10), 1887 => to_unsigned(356, 10), 1888 => to_unsigned(792, 10), 1889 => to_unsigned(170, 10), 1890 => to_unsigned(820, 10), 1891 => to_unsigned(135, 10), 1892 => to_unsigned(651, 10), 1893 => to_unsigned(252, 10), 1894 => to_unsigned(746, 10), 1895 => to_unsigned(914, 10), 1896 => to_unsigned(722, 10), 1897 => to_unsigned(287, 10), 1898 => to_unsigned(51, 10), 1899 => to_unsigned(550, 10), 1900 => to_unsigned(122, 10), 1901 => to_unsigned(419, 10), 1902 => to_unsigned(618, 10), 1903 => to_unsigned(734, 10), 1904 => to_unsigned(710, 10), 1905 => to_unsigned(491, 10), 1906 => to_unsigned(618, 10), 1907 => to_unsigned(436, 10), 1908 => to_unsigned(167, 10), 1909 => to_unsigned(92, 10), 1910 => to_unsigned(388, 10), 1911 => to_unsigned(985, 10), 1912 => to_unsigned(125, 10), 1913 => to_unsigned(666, 10), 1914 => to_unsigned(614, 10), 1915 => to_unsigned(652, 10), 1916 => to_unsigned(604, 10), 1917 => to_unsigned(528, 10), 1918 => to_unsigned(691, 10), 1919 => to_unsigned(935, 10), 1920 => to_unsigned(724, 10), 1921 => to_unsigned(186, 10), 1922 => to_unsigned(137, 10), 1923 => to_unsigned(1012, 10), 1924 => to_unsigned(831, 10), 1925 => to_unsigned(687, 10), 1926 => to_unsigned(727, 10), 1927 => to_unsigned(677, 10), 1928 => to_unsigned(711, 10), 1929 => to_unsigned(798, 10), 1930 => to_unsigned(781, 10), 1931 => to_unsigned(312, 10), 1932 => to_unsigned(130, 10), 1933 => to_unsigned(480, 10), 1934 => to_unsigned(180, 10), 1935 => to_unsigned(662, 10), 1936 => to_unsigned(734, 10), 1937 => to_unsigned(920, 10), 1938 => to_unsigned(94, 10), 1939 => to_unsigned(282, 10), 1940 => to_unsigned(313, 10), 1941 => to_unsigned(494, 10), 1942 => to_unsigned(232, 10), 1943 => to_unsigned(909, 10), 1944 => to_unsigned(198, 10), 1945 => to_unsigned(229, 10), 1946 => to_unsigned(195, 10), 1947 => to_unsigned(912, 10), 1948 => to_unsigned(525, 10), 1949 => to_unsigned(650, 10), 1950 => to_unsigned(208, 10), 1951 => to_unsigned(497, 10), 1952 => to_unsigned(917, 10), 1953 => to_unsigned(340, 10), 1954 => to_unsigned(208, 10), 1955 => to_unsigned(620, 10), 1956 => to_unsigned(548, 10), 1957 => to_unsigned(756, 10), 1958 => to_unsigned(51, 10), 1959 => to_unsigned(1010, 10), 1960 => to_unsigned(305, 10), 1961 => to_unsigned(528, 10), 1962 => to_unsigned(418, 10), 1963 => to_unsigned(489, 10), 1964 => to_unsigned(199, 10), 1965 => to_unsigned(479, 10), 1966 => to_unsigned(374, 10), 1967 => to_unsigned(362, 10), 1968 => to_unsigned(893, 10), 1969 => to_unsigned(423, 10), 1970 => to_unsigned(10, 10), 1971 => to_unsigned(594, 10), 1972 => to_unsigned(892, 10), 1973 => to_unsigned(539, 10), 1974 => to_unsigned(359, 10), 1975 => to_unsigned(256, 10), 1976 => to_unsigned(180, 10), 1977 => to_unsigned(841, 10), 1978 => to_unsigned(338, 10), 1979 => to_unsigned(901, 10), 1980 => to_unsigned(980, 10), 1981 => to_unsigned(651, 10), 1982 => to_unsigned(384, 10), 1983 => to_unsigned(777, 10), 1984 => to_unsigned(297, 10), 1985 => to_unsigned(520, 10), 1986 => to_unsigned(372, 10), 1987 => to_unsigned(197, 10), 1988 => to_unsigned(510, 10), 1989 => to_unsigned(25, 10), 1990 => to_unsigned(491, 10), 1991 => to_unsigned(549, 10), 1992 => to_unsigned(860, 10), 1993 => to_unsigned(446, 10), 1994 => to_unsigned(849, 10), 1995 => to_unsigned(172, 10), 1996 => to_unsigned(777, 10), 1997 => to_unsigned(975, 10), 1998 => to_unsigned(838, 10), 1999 => to_unsigned(315, 10), 2000 => to_unsigned(754, 10), 2001 => to_unsigned(394, 10), 2002 => to_unsigned(139, 10), 2003 => to_unsigned(262, 10), 2004 => to_unsigned(915, 10), 2005 => to_unsigned(863, 10), 2006 => to_unsigned(855, 10), 2007 => to_unsigned(131, 10), 2008 => to_unsigned(747, 10), 2009 => to_unsigned(366, 10), 2010 => to_unsigned(878, 10), 2011 => to_unsigned(375, 10), 2012 => to_unsigned(50, 10), 2013 => to_unsigned(389, 10), 2014 => to_unsigned(930, 10), 2015 => to_unsigned(246, 10), 2016 => to_unsigned(503, 10), 2017 => to_unsigned(235, 10), 2018 => to_unsigned(92, 10), 2019 => to_unsigned(784, 10), 2020 => to_unsigned(373, 10), 2021 => to_unsigned(44, 10), 2022 => to_unsigned(263, 10), 2023 => to_unsigned(100, 10), 2024 => to_unsigned(590, 10), 2025 => to_unsigned(177, 10), 2026 => to_unsigned(5, 10), 2027 => to_unsigned(726, 10), 2028 => to_unsigned(24, 10), 2029 => to_unsigned(949, 10), 2030 => to_unsigned(99, 10), 2031 => to_unsigned(141, 10), 2032 => to_unsigned(227, 10), 2033 => to_unsigned(518, 10), 2034 => to_unsigned(904, 10), 2035 => to_unsigned(643, 10), 2036 => to_unsigned(828, 10), 2037 => to_unsigned(637, 10), 2038 => to_unsigned(806, 10), 2039 => to_unsigned(686, 10), 2040 => to_unsigned(365, 10), 2041 => to_unsigned(129, 10), 2042 => to_unsigned(918, 10), 2043 => to_unsigned(433, 10), 2044 => to_unsigned(674, 10), 2045 => to_unsigned(141, 10), 2046 => to_unsigned(335, 10), 2047 => to_unsigned(435, 10)),
            7 => (0 => to_unsigned(341, 10), 1 => to_unsigned(15, 10), 2 => to_unsigned(773, 10), 3 => to_unsigned(317, 10), 4 => to_unsigned(28, 10), 5 => to_unsigned(470, 10), 6 => to_unsigned(515, 10), 7 => to_unsigned(614, 10), 8 => to_unsigned(624, 10), 9 => to_unsigned(181, 10), 10 => to_unsigned(720, 10), 11 => to_unsigned(947, 10), 12 => to_unsigned(826, 10), 13 => to_unsigned(384, 10), 14 => to_unsigned(10, 10), 15 => to_unsigned(885, 10), 16 => to_unsigned(983, 10), 17 => to_unsigned(158, 10), 18 => to_unsigned(850, 10), 19 => to_unsigned(5, 10), 20 => to_unsigned(436, 10), 21 => to_unsigned(520, 10), 22 => to_unsigned(14, 10), 23 => to_unsigned(284, 10), 24 => to_unsigned(654, 10), 25 => to_unsigned(441, 10), 26 => to_unsigned(660, 10), 27 => to_unsigned(909, 10), 28 => to_unsigned(910, 10), 29 => to_unsigned(965, 10), 30 => to_unsigned(609, 10), 31 => to_unsigned(423, 10), 32 => to_unsigned(369, 10), 33 => to_unsigned(533, 10), 34 => to_unsigned(35, 10), 35 => to_unsigned(22, 10), 36 => to_unsigned(481, 10), 37 => to_unsigned(1008, 10), 38 => to_unsigned(679, 10), 39 => to_unsigned(233, 10), 40 => to_unsigned(250, 10), 41 => to_unsigned(128, 10), 42 => to_unsigned(623, 10), 43 => to_unsigned(419, 10), 44 => to_unsigned(257, 10), 45 => to_unsigned(977, 10), 46 => to_unsigned(646, 10), 47 => to_unsigned(817, 10), 48 => to_unsigned(370, 10), 49 => to_unsigned(710, 10), 50 => to_unsigned(418, 10), 51 => to_unsigned(274, 10), 52 => to_unsigned(420, 10), 53 => to_unsigned(336, 10), 54 => to_unsigned(669, 10), 55 => to_unsigned(648, 10), 56 => to_unsigned(1000, 10), 57 => to_unsigned(811, 10), 58 => to_unsigned(928, 10), 59 => to_unsigned(930, 10), 60 => to_unsigned(913, 10), 61 => to_unsigned(443, 10), 62 => to_unsigned(381, 10), 63 => to_unsigned(624, 10), 64 => to_unsigned(69, 10), 65 => to_unsigned(265, 10), 66 => to_unsigned(522, 10), 67 => to_unsigned(556, 10), 68 => to_unsigned(489, 10), 69 => to_unsigned(489, 10), 70 => to_unsigned(976, 10), 71 => to_unsigned(499, 10), 72 => to_unsigned(472, 10), 73 => to_unsigned(24, 10), 74 => to_unsigned(598, 10), 75 => to_unsigned(836, 10), 76 => to_unsigned(262, 10), 77 => to_unsigned(916, 10), 78 => to_unsigned(832, 10), 79 => to_unsigned(816, 10), 80 => to_unsigned(750, 10), 81 => to_unsigned(438, 10), 82 => to_unsigned(459, 10), 83 => to_unsigned(359, 10), 84 => to_unsigned(141, 10), 85 => to_unsigned(479, 10), 86 => to_unsigned(273, 10), 87 => to_unsigned(711, 10), 88 => to_unsigned(575, 10), 89 => to_unsigned(59, 10), 90 => to_unsigned(330, 10), 91 => to_unsigned(956, 10), 92 => to_unsigned(1007, 10), 93 => to_unsigned(514, 10), 94 => to_unsigned(98, 10), 95 => to_unsigned(467, 10), 96 => to_unsigned(526, 10), 97 => to_unsigned(82, 10), 98 => to_unsigned(797, 10), 99 => to_unsigned(703, 10), 100 => to_unsigned(253, 10), 101 => to_unsigned(160, 10), 102 => to_unsigned(586, 10), 103 => to_unsigned(472, 10), 104 => to_unsigned(165, 10), 105 => to_unsigned(856, 10), 106 => to_unsigned(818, 10), 107 => to_unsigned(932, 10), 108 => to_unsigned(598, 10), 109 => to_unsigned(629, 10), 110 => to_unsigned(918, 10), 111 => to_unsigned(273, 10), 112 => to_unsigned(113, 10), 113 => to_unsigned(81, 10), 114 => to_unsigned(59, 10), 115 => to_unsigned(522, 10), 116 => to_unsigned(794, 10), 117 => to_unsigned(412, 10), 118 => to_unsigned(15, 10), 119 => to_unsigned(946, 10), 120 => to_unsigned(586, 10), 121 => to_unsigned(912, 10), 122 => to_unsigned(244, 10), 123 => to_unsigned(704, 10), 124 => to_unsigned(726, 10), 125 => to_unsigned(558, 10), 126 => to_unsigned(479, 10), 127 => to_unsigned(286, 10), 128 => to_unsigned(942, 10), 129 => to_unsigned(775, 10), 130 => to_unsigned(510, 10), 131 => to_unsigned(464, 10), 132 => to_unsigned(919, 10), 133 => to_unsigned(842, 10), 134 => to_unsigned(889, 10), 135 => to_unsigned(64, 10), 136 => to_unsigned(127, 10), 137 => to_unsigned(615, 10), 138 => to_unsigned(3, 10), 139 => to_unsigned(614, 10), 140 => to_unsigned(6, 10), 141 => to_unsigned(776, 10), 142 => to_unsigned(449, 10), 143 => to_unsigned(214, 10), 144 => to_unsigned(704, 10), 145 => to_unsigned(135, 10), 146 => to_unsigned(807, 10), 147 => to_unsigned(653, 10), 148 => to_unsigned(284, 10), 149 => to_unsigned(105, 10), 150 => to_unsigned(382, 10), 151 => to_unsigned(593, 10), 152 => to_unsigned(94, 10), 153 => to_unsigned(387, 10), 154 => to_unsigned(322, 10), 155 => to_unsigned(275, 10), 156 => to_unsigned(196, 10), 157 => to_unsigned(611, 10), 158 => to_unsigned(428, 10), 159 => to_unsigned(201, 10), 160 => to_unsigned(279, 10), 161 => to_unsigned(735, 10), 162 => to_unsigned(2, 10), 163 => to_unsigned(971, 10), 164 => to_unsigned(66, 10), 165 => to_unsigned(662, 10), 166 => to_unsigned(193, 10), 167 => to_unsigned(453, 10), 168 => to_unsigned(565, 10), 169 => to_unsigned(410, 10), 170 => to_unsigned(936, 10), 171 => to_unsigned(390, 10), 172 => to_unsigned(653, 10), 173 => to_unsigned(948, 10), 174 => to_unsigned(181, 10), 175 => to_unsigned(365, 10), 176 => to_unsigned(261, 10), 177 => to_unsigned(698, 10), 178 => to_unsigned(422, 10), 179 => to_unsigned(841, 10), 180 => to_unsigned(581, 10), 181 => to_unsigned(470, 10), 182 => to_unsigned(666, 10), 183 => to_unsigned(558, 10), 184 => to_unsigned(903, 10), 185 => to_unsigned(798, 10), 186 => to_unsigned(358, 10), 187 => to_unsigned(887, 10), 188 => to_unsigned(390, 10), 189 => to_unsigned(679, 10), 190 => to_unsigned(532, 10), 191 => to_unsigned(498, 10), 192 => to_unsigned(560, 10), 193 => to_unsigned(986, 10), 194 => to_unsigned(65, 10), 195 => to_unsigned(420, 10), 196 => to_unsigned(900, 10), 197 => to_unsigned(669, 10), 198 => to_unsigned(507, 10), 199 => to_unsigned(471, 10), 200 => to_unsigned(225, 10), 201 => to_unsigned(351, 10), 202 => to_unsigned(210, 10), 203 => to_unsigned(787, 10), 204 => to_unsigned(771, 10), 205 => to_unsigned(433, 10), 206 => to_unsigned(323, 10), 207 => to_unsigned(12, 10), 208 => to_unsigned(937, 10), 209 => to_unsigned(971, 10), 210 => to_unsigned(32, 10), 211 => to_unsigned(947, 10), 212 => to_unsigned(21, 10), 213 => to_unsigned(224, 10), 214 => to_unsigned(648, 10), 215 => to_unsigned(351, 10), 216 => to_unsigned(92, 10), 217 => to_unsigned(832, 10), 218 => to_unsigned(900, 10), 219 => to_unsigned(923, 10), 220 => to_unsigned(814, 10), 221 => to_unsigned(267, 10), 222 => to_unsigned(985, 10), 223 => to_unsigned(723, 10), 224 => to_unsigned(520, 10), 225 => to_unsigned(104, 10), 226 => to_unsigned(387, 10), 227 => to_unsigned(468, 10), 228 => to_unsigned(9, 10), 229 => to_unsigned(598, 10), 230 => to_unsigned(547, 10), 231 => to_unsigned(901, 10), 232 => to_unsigned(469, 10), 233 => to_unsigned(992, 10), 234 => to_unsigned(60, 10), 235 => to_unsigned(787, 10), 236 => to_unsigned(218, 10), 237 => to_unsigned(148, 10), 238 => to_unsigned(686, 10), 239 => to_unsigned(596, 10), 240 => to_unsigned(191, 10), 241 => to_unsigned(15, 10), 242 => to_unsigned(344, 10), 243 => to_unsigned(149, 10), 244 => to_unsigned(340, 10), 245 => to_unsigned(358, 10), 246 => to_unsigned(589, 10), 247 => to_unsigned(121, 10), 248 => to_unsigned(78, 10), 249 => to_unsigned(851, 10), 250 => to_unsigned(775, 10), 251 => to_unsigned(921, 10), 252 => to_unsigned(198, 10), 253 => to_unsigned(552, 10), 254 => to_unsigned(337, 10), 255 => to_unsigned(687, 10), 256 => to_unsigned(695, 10), 257 => to_unsigned(378, 10), 258 => to_unsigned(847, 10), 259 => to_unsigned(795, 10), 260 => to_unsigned(593, 10), 261 => to_unsigned(581, 10), 262 => to_unsigned(8, 10), 263 => to_unsigned(464, 10), 264 => to_unsigned(466, 10), 265 => to_unsigned(39, 10), 266 => to_unsigned(579, 10), 267 => to_unsigned(776, 10), 268 => to_unsigned(910, 10), 269 => to_unsigned(508, 10), 270 => to_unsigned(194, 10), 271 => to_unsigned(88, 10), 272 => to_unsigned(557, 10), 273 => to_unsigned(446, 10), 274 => to_unsigned(839, 10), 275 => to_unsigned(639, 10), 276 => to_unsigned(779, 10), 277 => to_unsigned(740, 10), 278 => to_unsigned(853, 10), 279 => to_unsigned(678, 10), 280 => to_unsigned(488, 10), 281 => to_unsigned(516, 10), 282 => to_unsigned(680, 10), 283 => to_unsigned(877, 10), 284 => to_unsigned(486, 10), 285 => to_unsigned(564, 10), 286 => to_unsigned(39, 10), 287 => to_unsigned(419, 10), 288 => to_unsigned(146, 10), 289 => to_unsigned(355, 10), 290 => to_unsigned(684, 10), 291 => to_unsigned(946, 10), 292 => to_unsigned(734, 10), 293 => to_unsigned(342, 10), 294 => to_unsigned(671, 10), 295 => to_unsigned(151, 10), 296 => to_unsigned(900, 10), 297 => to_unsigned(16, 10), 298 => to_unsigned(404, 10), 299 => to_unsigned(622, 10), 300 => to_unsigned(260, 10), 301 => to_unsigned(749, 10), 302 => to_unsigned(462, 10), 303 => to_unsigned(896, 10), 304 => to_unsigned(150, 10), 305 => to_unsigned(821, 10), 306 => to_unsigned(926, 10), 307 => to_unsigned(579, 10), 308 => to_unsigned(970, 10), 309 => to_unsigned(944, 10), 310 => to_unsigned(241, 10), 311 => to_unsigned(469, 10), 312 => to_unsigned(226, 10), 313 => to_unsigned(656, 10), 314 => to_unsigned(55, 10), 315 => to_unsigned(395, 10), 316 => to_unsigned(746, 10), 317 => to_unsigned(648, 10), 318 => to_unsigned(376, 10), 319 => to_unsigned(702, 10), 320 => to_unsigned(983, 10), 321 => to_unsigned(265, 10), 322 => to_unsigned(95, 10), 323 => to_unsigned(850, 10), 324 => to_unsigned(71, 10), 325 => to_unsigned(552, 10), 326 => to_unsigned(900, 10), 327 => to_unsigned(1001, 10), 328 => to_unsigned(580, 10), 329 => to_unsigned(895, 10), 330 => to_unsigned(131, 10), 331 => to_unsigned(133, 10), 332 => to_unsigned(427, 10), 333 => to_unsigned(984, 10), 334 => to_unsigned(340, 10), 335 => to_unsigned(474, 10), 336 => to_unsigned(276, 10), 337 => to_unsigned(81, 10), 338 => to_unsigned(453, 10), 339 => to_unsigned(711, 10), 340 => to_unsigned(900, 10), 341 => to_unsigned(740, 10), 342 => to_unsigned(930, 10), 343 => to_unsigned(1014, 10), 344 => to_unsigned(741, 10), 345 => to_unsigned(612, 10), 346 => to_unsigned(513, 10), 347 => to_unsigned(769, 10), 348 => to_unsigned(1014, 10), 349 => to_unsigned(935, 10), 350 => to_unsigned(627, 10), 351 => to_unsigned(436, 10), 352 => to_unsigned(338, 10), 353 => to_unsigned(499, 10), 354 => to_unsigned(120, 10), 355 => to_unsigned(84, 10), 356 => to_unsigned(86, 10), 357 => to_unsigned(797, 10), 358 => to_unsigned(714, 10), 359 => to_unsigned(531, 10), 360 => to_unsigned(295, 10), 361 => to_unsigned(708, 10), 362 => to_unsigned(168, 10), 363 => to_unsigned(446, 10), 364 => to_unsigned(856, 10), 365 => to_unsigned(912, 10), 366 => to_unsigned(1002, 10), 367 => to_unsigned(203, 10), 368 => to_unsigned(784, 10), 369 => to_unsigned(922, 10), 370 => to_unsigned(290, 10), 371 => to_unsigned(741, 10), 372 => to_unsigned(734, 10), 373 => to_unsigned(152, 10), 374 => to_unsigned(894, 10), 375 => to_unsigned(17, 10), 376 => to_unsigned(383, 10), 377 => to_unsigned(533, 10), 378 => to_unsigned(288, 10), 379 => to_unsigned(723, 10), 380 => to_unsigned(769, 10), 381 => to_unsigned(402, 10), 382 => to_unsigned(621, 10), 383 => to_unsigned(189, 10), 384 => to_unsigned(948, 10), 385 => to_unsigned(322, 10), 386 => to_unsigned(812, 10), 387 => to_unsigned(125, 10), 388 => to_unsigned(899, 10), 389 => to_unsigned(400, 10), 390 => to_unsigned(681, 10), 391 => to_unsigned(55, 10), 392 => to_unsigned(996, 10), 393 => to_unsigned(275, 10), 394 => to_unsigned(45, 10), 395 => to_unsigned(795, 10), 396 => to_unsigned(407, 10), 397 => to_unsigned(92, 10), 398 => to_unsigned(603, 10), 399 => to_unsigned(693, 10), 400 => to_unsigned(268, 10), 401 => to_unsigned(567, 10), 402 => to_unsigned(595, 10), 403 => to_unsigned(773, 10), 404 => to_unsigned(543, 10), 405 => to_unsigned(12, 10), 406 => to_unsigned(769, 10), 407 => to_unsigned(373, 10), 408 => to_unsigned(977, 10), 409 => to_unsigned(954, 10), 410 => to_unsigned(527, 10), 411 => to_unsigned(734, 10), 412 => to_unsigned(545, 10), 413 => to_unsigned(676, 10), 414 => to_unsigned(381, 10), 415 => to_unsigned(266, 10), 416 => to_unsigned(791, 10), 417 => to_unsigned(852, 10), 418 => to_unsigned(338, 10), 419 => to_unsigned(601, 10), 420 => to_unsigned(310, 10), 421 => to_unsigned(281, 10), 422 => to_unsigned(37, 10), 423 => to_unsigned(572, 10), 424 => to_unsigned(752, 10), 425 => to_unsigned(271, 10), 426 => to_unsigned(460, 10), 427 => to_unsigned(27, 10), 428 => to_unsigned(229, 10), 429 => to_unsigned(68, 10), 430 => to_unsigned(1002, 10), 431 => to_unsigned(529, 10), 432 => to_unsigned(1001, 10), 433 => to_unsigned(297, 10), 434 => to_unsigned(79, 10), 435 => to_unsigned(428, 10), 436 => to_unsigned(478, 10), 437 => to_unsigned(1020, 10), 438 => to_unsigned(306, 10), 439 => to_unsigned(478, 10), 440 => to_unsigned(44, 10), 441 => to_unsigned(524, 10), 442 => to_unsigned(207, 10), 443 => to_unsigned(209, 10), 444 => to_unsigned(729, 10), 445 => to_unsigned(477, 10), 446 => to_unsigned(833, 10), 447 => to_unsigned(1001, 10), 448 => to_unsigned(414, 10), 449 => to_unsigned(824, 10), 450 => to_unsigned(489, 10), 451 => to_unsigned(438, 10), 452 => to_unsigned(495, 10), 453 => to_unsigned(201, 10), 454 => to_unsigned(911, 10), 455 => to_unsigned(940, 10), 456 => to_unsigned(328, 10), 457 => to_unsigned(39, 10), 458 => to_unsigned(317, 10), 459 => to_unsigned(525, 10), 460 => to_unsigned(389, 10), 461 => to_unsigned(624, 10), 462 => to_unsigned(355, 10), 463 => to_unsigned(802, 10), 464 => to_unsigned(504, 10), 465 => to_unsigned(425, 10), 466 => to_unsigned(479, 10), 467 => to_unsigned(701, 10), 468 => to_unsigned(237, 10), 469 => to_unsigned(933, 10), 470 => to_unsigned(725, 10), 471 => to_unsigned(374, 10), 472 => to_unsigned(253, 10), 473 => to_unsigned(72, 10), 474 => to_unsigned(501, 10), 475 => to_unsigned(405, 10), 476 => to_unsigned(138, 10), 477 => to_unsigned(869, 10), 478 => to_unsigned(634, 10), 479 => to_unsigned(53, 10), 480 => to_unsigned(67, 10), 481 => to_unsigned(598, 10), 482 => to_unsigned(19, 10), 483 => to_unsigned(527, 10), 484 => to_unsigned(152, 10), 485 => to_unsigned(846, 10), 486 => to_unsigned(864, 10), 487 => to_unsigned(423, 10), 488 => to_unsigned(669, 10), 489 => to_unsigned(436, 10), 490 => to_unsigned(463, 10), 491 => to_unsigned(985, 10), 492 => to_unsigned(516, 10), 493 => to_unsigned(53, 10), 494 => to_unsigned(498, 10), 495 => to_unsigned(314, 10), 496 => to_unsigned(201, 10), 497 => to_unsigned(617, 10), 498 => to_unsigned(725, 10), 499 => to_unsigned(100, 10), 500 => to_unsigned(751, 10), 501 => to_unsigned(392, 10), 502 => to_unsigned(1001, 10), 503 => to_unsigned(551, 10), 504 => to_unsigned(294, 10), 505 => to_unsigned(299, 10), 506 => to_unsigned(614, 10), 507 => to_unsigned(472, 10), 508 => to_unsigned(1019, 10), 509 => to_unsigned(856, 10), 510 => to_unsigned(522, 10), 511 => to_unsigned(180, 10), 512 => to_unsigned(828, 10), 513 => to_unsigned(275, 10), 514 => to_unsigned(873, 10), 515 => to_unsigned(13, 10), 516 => to_unsigned(203, 10), 517 => to_unsigned(660, 10), 518 => to_unsigned(88, 10), 519 => to_unsigned(400, 10), 520 => to_unsigned(616, 10), 521 => to_unsigned(933, 10), 522 => to_unsigned(705, 10), 523 => to_unsigned(1017, 10), 524 => to_unsigned(752, 10), 525 => to_unsigned(219, 10), 526 => to_unsigned(339, 10), 527 => to_unsigned(140, 10), 528 => to_unsigned(835, 10), 529 => to_unsigned(825, 10), 530 => to_unsigned(561, 10), 531 => to_unsigned(726, 10), 532 => to_unsigned(973, 10), 533 => to_unsigned(157, 10), 534 => to_unsigned(1011, 10), 535 => to_unsigned(248, 10), 536 => to_unsigned(549, 10), 537 => to_unsigned(689, 10), 538 => to_unsigned(988, 10), 539 => to_unsigned(954, 10), 540 => to_unsigned(237, 10), 541 => to_unsigned(795, 10), 542 => to_unsigned(131, 10), 543 => to_unsigned(31, 10), 544 => to_unsigned(358, 10), 545 => to_unsigned(968, 10), 546 => to_unsigned(965, 10), 547 => to_unsigned(246, 10), 548 => to_unsigned(335, 10), 549 => to_unsigned(859, 10), 550 => to_unsigned(497, 10), 551 => to_unsigned(614, 10), 552 => to_unsigned(109, 10), 553 => to_unsigned(626, 10), 554 => to_unsigned(224, 10), 555 => to_unsigned(353, 10), 556 => to_unsigned(792, 10), 557 => to_unsigned(480, 10), 558 => to_unsigned(694, 10), 559 => to_unsigned(466, 10), 560 => to_unsigned(232, 10), 561 => to_unsigned(633, 10), 562 => to_unsigned(276, 10), 563 => to_unsigned(948, 10), 564 => to_unsigned(920, 10), 565 => to_unsigned(514, 10), 566 => to_unsigned(802, 10), 567 => to_unsigned(471, 10), 568 => to_unsigned(527, 10), 569 => to_unsigned(282, 10), 570 => to_unsigned(145, 10), 571 => to_unsigned(607, 10), 572 => to_unsigned(468, 10), 573 => to_unsigned(472, 10), 574 => to_unsigned(744, 10), 575 => to_unsigned(793, 10), 576 => to_unsigned(171, 10), 577 => to_unsigned(408, 10), 578 => to_unsigned(634, 10), 579 => to_unsigned(602, 10), 580 => to_unsigned(1020, 10), 581 => to_unsigned(459, 10), 582 => to_unsigned(219, 10), 583 => to_unsigned(412, 10), 584 => to_unsigned(272, 10), 585 => to_unsigned(294, 10), 586 => to_unsigned(59, 10), 587 => to_unsigned(636, 10), 588 => to_unsigned(163, 10), 589 => to_unsigned(300, 10), 590 => to_unsigned(223, 10), 591 => to_unsigned(499, 10), 592 => to_unsigned(679, 10), 593 => to_unsigned(825, 10), 594 => to_unsigned(712, 10), 595 => to_unsigned(74, 10), 596 => to_unsigned(421, 10), 597 => to_unsigned(62, 10), 598 => to_unsigned(75, 10), 599 => to_unsigned(405, 10), 600 => to_unsigned(822, 10), 601 => to_unsigned(898, 10), 602 => to_unsigned(489, 10), 603 => to_unsigned(294, 10), 604 => to_unsigned(259, 10), 605 => to_unsigned(597, 10), 606 => to_unsigned(803, 10), 607 => to_unsigned(227, 10), 608 => to_unsigned(888, 10), 609 => to_unsigned(964, 10), 610 => to_unsigned(566, 10), 611 => to_unsigned(563, 10), 612 => to_unsigned(269, 10), 613 => to_unsigned(68, 10), 614 => to_unsigned(439, 10), 615 => to_unsigned(584, 10), 616 => to_unsigned(116, 10), 617 => to_unsigned(850, 10), 618 => to_unsigned(991, 10), 619 => to_unsigned(206, 10), 620 => to_unsigned(608, 10), 621 => to_unsigned(421, 10), 622 => to_unsigned(581, 10), 623 => to_unsigned(1012, 10), 624 => to_unsigned(617, 10), 625 => to_unsigned(690, 10), 626 => to_unsigned(370, 10), 627 => to_unsigned(947, 10), 628 => to_unsigned(788, 10), 629 => to_unsigned(160, 10), 630 => to_unsigned(252, 10), 631 => to_unsigned(586, 10), 632 => to_unsigned(820, 10), 633 => to_unsigned(175, 10), 634 => to_unsigned(68, 10), 635 => to_unsigned(69, 10), 636 => to_unsigned(412, 10), 637 => to_unsigned(874, 10), 638 => to_unsigned(541, 10), 639 => to_unsigned(645, 10), 640 => to_unsigned(474, 10), 641 => to_unsigned(78, 10), 642 => to_unsigned(950, 10), 643 => to_unsigned(665, 10), 644 => to_unsigned(420, 10), 645 => to_unsigned(10, 10), 646 => to_unsigned(706, 10), 647 => to_unsigned(175, 10), 648 => to_unsigned(382, 10), 649 => to_unsigned(549, 10), 650 => to_unsigned(711, 10), 651 => to_unsigned(397, 10), 652 => to_unsigned(863, 10), 653 => to_unsigned(489, 10), 654 => to_unsigned(797, 10), 655 => to_unsigned(133, 10), 656 => to_unsigned(461, 10), 657 => to_unsigned(347, 10), 658 => to_unsigned(422, 10), 659 => to_unsigned(528, 10), 660 => to_unsigned(798, 10), 661 => to_unsigned(664, 10), 662 => to_unsigned(56, 10), 663 => to_unsigned(209, 10), 664 => to_unsigned(307, 10), 665 => to_unsigned(225, 10), 666 => to_unsigned(336, 10), 667 => to_unsigned(265, 10), 668 => to_unsigned(570, 10), 669 => to_unsigned(822, 10), 670 => to_unsigned(961, 10), 671 => to_unsigned(46, 10), 672 => to_unsigned(363, 10), 673 => to_unsigned(414, 10), 674 => to_unsigned(733, 10), 675 => to_unsigned(658, 10), 676 => to_unsigned(83, 10), 677 => to_unsigned(52, 10), 678 => to_unsigned(305, 10), 679 => to_unsigned(764, 10), 680 => to_unsigned(718, 10), 681 => to_unsigned(250, 10), 682 => to_unsigned(842, 10), 683 => to_unsigned(754, 10), 684 => to_unsigned(973, 10), 685 => to_unsigned(67, 10), 686 => to_unsigned(735, 10), 687 => to_unsigned(198, 10), 688 => to_unsigned(951, 10), 689 => to_unsigned(975, 10), 690 => to_unsigned(976, 10), 691 => to_unsigned(629, 10), 692 => to_unsigned(123, 10), 693 => to_unsigned(34, 10), 694 => to_unsigned(719, 10), 695 => to_unsigned(195, 10), 696 => to_unsigned(950, 10), 697 => to_unsigned(619, 10), 698 => to_unsigned(18, 10), 699 => to_unsigned(286, 10), 700 => to_unsigned(299, 10), 701 => to_unsigned(171, 10), 702 => to_unsigned(915, 10), 703 => to_unsigned(433, 10), 704 => to_unsigned(69, 10), 705 => to_unsigned(369, 10), 706 => to_unsigned(326, 10), 707 => to_unsigned(459, 10), 708 => to_unsigned(259, 10), 709 => to_unsigned(913, 10), 710 => to_unsigned(915, 10), 711 => to_unsigned(838, 10), 712 => to_unsigned(377, 10), 713 => to_unsigned(153, 10), 714 => to_unsigned(757, 10), 715 => to_unsigned(600, 10), 716 => to_unsigned(66, 10), 717 => to_unsigned(150, 10), 718 => to_unsigned(246, 10), 719 => to_unsigned(849, 10), 720 => to_unsigned(751, 10), 721 => to_unsigned(758, 10), 722 => to_unsigned(278, 10), 723 => to_unsigned(398, 10), 724 => to_unsigned(612, 10), 725 => to_unsigned(274, 10), 726 => to_unsigned(850, 10), 727 => to_unsigned(495, 10), 728 => to_unsigned(725, 10), 729 => to_unsigned(914, 10), 730 => to_unsigned(591, 10), 731 => to_unsigned(278, 10), 732 => to_unsigned(375, 10), 733 => to_unsigned(398, 10), 734 => to_unsigned(966, 10), 735 => to_unsigned(500, 10), 736 => to_unsigned(148, 10), 737 => to_unsigned(332, 10), 738 => to_unsigned(38, 10), 739 => to_unsigned(22, 10), 740 => to_unsigned(554, 10), 741 => to_unsigned(67, 10), 742 => to_unsigned(183, 10), 743 => to_unsigned(281, 10), 744 => to_unsigned(546, 10), 745 => to_unsigned(926, 10), 746 => to_unsigned(962, 10), 747 => to_unsigned(619, 10), 748 => to_unsigned(657, 10), 749 => to_unsigned(884, 10), 750 => to_unsigned(285, 10), 751 => to_unsigned(24, 10), 752 => to_unsigned(369, 10), 753 => to_unsigned(107, 10), 754 => to_unsigned(980, 10), 755 => to_unsigned(828, 10), 756 => to_unsigned(915, 10), 757 => to_unsigned(818, 10), 758 => to_unsigned(814, 10), 759 => to_unsigned(205, 10), 760 => to_unsigned(431, 10), 761 => to_unsigned(692, 10), 762 => to_unsigned(374, 10), 763 => to_unsigned(15, 10), 764 => to_unsigned(317, 10), 765 => to_unsigned(747, 10), 766 => to_unsigned(900, 10), 767 => to_unsigned(879, 10), 768 => to_unsigned(466, 10), 769 => to_unsigned(931, 10), 770 => to_unsigned(159, 10), 771 => to_unsigned(928, 10), 772 => to_unsigned(261, 10), 773 => to_unsigned(733, 10), 774 => to_unsigned(379, 10), 775 => to_unsigned(861, 10), 776 => to_unsigned(590, 10), 777 => to_unsigned(292, 10), 778 => to_unsigned(769, 10), 779 => to_unsigned(145, 10), 780 => to_unsigned(72, 10), 781 => to_unsigned(536, 10), 782 => to_unsigned(316, 10), 783 => to_unsigned(789, 10), 784 => to_unsigned(536, 10), 785 => to_unsigned(564, 10), 786 => to_unsigned(130, 10), 787 => to_unsigned(238, 10), 788 => to_unsigned(458, 10), 789 => to_unsigned(722, 10), 790 => to_unsigned(622, 10), 791 => to_unsigned(434, 10), 792 => to_unsigned(991, 10), 793 => to_unsigned(562, 10), 794 => to_unsigned(963, 10), 795 => to_unsigned(253, 10), 796 => to_unsigned(170, 10), 797 => to_unsigned(827, 10), 798 => to_unsigned(328, 10), 799 => to_unsigned(102, 10), 800 => to_unsigned(756, 10), 801 => to_unsigned(1015, 10), 802 => to_unsigned(813, 10), 803 => to_unsigned(96, 10), 804 => to_unsigned(847, 10), 805 => to_unsigned(80, 10), 806 => to_unsigned(391, 10), 807 => to_unsigned(95, 10), 808 => to_unsigned(670, 10), 809 => to_unsigned(869, 10), 810 => to_unsigned(641, 10), 811 => to_unsigned(20, 10), 812 => to_unsigned(345, 10), 813 => to_unsigned(179, 10), 814 => to_unsigned(236, 10), 815 => to_unsigned(629, 10), 816 => to_unsigned(587, 10), 817 => to_unsigned(921, 10), 818 => to_unsigned(639, 10), 819 => to_unsigned(938, 10), 820 => to_unsigned(639, 10), 821 => to_unsigned(819, 10), 822 => to_unsigned(166, 10), 823 => to_unsigned(902, 10), 824 => to_unsigned(406, 10), 825 => to_unsigned(356, 10), 826 => to_unsigned(161, 10), 827 => to_unsigned(491, 10), 828 => to_unsigned(394, 10), 829 => to_unsigned(817, 10), 830 => to_unsigned(35, 10), 831 => to_unsigned(442, 10), 832 => to_unsigned(59, 10), 833 => to_unsigned(543, 10), 834 => to_unsigned(904, 10), 835 => to_unsigned(644, 10), 836 => to_unsigned(521, 10), 837 => to_unsigned(128, 10), 838 => to_unsigned(342, 10), 839 => to_unsigned(104, 10), 840 => to_unsigned(822, 10), 841 => to_unsigned(601, 10), 842 => to_unsigned(810, 10), 843 => to_unsigned(806, 10), 844 => to_unsigned(138, 10), 845 => to_unsigned(871, 10), 846 => to_unsigned(247, 10), 847 => to_unsigned(861, 10), 848 => to_unsigned(301, 10), 849 => to_unsigned(18, 10), 850 => to_unsigned(533, 10), 851 => to_unsigned(693, 10), 852 => to_unsigned(394, 10), 853 => to_unsigned(421, 10), 854 => to_unsigned(430, 10), 855 => to_unsigned(307, 10), 856 => to_unsigned(133, 10), 857 => to_unsigned(502, 10), 858 => to_unsigned(259, 10), 859 => to_unsigned(1007, 10), 860 => to_unsigned(821, 10), 861 => to_unsigned(90, 10), 862 => to_unsigned(708, 10), 863 => to_unsigned(846, 10), 864 => to_unsigned(378, 10), 865 => to_unsigned(158, 10), 866 => to_unsigned(1022, 10), 867 => to_unsigned(834, 10), 868 => to_unsigned(63, 10), 869 => to_unsigned(1010, 10), 870 => to_unsigned(621, 10), 871 => to_unsigned(217, 10), 872 => to_unsigned(854, 10), 873 => to_unsigned(955, 10), 874 => to_unsigned(499, 10), 875 => to_unsigned(133, 10), 876 => to_unsigned(937, 10), 877 => to_unsigned(465, 10), 878 => to_unsigned(270, 10), 879 => to_unsigned(602, 10), 880 => to_unsigned(559, 10), 881 => to_unsigned(797, 10), 882 => to_unsigned(77, 10), 883 => to_unsigned(93, 10), 884 => to_unsigned(667, 10), 885 => to_unsigned(533, 10), 886 => to_unsigned(1003, 10), 887 => to_unsigned(550, 10), 888 => to_unsigned(320, 10), 889 => to_unsigned(563, 10), 890 => to_unsigned(810, 10), 891 => to_unsigned(55, 10), 892 => to_unsigned(717, 10), 893 => to_unsigned(467, 10), 894 => to_unsigned(274, 10), 895 => to_unsigned(610, 10), 896 => to_unsigned(476, 10), 897 => to_unsigned(952, 10), 898 => to_unsigned(503, 10), 899 => to_unsigned(160, 10), 900 => to_unsigned(617, 10), 901 => to_unsigned(159, 10), 902 => to_unsigned(703, 10), 903 => to_unsigned(259, 10), 904 => to_unsigned(908, 10), 905 => to_unsigned(54, 10), 906 => to_unsigned(521, 10), 907 => to_unsigned(567, 10), 908 => to_unsigned(374, 10), 909 => to_unsigned(1023, 10), 910 => to_unsigned(798, 10), 911 => to_unsigned(172, 10), 912 => to_unsigned(782, 10), 913 => to_unsigned(100, 10), 914 => to_unsigned(105, 10), 915 => to_unsigned(769, 10), 916 => to_unsigned(105, 10), 917 => to_unsigned(452, 10), 918 => to_unsigned(28, 10), 919 => to_unsigned(506, 10), 920 => to_unsigned(15, 10), 921 => to_unsigned(249, 10), 922 => to_unsigned(970, 10), 923 => to_unsigned(405, 10), 924 => to_unsigned(26, 10), 925 => to_unsigned(481, 10), 926 => to_unsigned(610, 10), 927 => to_unsigned(715, 10), 928 => to_unsigned(739, 10), 929 => to_unsigned(761, 10), 930 => to_unsigned(892, 10), 931 => to_unsigned(559, 10), 932 => to_unsigned(593, 10), 933 => to_unsigned(582, 10), 934 => to_unsigned(912, 10), 935 => to_unsigned(179, 10), 936 => to_unsigned(384, 10), 937 => to_unsigned(776, 10), 938 => to_unsigned(400, 10), 939 => to_unsigned(392, 10), 940 => to_unsigned(460, 10), 941 => to_unsigned(681, 10), 942 => to_unsigned(418, 10), 943 => to_unsigned(489, 10), 944 => to_unsigned(181, 10), 945 => to_unsigned(84, 10), 946 => to_unsigned(363, 10), 947 => to_unsigned(116, 10), 948 => to_unsigned(534, 10), 949 => to_unsigned(421, 10), 950 => to_unsigned(270, 10), 951 => to_unsigned(627, 10), 952 => to_unsigned(294, 10), 953 => to_unsigned(800, 10), 954 => to_unsigned(191, 10), 955 => to_unsigned(470, 10), 956 => to_unsigned(717, 10), 957 => to_unsigned(423, 10), 958 => to_unsigned(652, 10), 959 => to_unsigned(239, 10), 960 => to_unsigned(386, 10), 961 => to_unsigned(303, 10), 962 => to_unsigned(536, 10), 963 => to_unsigned(954, 10), 964 => to_unsigned(794, 10), 965 => to_unsigned(150, 10), 966 => to_unsigned(2, 10), 967 => to_unsigned(948, 10), 968 => to_unsigned(798, 10), 969 => to_unsigned(681, 10), 970 => to_unsigned(164, 10), 971 => to_unsigned(552, 10), 972 => to_unsigned(204, 10), 973 => to_unsigned(713, 10), 974 => to_unsigned(235, 10), 975 => to_unsigned(88, 10), 976 => to_unsigned(122, 10), 977 => to_unsigned(884, 10), 978 => to_unsigned(791, 10), 979 => to_unsigned(885, 10), 980 => to_unsigned(417, 10), 981 => to_unsigned(668, 10), 982 => to_unsigned(97, 10), 983 => to_unsigned(234, 10), 984 => to_unsigned(660, 10), 985 => to_unsigned(70, 10), 986 => to_unsigned(498, 10), 987 => to_unsigned(486, 10), 988 => to_unsigned(244, 10), 989 => to_unsigned(432, 10), 990 => to_unsigned(955, 10), 991 => to_unsigned(901, 10), 992 => to_unsigned(100, 10), 993 => to_unsigned(914, 10), 994 => to_unsigned(933, 10), 995 => to_unsigned(734, 10), 996 => to_unsigned(924, 10), 997 => to_unsigned(393, 10), 998 => to_unsigned(144, 10), 999 => to_unsigned(501, 10), 1000 => to_unsigned(216, 10), 1001 => to_unsigned(340, 10), 1002 => to_unsigned(521, 10), 1003 => to_unsigned(152, 10), 1004 => to_unsigned(569, 10), 1005 => to_unsigned(955, 10), 1006 => to_unsigned(467, 10), 1007 => to_unsigned(525, 10), 1008 => to_unsigned(28, 10), 1009 => to_unsigned(390, 10), 1010 => to_unsigned(61, 10), 1011 => to_unsigned(91, 10), 1012 => to_unsigned(435, 10), 1013 => to_unsigned(176, 10), 1014 => to_unsigned(830, 10), 1015 => to_unsigned(784, 10), 1016 => to_unsigned(223, 10), 1017 => to_unsigned(34, 10), 1018 => to_unsigned(483, 10), 1019 => to_unsigned(222, 10), 1020 => to_unsigned(585, 10), 1021 => to_unsigned(280, 10), 1022 => to_unsigned(851, 10), 1023 => to_unsigned(875, 10), 1024 => to_unsigned(700, 10), 1025 => to_unsigned(756, 10), 1026 => to_unsigned(336, 10), 1027 => to_unsigned(1014, 10), 1028 => to_unsigned(946, 10), 1029 => to_unsigned(704, 10), 1030 => to_unsigned(648, 10), 1031 => to_unsigned(958, 10), 1032 => to_unsigned(468, 10), 1033 => to_unsigned(79, 10), 1034 => to_unsigned(576, 10), 1035 => to_unsigned(900, 10), 1036 => to_unsigned(651, 10), 1037 => to_unsigned(187, 10), 1038 => to_unsigned(694, 10), 1039 => to_unsigned(965, 10), 1040 => to_unsigned(192, 10), 1041 => to_unsigned(568, 10), 1042 => to_unsigned(451, 10), 1043 => to_unsigned(575, 10), 1044 => to_unsigned(72, 10), 1045 => to_unsigned(39, 10), 1046 => to_unsigned(117, 10), 1047 => to_unsigned(516, 10), 1048 => to_unsigned(352, 10), 1049 => to_unsigned(898, 10), 1050 => to_unsigned(693, 10), 1051 => to_unsigned(106, 10), 1052 => to_unsigned(336, 10), 1053 => to_unsigned(468, 10), 1054 => to_unsigned(280, 10), 1055 => to_unsigned(84, 10), 1056 => to_unsigned(590, 10), 1057 => to_unsigned(1018, 10), 1058 => to_unsigned(784, 10), 1059 => to_unsigned(218, 10), 1060 => to_unsigned(956, 10), 1061 => to_unsigned(715, 10), 1062 => to_unsigned(1012, 10), 1063 => to_unsigned(681, 10), 1064 => to_unsigned(669, 10), 1065 => to_unsigned(758, 10), 1066 => to_unsigned(579, 10), 1067 => to_unsigned(446, 10), 1068 => to_unsigned(277, 10), 1069 => to_unsigned(22, 10), 1070 => to_unsigned(439, 10), 1071 => to_unsigned(398, 10), 1072 => to_unsigned(448, 10), 1073 => to_unsigned(35, 10), 1074 => to_unsigned(457, 10), 1075 => to_unsigned(319, 10), 1076 => to_unsigned(782, 10), 1077 => to_unsigned(60, 10), 1078 => to_unsigned(760, 10), 1079 => to_unsigned(735, 10), 1080 => to_unsigned(210, 10), 1081 => to_unsigned(448, 10), 1082 => to_unsigned(598, 10), 1083 => to_unsigned(889, 10), 1084 => to_unsigned(109, 10), 1085 => to_unsigned(33, 10), 1086 => to_unsigned(310, 10), 1087 => to_unsigned(414, 10), 1088 => to_unsigned(15, 10), 1089 => to_unsigned(543, 10), 1090 => to_unsigned(940, 10), 1091 => to_unsigned(34, 10), 1092 => to_unsigned(137, 10), 1093 => to_unsigned(185, 10), 1094 => to_unsigned(206, 10), 1095 => to_unsigned(280, 10), 1096 => to_unsigned(710, 10), 1097 => to_unsigned(600, 10), 1098 => to_unsigned(617, 10), 1099 => to_unsigned(518, 10), 1100 => to_unsigned(918, 10), 1101 => to_unsigned(234, 10), 1102 => to_unsigned(335, 10), 1103 => to_unsigned(39, 10), 1104 => to_unsigned(181, 10), 1105 => to_unsigned(310, 10), 1106 => to_unsigned(448, 10), 1107 => to_unsigned(513, 10), 1108 => to_unsigned(920, 10), 1109 => to_unsigned(883, 10), 1110 => to_unsigned(385, 10), 1111 => to_unsigned(146, 10), 1112 => to_unsigned(778, 10), 1113 => to_unsigned(112, 10), 1114 => to_unsigned(513, 10), 1115 => to_unsigned(229, 10), 1116 => to_unsigned(791, 10), 1117 => to_unsigned(318, 10), 1118 => to_unsigned(596, 10), 1119 => to_unsigned(839, 10), 1120 => to_unsigned(1011, 10), 1121 => to_unsigned(131, 10), 1122 => to_unsigned(26, 10), 1123 => to_unsigned(526, 10), 1124 => to_unsigned(3, 10), 1125 => to_unsigned(367, 10), 1126 => to_unsigned(425, 10), 1127 => to_unsigned(1012, 10), 1128 => to_unsigned(424, 10), 1129 => to_unsigned(732, 10), 1130 => to_unsigned(150, 10), 1131 => to_unsigned(712, 10), 1132 => to_unsigned(896, 10), 1133 => to_unsigned(545, 10), 1134 => to_unsigned(337, 10), 1135 => to_unsigned(754, 10), 1136 => to_unsigned(461, 10), 1137 => to_unsigned(380, 10), 1138 => to_unsigned(745, 10), 1139 => to_unsigned(789, 10), 1140 => to_unsigned(421, 10), 1141 => to_unsigned(842, 10), 1142 => to_unsigned(825, 10), 1143 => to_unsigned(724, 10), 1144 => to_unsigned(115, 10), 1145 => to_unsigned(823, 10), 1146 => to_unsigned(658, 10), 1147 => to_unsigned(312, 10), 1148 => to_unsigned(11, 10), 1149 => to_unsigned(252, 10), 1150 => to_unsigned(447, 10), 1151 => to_unsigned(953, 10), 1152 => to_unsigned(186, 10), 1153 => to_unsigned(455, 10), 1154 => to_unsigned(484, 10), 1155 => to_unsigned(71, 10), 1156 => to_unsigned(685, 10), 1157 => to_unsigned(790, 10), 1158 => to_unsigned(207, 10), 1159 => to_unsigned(419, 10), 1160 => to_unsigned(628, 10), 1161 => to_unsigned(839, 10), 1162 => to_unsigned(917, 10), 1163 => to_unsigned(66, 10), 1164 => to_unsigned(263, 10), 1165 => to_unsigned(620, 10), 1166 => to_unsigned(686, 10), 1167 => to_unsigned(536, 10), 1168 => to_unsigned(789, 10), 1169 => to_unsigned(1020, 10), 1170 => to_unsigned(379, 10), 1171 => to_unsigned(337, 10), 1172 => to_unsigned(251, 10), 1173 => to_unsigned(278, 10), 1174 => to_unsigned(22, 10), 1175 => to_unsigned(164, 10), 1176 => to_unsigned(384, 10), 1177 => to_unsigned(712, 10), 1178 => to_unsigned(474, 10), 1179 => to_unsigned(370, 10), 1180 => to_unsigned(73, 10), 1181 => to_unsigned(725, 10), 1182 => to_unsigned(292, 10), 1183 => to_unsigned(776, 10), 1184 => to_unsigned(322, 10), 1185 => to_unsigned(423, 10), 1186 => to_unsigned(823, 10), 1187 => to_unsigned(859, 10), 1188 => to_unsigned(580, 10), 1189 => to_unsigned(497, 10), 1190 => to_unsigned(254, 10), 1191 => to_unsigned(313, 10), 1192 => to_unsigned(581, 10), 1193 => to_unsigned(108, 10), 1194 => to_unsigned(863, 10), 1195 => to_unsigned(846, 10), 1196 => to_unsigned(180, 10), 1197 => to_unsigned(280, 10), 1198 => to_unsigned(591, 10), 1199 => to_unsigned(119, 10), 1200 => to_unsigned(308, 10), 1201 => to_unsigned(643, 10), 1202 => to_unsigned(1003, 10), 1203 => to_unsigned(240, 10), 1204 => to_unsigned(916, 10), 1205 => to_unsigned(866, 10), 1206 => to_unsigned(647, 10), 1207 => to_unsigned(866, 10), 1208 => to_unsigned(890, 10), 1209 => to_unsigned(661, 10), 1210 => to_unsigned(516, 10), 1211 => to_unsigned(342, 10), 1212 => to_unsigned(521, 10), 1213 => to_unsigned(754, 10), 1214 => to_unsigned(1012, 10), 1215 => to_unsigned(725, 10), 1216 => to_unsigned(44, 10), 1217 => to_unsigned(62, 10), 1218 => to_unsigned(596, 10), 1219 => to_unsigned(899, 10), 1220 => to_unsigned(137, 10), 1221 => to_unsigned(473, 10), 1222 => to_unsigned(816, 10), 1223 => to_unsigned(190, 10), 1224 => to_unsigned(234, 10), 1225 => to_unsigned(521, 10), 1226 => to_unsigned(496, 10), 1227 => to_unsigned(141, 10), 1228 => to_unsigned(752, 10), 1229 => to_unsigned(782, 10), 1230 => to_unsigned(198, 10), 1231 => to_unsigned(675, 10), 1232 => to_unsigned(729, 10), 1233 => to_unsigned(594, 10), 1234 => to_unsigned(748, 10), 1235 => to_unsigned(393, 10), 1236 => to_unsigned(859, 10), 1237 => to_unsigned(823, 10), 1238 => to_unsigned(772, 10), 1239 => to_unsigned(769, 10), 1240 => to_unsigned(355, 10), 1241 => to_unsigned(903, 10), 1242 => to_unsigned(448, 10), 1243 => to_unsigned(823, 10), 1244 => to_unsigned(638, 10), 1245 => to_unsigned(71, 10), 1246 => to_unsigned(365, 10), 1247 => to_unsigned(349, 10), 1248 => to_unsigned(580, 10), 1249 => to_unsigned(774, 10), 1250 => to_unsigned(592, 10), 1251 => to_unsigned(987, 10), 1252 => to_unsigned(579, 10), 1253 => to_unsigned(43, 10), 1254 => to_unsigned(577, 10), 1255 => to_unsigned(559, 10), 1256 => to_unsigned(610, 10), 1257 => to_unsigned(494, 10), 1258 => to_unsigned(913, 10), 1259 => to_unsigned(293, 10), 1260 => to_unsigned(749, 10), 1261 => to_unsigned(826, 10), 1262 => to_unsigned(549, 10), 1263 => to_unsigned(304, 10), 1264 => to_unsigned(1019, 10), 1265 => to_unsigned(934, 10), 1266 => to_unsigned(1005, 10), 1267 => to_unsigned(557, 10), 1268 => to_unsigned(506, 10), 1269 => to_unsigned(36, 10), 1270 => to_unsigned(343, 10), 1271 => to_unsigned(761, 10), 1272 => to_unsigned(666, 10), 1273 => to_unsigned(929, 10), 1274 => to_unsigned(810, 10), 1275 => to_unsigned(883, 10), 1276 => to_unsigned(223, 10), 1277 => to_unsigned(209, 10), 1278 => to_unsigned(405, 10), 1279 => to_unsigned(117, 10), 1280 => to_unsigned(748, 10), 1281 => to_unsigned(927, 10), 1282 => to_unsigned(907, 10), 1283 => to_unsigned(834, 10), 1284 => to_unsigned(298, 10), 1285 => to_unsigned(609, 10), 1286 => to_unsigned(790, 10), 1287 => to_unsigned(395, 10), 1288 => to_unsigned(488, 10), 1289 => to_unsigned(507, 10), 1290 => to_unsigned(941, 10), 1291 => to_unsigned(688, 10), 1292 => to_unsigned(862, 10), 1293 => to_unsigned(787, 10), 1294 => to_unsigned(294, 10), 1295 => to_unsigned(870, 10), 1296 => to_unsigned(964, 10), 1297 => to_unsigned(373, 10), 1298 => to_unsigned(269, 10), 1299 => to_unsigned(813, 10), 1300 => to_unsigned(624, 10), 1301 => to_unsigned(495, 10), 1302 => to_unsigned(90, 10), 1303 => to_unsigned(1018, 10), 1304 => to_unsigned(373, 10), 1305 => to_unsigned(38, 10), 1306 => to_unsigned(350, 10), 1307 => to_unsigned(526, 10), 1308 => to_unsigned(444, 10), 1309 => to_unsigned(611, 10), 1310 => to_unsigned(607, 10), 1311 => to_unsigned(182, 10), 1312 => to_unsigned(202, 10), 1313 => to_unsigned(611, 10), 1314 => to_unsigned(1002, 10), 1315 => to_unsigned(462, 10), 1316 => to_unsigned(275, 10), 1317 => to_unsigned(425, 10), 1318 => to_unsigned(795, 10), 1319 => to_unsigned(490, 10), 1320 => to_unsigned(389, 10), 1321 => to_unsigned(439, 10), 1322 => to_unsigned(728, 10), 1323 => to_unsigned(584, 10), 1324 => to_unsigned(1006, 10), 1325 => to_unsigned(787, 10), 1326 => to_unsigned(293, 10), 1327 => to_unsigned(333, 10), 1328 => to_unsigned(222, 10), 1329 => to_unsigned(879, 10), 1330 => to_unsigned(0, 10), 1331 => to_unsigned(651, 10), 1332 => to_unsigned(34, 10), 1333 => to_unsigned(12, 10), 1334 => to_unsigned(563, 10), 1335 => to_unsigned(667, 10), 1336 => to_unsigned(627, 10), 1337 => to_unsigned(377, 10), 1338 => to_unsigned(679, 10), 1339 => to_unsigned(544, 10), 1340 => to_unsigned(411, 10), 1341 => to_unsigned(774, 10), 1342 => to_unsigned(694, 10), 1343 => to_unsigned(604, 10), 1344 => to_unsigned(273, 10), 1345 => to_unsigned(708, 10), 1346 => to_unsigned(152, 10), 1347 => to_unsigned(731, 10), 1348 => to_unsigned(18, 10), 1349 => to_unsigned(82, 10), 1350 => to_unsigned(990, 10), 1351 => to_unsigned(901, 10), 1352 => to_unsigned(158, 10), 1353 => to_unsigned(744, 10), 1354 => to_unsigned(511, 10), 1355 => to_unsigned(587, 10), 1356 => to_unsigned(953, 10), 1357 => to_unsigned(997, 10), 1358 => to_unsigned(62, 10), 1359 => to_unsigned(316, 10), 1360 => to_unsigned(439, 10), 1361 => to_unsigned(734, 10), 1362 => to_unsigned(129, 10), 1363 => to_unsigned(278, 10), 1364 => to_unsigned(517, 10), 1365 => to_unsigned(228, 10), 1366 => to_unsigned(722, 10), 1367 => to_unsigned(770, 10), 1368 => to_unsigned(304, 10), 1369 => to_unsigned(46, 10), 1370 => to_unsigned(498, 10), 1371 => to_unsigned(427, 10), 1372 => to_unsigned(445, 10), 1373 => to_unsigned(521, 10), 1374 => to_unsigned(418, 10), 1375 => to_unsigned(881, 10), 1376 => to_unsigned(841, 10), 1377 => to_unsigned(907, 10), 1378 => to_unsigned(423, 10), 1379 => to_unsigned(551, 10), 1380 => to_unsigned(993, 10), 1381 => to_unsigned(22, 10), 1382 => to_unsigned(488, 10), 1383 => to_unsigned(436, 10), 1384 => to_unsigned(755, 10), 1385 => to_unsigned(105, 10), 1386 => to_unsigned(449, 10), 1387 => to_unsigned(543, 10), 1388 => to_unsigned(1021, 10), 1389 => to_unsigned(531, 10), 1390 => to_unsigned(312, 10), 1391 => to_unsigned(538, 10), 1392 => to_unsigned(764, 10), 1393 => to_unsigned(190, 10), 1394 => to_unsigned(20, 10), 1395 => to_unsigned(997, 10), 1396 => to_unsigned(292, 10), 1397 => to_unsigned(833, 10), 1398 => to_unsigned(877, 10), 1399 => to_unsigned(274, 10), 1400 => to_unsigned(71, 10), 1401 => to_unsigned(611, 10), 1402 => to_unsigned(577, 10), 1403 => to_unsigned(248, 10), 1404 => to_unsigned(635, 10), 1405 => to_unsigned(442, 10), 1406 => to_unsigned(684, 10), 1407 => to_unsigned(221, 10), 1408 => to_unsigned(844, 10), 1409 => to_unsigned(1016, 10), 1410 => to_unsigned(574, 10), 1411 => to_unsigned(183, 10), 1412 => to_unsigned(789, 10), 1413 => to_unsigned(418, 10), 1414 => to_unsigned(421, 10), 1415 => to_unsigned(194, 10), 1416 => to_unsigned(800, 10), 1417 => to_unsigned(888, 10), 1418 => to_unsigned(375, 10), 1419 => to_unsigned(246, 10), 1420 => to_unsigned(964, 10), 1421 => to_unsigned(878, 10), 1422 => to_unsigned(222, 10), 1423 => to_unsigned(693, 10), 1424 => to_unsigned(244, 10), 1425 => to_unsigned(435, 10), 1426 => to_unsigned(531, 10), 1427 => to_unsigned(321, 10), 1428 => to_unsigned(235, 10), 1429 => to_unsigned(281, 10), 1430 => to_unsigned(48, 10), 1431 => to_unsigned(988, 10), 1432 => to_unsigned(906, 10), 1433 => to_unsigned(652, 10), 1434 => to_unsigned(845, 10), 1435 => to_unsigned(446, 10), 1436 => to_unsigned(70, 10), 1437 => to_unsigned(866, 10), 1438 => to_unsigned(574, 10), 1439 => to_unsigned(424, 10), 1440 => to_unsigned(141, 10), 1441 => to_unsigned(594, 10), 1442 => to_unsigned(373, 10), 1443 => to_unsigned(972, 10), 1444 => to_unsigned(924, 10), 1445 => to_unsigned(632, 10), 1446 => to_unsigned(15, 10), 1447 => to_unsigned(523, 10), 1448 => to_unsigned(705, 10), 1449 => to_unsigned(874, 10), 1450 => to_unsigned(524, 10), 1451 => to_unsigned(649, 10), 1452 => to_unsigned(415, 10), 1453 => to_unsigned(659, 10), 1454 => to_unsigned(297, 10), 1455 => to_unsigned(497, 10), 1456 => to_unsigned(598, 10), 1457 => to_unsigned(415, 10), 1458 => to_unsigned(346, 10), 1459 => to_unsigned(485, 10), 1460 => to_unsigned(159, 10), 1461 => to_unsigned(749, 10), 1462 => to_unsigned(41, 10), 1463 => to_unsigned(31, 10), 1464 => to_unsigned(382, 10), 1465 => to_unsigned(467, 10), 1466 => to_unsigned(531, 10), 1467 => to_unsigned(748, 10), 1468 => to_unsigned(232, 10), 1469 => to_unsigned(88, 10), 1470 => to_unsigned(302, 10), 1471 => to_unsigned(684, 10), 1472 => to_unsigned(556, 10), 1473 => to_unsigned(141, 10), 1474 => to_unsigned(810, 10), 1475 => to_unsigned(799, 10), 1476 => to_unsigned(102, 10), 1477 => to_unsigned(134, 10), 1478 => to_unsigned(748, 10), 1479 => to_unsigned(456, 10), 1480 => to_unsigned(973, 10), 1481 => to_unsigned(689, 10), 1482 => to_unsigned(743, 10), 1483 => to_unsigned(172, 10), 1484 => to_unsigned(442, 10), 1485 => to_unsigned(451, 10), 1486 => to_unsigned(376, 10), 1487 => to_unsigned(426, 10), 1488 => to_unsigned(202, 10), 1489 => to_unsigned(582, 10), 1490 => to_unsigned(148, 10), 1491 => to_unsigned(392, 10), 1492 => to_unsigned(284, 10), 1493 => to_unsigned(181, 10), 1494 => to_unsigned(208, 10), 1495 => to_unsigned(411, 10), 1496 => to_unsigned(506, 10), 1497 => to_unsigned(442, 10), 1498 => to_unsigned(419, 10), 1499 => to_unsigned(621, 10), 1500 => to_unsigned(664, 10), 1501 => to_unsigned(769, 10), 1502 => to_unsigned(641, 10), 1503 => to_unsigned(820, 10), 1504 => to_unsigned(702, 10), 1505 => to_unsigned(117, 10), 1506 => to_unsigned(153, 10), 1507 => to_unsigned(154, 10), 1508 => to_unsigned(961, 10), 1509 => to_unsigned(971, 10), 1510 => to_unsigned(96, 10), 1511 => to_unsigned(204, 10), 1512 => to_unsigned(698, 10), 1513 => to_unsigned(92, 10), 1514 => to_unsigned(321, 10), 1515 => to_unsigned(454, 10), 1516 => to_unsigned(843, 10), 1517 => to_unsigned(71, 10), 1518 => to_unsigned(197, 10), 1519 => to_unsigned(12, 10), 1520 => to_unsigned(32, 10), 1521 => to_unsigned(90, 10), 1522 => to_unsigned(751, 10), 1523 => to_unsigned(704, 10), 1524 => to_unsigned(597, 10), 1525 => to_unsigned(984, 10), 1526 => to_unsigned(845, 10), 1527 => to_unsigned(294, 10), 1528 => to_unsigned(280, 10), 1529 => to_unsigned(370, 10), 1530 => to_unsigned(430, 10), 1531 => to_unsigned(101, 10), 1532 => to_unsigned(585, 10), 1533 => to_unsigned(543, 10), 1534 => to_unsigned(689, 10), 1535 => to_unsigned(4, 10), 1536 => to_unsigned(347, 10), 1537 => to_unsigned(701, 10), 1538 => to_unsigned(28, 10), 1539 => to_unsigned(848, 10), 1540 => to_unsigned(692, 10), 1541 => to_unsigned(663, 10), 1542 => to_unsigned(339, 10), 1543 => to_unsigned(367, 10), 1544 => to_unsigned(200, 10), 1545 => to_unsigned(368, 10), 1546 => to_unsigned(532, 10), 1547 => to_unsigned(307, 10), 1548 => to_unsigned(759, 10), 1549 => to_unsigned(253, 10), 1550 => to_unsigned(557, 10), 1551 => to_unsigned(490, 10), 1552 => to_unsigned(536, 10), 1553 => to_unsigned(700, 10), 1554 => to_unsigned(627, 10), 1555 => to_unsigned(278, 10), 1556 => to_unsigned(531, 10), 1557 => to_unsigned(411, 10), 1558 => to_unsigned(386, 10), 1559 => to_unsigned(637, 10), 1560 => to_unsigned(818, 10), 1561 => to_unsigned(1014, 10), 1562 => to_unsigned(852, 10), 1563 => to_unsigned(205, 10), 1564 => to_unsigned(1023, 10), 1565 => to_unsigned(931, 10), 1566 => to_unsigned(889, 10), 1567 => to_unsigned(294, 10), 1568 => to_unsigned(976, 10), 1569 => to_unsigned(685, 10), 1570 => to_unsigned(160, 10), 1571 => to_unsigned(194, 10), 1572 => to_unsigned(530, 10), 1573 => to_unsigned(217, 10), 1574 => to_unsigned(939, 10), 1575 => to_unsigned(515, 10), 1576 => to_unsigned(147, 10), 1577 => to_unsigned(816, 10), 1578 => to_unsigned(312, 10), 1579 => to_unsigned(913, 10), 1580 => to_unsigned(788, 10), 1581 => to_unsigned(981, 10), 1582 => to_unsigned(424, 10), 1583 => to_unsigned(1001, 10), 1584 => to_unsigned(48, 10), 1585 => to_unsigned(966, 10), 1586 => to_unsigned(272, 10), 1587 => to_unsigned(193, 10), 1588 => to_unsigned(460, 10), 1589 => to_unsigned(942, 10), 1590 => to_unsigned(181, 10), 1591 => to_unsigned(272, 10), 1592 => to_unsigned(661, 10), 1593 => to_unsigned(754, 10), 1594 => to_unsigned(333, 10), 1595 => to_unsigned(514, 10), 1596 => to_unsigned(195, 10), 1597 => to_unsigned(913, 10), 1598 => to_unsigned(841, 10), 1599 => to_unsigned(567, 10), 1600 => to_unsigned(804, 10), 1601 => to_unsigned(269, 10), 1602 => to_unsigned(17, 10), 1603 => to_unsigned(957, 10), 1604 => to_unsigned(692, 10), 1605 => to_unsigned(380, 10), 1606 => to_unsigned(417, 10), 1607 => to_unsigned(962, 10), 1608 => to_unsigned(277, 10), 1609 => to_unsigned(433, 10), 1610 => to_unsigned(998, 10), 1611 => to_unsigned(946, 10), 1612 => to_unsigned(238, 10), 1613 => to_unsigned(914, 10), 1614 => to_unsigned(218, 10), 1615 => to_unsigned(76, 10), 1616 => to_unsigned(960, 10), 1617 => to_unsigned(575, 10), 1618 => to_unsigned(501, 10), 1619 => to_unsigned(143, 10), 1620 => to_unsigned(628, 10), 1621 => to_unsigned(518, 10), 1622 => to_unsigned(775, 10), 1623 => to_unsigned(307, 10), 1624 => to_unsigned(100, 10), 1625 => to_unsigned(888, 10), 1626 => to_unsigned(559, 10), 1627 => to_unsigned(17, 10), 1628 => to_unsigned(390, 10), 1629 => to_unsigned(657, 10), 1630 => to_unsigned(452, 10), 1631 => to_unsigned(15, 10), 1632 => to_unsigned(720, 10), 1633 => to_unsigned(753, 10), 1634 => to_unsigned(554, 10), 1635 => to_unsigned(974, 10), 1636 => to_unsigned(709, 10), 1637 => to_unsigned(716, 10), 1638 => to_unsigned(467, 10), 1639 => to_unsigned(613, 10), 1640 => to_unsigned(846, 10), 1641 => to_unsigned(470, 10), 1642 => to_unsigned(234, 10), 1643 => to_unsigned(197, 10), 1644 => to_unsigned(193, 10), 1645 => to_unsigned(373, 10), 1646 => to_unsigned(579, 10), 1647 => to_unsigned(958, 10), 1648 => to_unsigned(333, 10), 1649 => to_unsigned(511, 10), 1650 => to_unsigned(186, 10), 1651 => to_unsigned(281, 10), 1652 => to_unsigned(255, 10), 1653 => to_unsigned(774, 10), 1654 => to_unsigned(142, 10), 1655 => to_unsigned(781, 10), 1656 => to_unsigned(717, 10), 1657 => to_unsigned(989, 10), 1658 => to_unsigned(384, 10), 1659 => to_unsigned(959, 10), 1660 => to_unsigned(105, 10), 1661 => to_unsigned(347, 10), 1662 => to_unsigned(606, 10), 1663 => to_unsigned(29, 10), 1664 => to_unsigned(405, 10), 1665 => to_unsigned(532, 10), 1666 => to_unsigned(411, 10), 1667 => to_unsigned(933, 10), 1668 => to_unsigned(532, 10), 1669 => to_unsigned(177, 10), 1670 => to_unsigned(217, 10), 1671 => to_unsigned(120, 10), 1672 => to_unsigned(629, 10), 1673 => to_unsigned(803, 10), 1674 => to_unsigned(52, 10), 1675 => to_unsigned(108, 10), 1676 => to_unsigned(98, 10), 1677 => to_unsigned(760, 10), 1678 => to_unsigned(384, 10), 1679 => to_unsigned(80, 10), 1680 => to_unsigned(793, 10), 1681 => to_unsigned(25, 10), 1682 => to_unsigned(353, 10), 1683 => to_unsigned(686, 10), 1684 => to_unsigned(462, 10), 1685 => to_unsigned(818, 10), 1686 => to_unsigned(235, 10), 1687 => to_unsigned(447, 10), 1688 => to_unsigned(196, 10), 1689 => to_unsigned(263, 10), 1690 => to_unsigned(10, 10), 1691 => to_unsigned(35, 10), 1692 => to_unsigned(946, 10), 1693 => to_unsigned(828, 10), 1694 => to_unsigned(201, 10), 1695 => to_unsigned(897, 10), 1696 => to_unsigned(502, 10), 1697 => to_unsigned(454, 10), 1698 => to_unsigned(525, 10), 1699 => to_unsigned(199, 10), 1700 => to_unsigned(301, 10), 1701 => to_unsigned(433, 10), 1702 => to_unsigned(154, 10), 1703 => to_unsigned(340, 10), 1704 => to_unsigned(899, 10), 1705 => to_unsigned(324, 10), 1706 => to_unsigned(486, 10), 1707 => to_unsigned(982, 10), 1708 => to_unsigned(674, 10), 1709 => to_unsigned(584, 10), 1710 => to_unsigned(874, 10), 1711 => to_unsigned(643, 10), 1712 => to_unsigned(192, 10), 1713 => to_unsigned(766, 10), 1714 => to_unsigned(598, 10), 1715 => to_unsigned(513, 10), 1716 => to_unsigned(551, 10), 1717 => to_unsigned(339, 10), 1718 => to_unsigned(177, 10), 1719 => to_unsigned(436, 10), 1720 => to_unsigned(69, 10), 1721 => to_unsigned(426, 10), 1722 => to_unsigned(832, 10), 1723 => to_unsigned(299, 10), 1724 => to_unsigned(426, 10), 1725 => to_unsigned(524, 10), 1726 => to_unsigned(854, 10), 1727 => to_unsigned(362, 10), 1728 => to_unsigned(942, 10), 1729 => to_unsigned(558, 10), 1730 => to_unsigned(586, 10), 1731 => to_unsigned(293, 10), 1732 => to_unsigned(704, 10), 1733 => to_unsigned(755, 10), 1734 => to_unsigned(290, 10), 1735 => to_unsigned(648, 10), 1736 => to_unsigned(80, 10), 1737 => to_unsigned(62, 10), 1738 => to_unsigned(334, 10), 1739 => to_unsigned(406, 10), 1740 => to_unsigned(101, 10), 1741 => to_unsigned(981, 10), 1742 => to_unsigned(563, 10), 1743 => to_unsigned(554, 10), 1744 => to_unsigned(134, 10), 1745 => to_unsigned(162, 10), 1746 => to_unsigned(519, 10), 1747 => to_unsigned(918, 10), 1748 => to_unsigned(584, 10), 1749 => to_unsigned(521, 10), 1750 => to_unsigned(263, 10), 1751 => to_unsigned(311, 10), 1752 => to_unsigned(862, 10), 1753 => to_unsigned(744, 10), 1754 => to_unsigned(18, 10), 1755 => to_unsigned(524, 10), 1756 => to_unsigned(191, 10), 1757 => to_unsigned(232, 10), 1758 => to_unsigned(412, 10), 1759 => to_unsigned(1001, 10), 1760 => to_unsigned(39, 10), 1761 => to_unsigned(191, 10), 1762 => to_unsigned(882, 10), 1763 => to_unsigned(650, 10), 1764 => to_unsigned(706, 10), 1765 => to_unsigned(1010, 10), 1766 => to_unsigned(355, 10), 1767 => to_unsigned(66, 10), 1768 => to_unsigned(505, 10), 1769 => to_unsigned(220, 10), 1770 => to_unsigned(358, 10), 1771 => to_unsigned(17, 10), 1772 => to_unsigned(922, 10), 1773 => to_unsigned(564, 10), 1774 => to_unsigned(682, 10), 1775 => to_unsigned(922, 10), 1776 => to_unsigned(51, 10), 1777 => to_unsigned(714, 10), 1778 => to_unsigned(156, 10), 1779 => to_unsigned(733, 10), 1780 => to_unsigned(102, 10), 1781 => to_unsigned(569, 10), 1782 => to_unsigned(604, 10), 1783 => to_unsigned(326, 10), 1784 => to_unsigned(334, 10), 1785 => to_unsigned(251, 10), 1786 => to_unsigned(1004, 10), 1787 => to_unsigned(456, 10), 1788 => to_unsigned(926, 10), 1789 => to_unsigned(519, 10), 1790 => to_unsigned(468, 10), 1791 => to_unsigned(858, 10), 1792 => to_unsigned(221, 10), 1793 => to_unsigned(458, 10), 1794 => to_unsigned(764, 10), 1795 => to_unsigned(678, 10), 1796 => to_unsigned(23, 10), 1797 => to_unsigned(472, 10), 1798 => to_unsigned(817, 10), 1799 => to_unsigned(604, 10), 1800 => to_unsigned(385, 10), 1801 => to_unsigned(909, 10), 1802 => to_unsigned(194, 10), 1803 => to_unsigned(297, 10), 1804 => to_unsigned(560, 10), 1805 => to_unsigned(172, 10), 1806 => to_unsigned(251, 10), 1807 => to_unsigned(974, 10), 1808 => to_unsigned(105, 10), 1809 => to_unsigned(787, 10), 1810 => to_unsigned(484, 10), 1811 => to_unsigned(607, 10), 1812 => to_unsigned(623, 10), 1813 => to_unsigned(283, 10), 1814 => to_unsigned(734, 10), 1815 => to_unsigned(1, 10), 1816 => to_unsigned(81, 10), 1817 => to_unsigned(405, 10), 1818 => to_unsigned(457, 10), 1819 => to_unsigned(783, 10), 1820 => to_unsigned(92, 10), 1821 => to_unsigned(19, 10), 1822 => to_unsigned(956, 10), 1823 => to_unsigned(149, 10), 1824 => to_unsigned(86, 10), 1825 => to_unsigned(484, 10), 1826 => to_unsigned(376, 10), 1827 => to_unsigned(144, 10), 1828 => to_unsigned(371, 10), 1829 => to_unsigned(690, 10), 1830 => to_unsigned(235, 10), 1831 => to_unsigned(357, 10), 1832 => to_unsigned(345, 10), 1833 => to_unsigned(506, 10), 1834 => to_unsigned(244, 10), 1835 => to_unsigned(93, 10), 1836 => to_unsigned(719, 10), 1837 => to_unsigned(153, 10), 1838 => to_unsigned(639, 10), 1839 => to_unsigned(298, 10), 1840 => to_unsigned(828, 10), 1841 => to_unsigned(1023, 10), 1842 => to_unsigned(97, 10), 1843 => to_unsigned(192, 10), 1844 => to_unsigned(254, 10), 1845 => to_unsigned(1010, 10), 1846 => to_unsigned(343, 10), 1847 => to_unsigned(314, 10), 1848 => to_unsigned(707, 10), 1849 => to_unsigned(983, 10), 1850 => to_unsigned(670, 10), 1851 => to_unsigned(350, 10), 1852 => to_unsigned(188, 10), 1853 => to_unsigned(113, 10), 1854 => to_unsigned(732, 10), 1855 => to_unsigned(835, 10), 1856 => to_unsigned(553, 10), 1857 => to_unsigned(778, 10), 1858 => to_unsigned(46, 10), 1859 => to_unsigned(165, 10), 1860 => to_unsigned(887, 10), 1861 => to_unsigned(3, 10), 1862 => to_unsigned(486, 10), 1863 => to_unsigned(422, 10), 1864 => to_unsigned(788, 10), 1865 => to_unsigned(704, 10), 1866 => to_unsigned(737, 10), 1867 => to_unsigned(1005, 10), 1868 => to_unsigned(698, 10), 1869 => to_unsigned(750, 10), 1870 => to_unsigned(633, 10), 1871 => to_unsigned(883, 10), 1872 => to_unsigned(558, 10), 1873 => to_unsigned(392, 10), 1874 => to_unsigned(523, 10), 1875 => to_unsigned(361, 10), 1876 => to_unsigned(465, 10), 1877 => to_unsigned(713, 10), 1878 => to_unsigned(549, 10), 1879 => to_unsigned(778, 10), 1880 => to_unsigned(161, 10), 1881 => to_unsigned(68, 10), 1882 => to_unsigned(234, 10), 1883 => to_unsigned(911, 10), 1884 => to_unsigned(218, 10), 1885 => to_unsigned(98, 10), 1886 => to_unsigned(137, 10), 1887 => to_unsigned(338, 10), 1888 => to_unsigned(531, 10), 1889 => to_unsigned(128, 10), 1890 => to_unsigned(416, 10), 1891 => to_unsigned(720, 10), 1892 => to_unsigned(673, 10), 1893 => to_unsigned(230, 10), 1894 => to_unsigned(503, 10), 1895 => to_unsigned(664, 10), 1896 => to_unsigned(313, 10), 1897 => to_unsigned(794, 10), 1898 => to_unsigned(994, 10), 1899 => to_unsigned(396, 10), 1900 => to_unsigned(130, 10), 1901 => to_unsigned(549, 10), 1902 => to_unsigned(140, 10), 1903 => to_unsigned(802, 10), 1904 => to_unsigned(729, 10), 1905 => to_unsigned(371, 10), 1906 => to_unsigned(659, 10), 1907 => to_unsigned(692, 10), 1908 => to_unsigned(13, 10), 1909 => to_unsigned(769, 10), 1910 => to_unsigned(580, 10), 1911 => to_unsigned(84, 10), 1912 => to_unsigned(282, 10), 1913 => to_unsigned(89, 10), 1914 => to_unsigned(407, 10), 1915 => to_unsigned(741, 10), 1916 => to_unsigned(166, 10), 1917 => to_unsigned(575, 10), 1918 => to_unsigned(948, 10), 1919 => to_unsigned(908, 10), 1920 => to_unsigned(86, 10), 1921 => to_unsigned(926, 10), 1922 => to_unsigned(203, 10), 1923 => to_unsigned(939, 10), 1924 => to_unsigned(245, 10), 1925 => to_unsigned(60, 10), 1926 => to_unsigned(315, 10), 1927 => to_unsigned(216, 10), 1928 => to_unsigned(541, 10), 1929 => to_unsigned(831, 10), 1930 => to_unsigned(702, 10), 1931 => to_unsigned(719, 10), 1932 => to_unsigned(236, 10), 1933 => to_unsigned(479, 10), 1934 => to_unsigned(477, 10), 1935 => to_unsigned(643, 10), 1936 => to_unsigned(669, 10), 1937 => to_unsigned(374, 10), 1938 => to_unsigned(225, 10), 1939 => to_unsigned(451, 10), 1940 => to_unsigned(796, 10), 1941 => to_unsigned(873, 10), 1942 => to_unsigned(977, 10), 1943 => to_unsigned(367, 10), 1944 => to_unsigned(1023, 10), 1945 => to_unsigned(595, 10), 1946 => to_unsigned(931, 10), 1947 => to_unsigned(411, 10), 1948 => to_unsigned(213, 10), 1949 => to_unsigned(247, 10), 1950 => to_unsigned(943, 10), 1951 => to_unsigned(1011, 10), 1952 => to_unsigned(328, 10), 1953 => to_unsigned(258, 10), 1954 => to_unsigned(310, 10), 1955 => to_unsigned(965, 10), 1956 => to_unsigned(985, 10), 1957 => to_unsigned(291, 10), 1958 => to_unsigned(9, 10), 1959 => to_unsigned(663, 10), 1960 => to_unsigned(624, 10), 1961 => to_unsigned(79, 10), 1962 => to_unsigned(217, 10), 1963 => to_unsigned(853, 10), 1964 => to_unsigned(108, 10), 1965 => to_unsigned(55, 10), 1966 => to_unsigned(385, 10), 1967 => to_unsigned(347, 10), 1968 => to_unsigned(434, 10), 1969 => to_unsigned(988, 10), 1970 => to_unsigned(372, 10), 1971 => to_unsigned(842, 10), 1972 => to_unsigned(1011, 10), 1973 => to_unsigned(343, 10), 1974 => to_unsigned(450, 10), 1975 => to_unsigned(82, 10), 1976 => to_unsigned(163, 10), 1977 => to_unsigned(902, 10), 1978 => to_unsigned(875, 10), 1979 => to_unsigned(842, 10), 1980 => to_unsigned(103, 10), 1981 => to_unsigned(742, 10), 1982 => to_unsigned(1002, 10), 1983 => to_unsigned(227, 10), 1984 => to_unsigned(355, 10), 1985 => to_unsigned(542, 10), 1986 => to_unsigned(775, 10), 1987 => to_unsigned(926, 10), 1988 => to_unsigned(340, 10), 1989 => to_unsigned(749, 10), 1990 => to_unsigned(1010, 10), 1991 => to_unsigned(404, 10), 1992 => to_unsigned(118, 10), 1993 => to_unsigned(877, 10), 1994 => to_unsigned(545, 10), 1995 => to_unsigned(1005, 10), 1996 => to_unsigned(518, 10), 1997 => to_unsigned(918, 10), 1998 => to_unsigned(375, 10), 1999 => to_unsigned(467, 10), 2000 => to_unsigned(824, 10), 2001 => to_unsigned(33, 10), 2002 => to_unsigned(278, 10), 2003 => to_unsigned(444, 10), 2004 => to_unsigned(461, 10), 2005 => to_unsigned(383, 10), 2006 => to_unsigned(692, 10), 2007 => to_unsigned(479, 10), 2008 => to_unsigned(468, 10), 2009 => to_unsigned(654, 10), 2010 => to_unsigned(286, 10), 2011 => to_unsigned(16, 10), 2012 => to_unsigned(70, 10), 2013 => to_unsigned(656, 10), 2014 => to_unsigned(33, 10), 2015 => to_unsigned(126, 10), 2016 => to_unsigned(358, 10), 2017 => to_unsigned(635, 10), 2018 => to_unsigned(799, 10), 2019 => to_unsigned(182, 10), 2020 => to_unsigned(337, 10), 2021 => to_unsigned(254, 10), 2022 => to_unsigned(772, 10), 2023 => to_unsigned(353, 10), 2024 => to_unsigned(871, 10), 2025 => to_unsigned(311, 10), 2026 => to_unsigned(207, 10), 2027 => to_unsigned(943, 10), 2028 => to_unsigned(839, 10), 2029 => to_unsigned(61, 10), 2030 => to_unsigned(553, 10), 2031 => to_unsigned(182, 10), 2032 => to_unsigned(820, 10), 2033 => to_unsigned(324, 10), 2034 => to_unsigned(811, 10), 2035 => to_unsigned(702, 10), 2036 => to_unsigned(39, 10), 2037 => to_unsigned(494, 10), 2038 => to_unsigned(864, 10), 2039 => to_unsigned(211, 10), 2040 => to_unsigned(89, 10), 2041 => to_unsigned(719, 10), 2042 => to_unsigned(652, 10), 2043 => to_unsigned(148, 10), 2044 => to_unsigned(892, 10), 2045 => to_unsigned(683, 10), 2046 => to_unsigned(973, 10), 2047 => to_unsigned(397, 10)),
            8 => (0 => to_unsigned(817, 10), 1 => to_unsigned(142, 10), 2 => to_unsigned(192, 10), 3 => to_unsigned(293, 10), 4 => to_unsigned(983, 10), 5 => to_unsigned(549, 10), 6 => to_unsigned(677, 10), 7 => to_unsigned(260, 10), 8 => to_unsigned(605, 10), 9 => to_unsigned(535, 10), 10 => to_unsigned(366, 10), 11 => to_unsigned(873, 10), 12 => to_unsigned(273, 10), 13 => to_unsigned(686, 10), 14 => to_unsigned(578, 10), 15 => to_unsigned(51, 10), 16 => to_unsigned(243, 10), 17 => to_unsigned(523, 10), 18 => to_unsigned(944, 10), 19 => to_unsigned(374, 10), 20 => to_unsigned(767, 10), 21 => to_unsigned(319, 10), 22 => to_unsigned(132, 10), 23 => to_unsigned(6, 10), 24 => to_unsigned(298, 10), 25 => to_unsigned(678, 10), 26 => to_unsigned(72, 10), 27 => to_unsigned(68, 10), 28 => to_unsigned(556, 10), 29 => to_unsigned(559, 10), 30 => to_unsigned(991, 10), 31 => to_unsigned(567, 10), 32 => to_unsigned(688, 10), 33 => to_unsigned(114, 10), 34 => to_unsigned(830, 10), 35 => to_unsigned(217, 10), 36 => to_unsigned(649, 10), 37 => to_unsigned(363, 10), 38 => to_unsigned(317, 10), 39 => to_unsigned(318, 10), 40 => to_unsigned(561, 10), 41 => to_unsigned(304, 10), 42 => to_unsigned(868, 10), 43 => to_unsigned(379, 10), 44 => to_unsigned(526, 10), 45 => to_unsigned(225, 10), 46 => to_unsigned(523, 10), 47 => to_unsigned(401, 10), 48 => to_unsigned(674, 10), 49 => to_unsigned(692, 10), 50 => to_unsigned(446, 10), 51 => to_unsigned(994, 10), 52 => to_unsigned(999, 10), 53 => to_unsigned(15, 10), 54 => to_unsigned(325, 10), 55 => to_unsigned(670, 10), 56 => to_unsigned(728, 10), 57 => to_unsigned(930, 10), 58 => to_unsigned(959, 10), 59 => to_unsigned(701, 10), 60 => to_unsigned(964, 10), 61 => to_unsigned(85, 10), 62 => to_unsigned(612, 10), 63 => to_unsigned(1014, 10), 64 => to_unsigned(929, 10), 65 => to_unsigned(510, 10), 66 => to_unsigned(644, 10), 67 => to_unsigned(150, 10), 68 => to_unsigned(808, 10), 69 => to_unsigned(787, 10), 70 => to_unsigned(928, 10), 71 => to_unsigned(681, 10), 72 => to_unsigned(97, 10), 73 => to_unsigned(403, 10), 74 => to_unsigned(927, 10), 75 => to_unsigned(107, 10), 76 => to_unsigned(410, 10), 77 => to_unsigned(70, 10), 78 => to_unsigned(87, 10), 79 => to_unsigned(207, 10), 80 => to_unsigned(40, 10), 81 => to_unsigned(564, 10), 82 => to_unsigned(69, 10), 83 => to_unsigned(447, 10), 84 => to_unsigned(764, 10), 85 => to_unsigned(890, 10), 86 => to_unsigned(397, 10), 87 => to_unsigned(769, 10), 88 => to_unsigned(323, 10), 89 => to_unsigned(872, 10), 90 => to_unsigned(773, 10), 91 => to_unsigned(932, 10), 92 => to_unsigned(777, 10), 93 => to_unsigned(329, 10), 94 => to_unsigned(300, 10), 95 => to_unsigned(652, 10), 96 => to_unsigned(933, 10), 97 => to_unsigned(933, 10), 98 => to_unsigned(737, 10), 99 => to_unsigned(844, 10), 100 => to_unsigned(664, 10), 101 => to_unsigned(440, 10), 102 => to_unsigned(356, 10), 103 => to_unsigned(305, 10), 104 => to_unsigned(169, 10), 105 => to_unsigned(793, 10), 106 => to_unsigned(116, 10), 107 => to_unsigned(156, 10), 108 => to_unsigned(725, 10), 109 => to_unsigned(738, 10), 110 => to_unsigned(466, 10), 111 => to_unsigned(314, 10), 112 => to_unsigned(565, 10), 113 => to_unsigned(915, 10), 114 => to_unsigned(209, 10), 115 => to_unsigned(181, 10), 116 => to_unsigned(269, 10), 117 => to_unsigned(616, 10), 118 => to_unsigned(401, 10), 119 => to_unsigned(258, 10), 120 => to_unsigned(103, 10), 121 => to_unsigned(861, 10), 122 => to_unsigned(699, 10), 123 => to_unsigned(1003, 10), 124 => to_unsigned(974, 10), 125 => to_unsigned(147, 10), 126 => to_unsigned(805, 10), 127 => to_unsigned(962, 10), 128 => to_unsigned(617, 10), 129 => to_unsigned(73, 10), 130 => to_unsigned(356, 10), 131 => to_unsigned(18, 10), 132 => to_unsigned(480, 10), 133 => to_unsigned(176, 10), 134 => to_unsigned(321, 10), 135 => to_unsigned(529, 10), 136 => to_unsigned(1003, 10), 137 => to_unsigned(825, 10), 138 => to_unsigned(233, 10), 139 => to_unsigned(106, 10), 140 => to_unsigned(824, 10), 141 => to_unsigned(629, 10), 142 => to_unsigned(43, 10), 143 => to_unsigned(585, 10), 144 => to_unsigned(866, 10), 145 => to_unsigned(77, 10), 146 => to_unsigned(618, 10), 147 => to_unsigned(849, 10), 148 => to_unsigned(431, 10), 149 => to_unsigned(687, 10), 150 => to_unsigned(46, 10), 151 => to_unsigned(509, 10), 152 => to_unsigned(698, 10), 153 => to_unsigned(1005, 10), 154 => to_unsigned(693, 10), 155 => to_unsigned(12, 10), 156 => to_unsigned(957, 10), 157 => to_unsigned(946, 10), 158 => to_unsigned(897, 10), 159 => to_unsigned(461, 10), 160 => to_unsigned(284, 10), 161 => to_unsigned(266, 10), 162 => to_unsigned(249, 10), 163 => to_unsigned(278, 10), 164 => to_unsigned(202, 10), 165 => to_unsigned(783, 10), 166 => to_unsigned(66, 10), 167 => to_unsigned(221, 10), 168 => to_unsigned(831, 10), 169 => to_unsigned(27, 10), 170 => to_unsigned(192, 10), 171 => to_unsigned(848, 10), 172 => to_unsigned(480, 10), 173 => to_unsigned(233, 10), 174 => to_unsigned(506, 10), 175 => to_unsigned(666, 10), 176 => to_unsigned(790, 10), 177 => to_unsigned(377, 10), 178 => to_unsigned(448, 10), 179 => to_unsigned(950, 10), 180 => to_unsigned(609, 10), 181 => to_unsigned(659, 10), 182 => to_unsigned(772, 10), 183 => to_unsigned(16, 10), 184 => to_unsigned(736, 10), 185 => to_unsigned(526, 10), 186 => to_unsigned(366, 10), 187 => to_unsigned(716, 10), 188 => to_unsigned(405, 10), 189 => to_unsigned(811, 10), 190 => to_unsigned(29, 10), 191 => to_unsigned(1021, 10), 192 => to_unsigned(409, 10), 193 => to_unsigned(847, 10), 194 => to_unsigned(240, 10), 195 => to_unsigned(29, 10), 196 => to_unsigned(609, 10), 197 => to_unsigned(975, 10), 198 => to_unsigned(160, 10), 199 => to_unsigned(536, 10), 200 => to_unsigned(73, 10), 201 => to_unsigned(732, 10), 202 => to_unsigned(148, 10), 203 => to_unsigned(666, 10), 204 => to_unsigned(708, 10), 205 => to_unsigned(13, 10), 206 => to_unsigned(617, 10), 207 => to_unsigned(788, 10), 208 => to_unsigned(184, 10), 209 => to_unsigned(126, 10), 210 => to_unsigned(1011, 10), 211 => to_unsigned(48, 10), 212 => to_unsigned(744, 10), 213 => to_unsigned(55, 10), 214 => to_unsigned(146, 10), 215 => to_unsigned(359, 10), 216 => to_unsigned(493, 10), 217 => to_unsigned(708, 10), 218 => to_unsigned(934, 10), 219 => to_unsigned(42, 10), 220 => to_unsigned(599, 10), 221 => to_unsigned(398, 10), 222 => to_unsigned(22, 10), 223 => to_unsigned(957, 10), 224 => to_unsigned(8, 10), 225 => to_unsigned(900, 10), 226 => to_unsigned(821, 10), 227 => to_unsigned(599, 10), 228 => to_unsigned(775, 10), 229 => to_unsigned(822, 10), 230 => to_unsigned(919, 10), 231 => to_unsigned(73, 10), 232 => to_unsigned(714, 10), 233 => to_unsigned(610, 10), 234 => to_unsigned(48, 10), 235 => to_unsigned(858, 10), 236 => to_unsigned(565, 10), 237 => to_unsigned(649, 10), 238 => to_unsigned(224, 10), 239 => to_unsigned(34, 10), 240 => to_unsigned(1008, 10), 241 => to_unsigned(329, 10), 242 => to_unsigned(352, 10), 243 => to_unsigned(232, 10), 244 => to_unsigned(830, 10), 245 => to_unsigned(834, 10), 246 => to_unsigned(672, 10), 247 => to_unsigned(431, 10), 248 => to_unsigned(37, 10), 249 => to_unsigned(574, 10), 250 => to_unsigned(835, 10), 251 => to_unsigned(512, 10), 252 => to_unsigned(798, 10), 253 => to_unsigned(460, 10), 254 => to_unsigned(7, 10), 255 => to_unsigned(628, 10), 256 => to_unsigned(551, 10), 257 => to_unsigned(518, 10), 258 => to_unsigned(709, 10), 259 => to_unsigned(426, 10), 260 => to_unsigned(177, 10), 261 => to_unsigned(235, 10), 262 => to_unsigned(823, 10), 263 => to_unsigned(387, 10), 264 => to_unsigned(546, 10), 265 => to_unsigned(452, 10), 266 => to_unsigned(749, 10), 267 => to_unsigned(625, 10), 268 => to_unsigned(558, 10), 269 => to_unsigned(866, 10), 270 => to_unsigned(967, 10), 271 => to_unsigned(300, 10), 272 => to_unsigned(946, 10), 273 => to_unsigned(542, 10), 274 => to_unsigned(1, 10), 275 => to_unsigned(549, 10), 276 => to_unsigned(279, 10), 277 => to_unsigned(950, 10), 278 => to_unsigned(443, 10), 279 => to_unsigned(140, 10), 280 => to_unsigned(131, 10), 281 => to_unsigned(644, 10), 282 => to_unsigned(260, 10), 283 => to_unsigned(483, 10), 284 => to_unsigned(787, 10), 285 => to_unsigned(684, 10), 286 => to_unsigned(510, 10), 287 => to_unsigned(490, 10), 288 => to_unsigned(314, 10), 289 => to_unsigned(583, 10), 290 => to_unsigned(65, 10), 291 => to_unsigned(995, 10), 292 => to_unsigned(516, 10), 293 => to_unsigned(733, 10), 294 => to_unsigned(563, 10), 295 => to_unsigned(51, 10), 296 => to_unsigned(258, 10), 297 => to_unsigned(307, 10), 298 => to_unsigned(837, 10), 299 => to_unsigned(242, 10), 300 => to_unsigned(392, 10), 301 => to_unsigned(502, 10), 302 => to_unsigned(314, 10), 303 => to_unsigned(990, 10), 304 => to_unsigned(165, 10), 305 => to_unsigned(704, 10), 306 => to_unsigned(679, 10), 307 => to_unsigned(239, 10), 308 => to_unsigned(542, 10), 309 => to_unsigned(570, 10), 310 => to_unsigned(228, 10), 311 => to_unsigned(604, 10), 312 => to_unsigned(709, 10), 313 => to_unsigned(1019, 10), 314 => to_unsigned(961, 10), 315 => to_unsigned(428, 10), 316 => to_unsigned(388, 10), 317 => to_unsigned(148, 10), 318 => to_unsigned(258, 10), 319 => to_unsigned(257, 10), 320 => to_unsigned(13, 10), 321 => to_unsigned(549, 10), 322 => to_unsigned(854, 10), 323 => to_unsigned(683, 10), 324 => to_unsigned(96, 10), 325 => to_unsigned(667, 10), 326 => to_unsigned(846, 10), 327 => to_unsigned(650, 10), 328 => to_unsigned(220, 10), 329 => to_unsigned(287, 10), 330 => to_unsigned(340, 10), 331 => to_unsigned(383, 10), 332 => to_unsigned(441, 10), 333 => to_unsigned(628, 10), 334 => to_unsigned(76, 10), 335 => to_unsigned(202, 10), 336 => to_unsigned(1008, 10), 337 => to_unsigned(919, 10), 338 => to_unsigned(645, 10), 339 => to_unsigned(789, 10), 340 => to_unsigned(432, 10), 341 => to_unsigned(807, 10), 342 => to_unsigned(595, 10), 343 => to_unsigned(922, 10), 344 => to_unsigned(619, 10), 345 => to_unsigned(244, 10), 346 => to_unsigned(496, 10), 347 => to_unsigned(539, 10), 348 => to_unsigned(731, 10), 349 => to_unsigned(241, 10), 350 => to_unsigned(55, 10), 351 => to_unsigned(397, 10), 352 => to_unsigned(135, 10), 353 => to_unsigned(970, 10), 354 => to_unsigned(408, 10), 355 => to_unsigned(719, 10), 356 => to_unsigned(938, 10), 357 => to_unsigned(235, 10), 358 => to_unsigned(735, 10), 359 => to_unsigned(821, 10), 360 => to_unsigned(527, 10), 361 => to_unsigned(329, 10), 362 => to_unsigned(675, 10), 363 => to_unsigned(428, 10), 364 => to_unsigned(291, 10), 365 => to_unsigned(57, 10), 366 => to_unsigned(98, 10), 367 => to_unsigned(289, 10), 368 => to_unsigned(913, 10), 369 => to_unsigned(78, 10), 370 => to_unsigned(278, 10), 371 => to_unsigned(11, 10), 372 => to_unsigned(410, 10), 373 => to_unsigned(987, 10), 374 => to_unsigned(483, 10), 375 => to_unsigned(229, 10), 376 => to_unsigned(751, 10), 377 => to_unsigned(821, 10), 378 => to_unsigned(558, 10), 379 => to_unsigned(683, 10), 380 => to_unsigned(540, 10), 381 => to_unsigned(250, 10), 382 => to_unsigned(639, 10), 383 => to_unsigned(229, 10), 384 => to_unsigned(368, 10), 385 => to_unsigned(30, 10), 386 => to_unsigned(687, 10), 387 => to_unsigned(255, 10), 388 => to_unsigned(837, 10), 389 => to_unsigned(41, 10), 390 => to_unsigned(362, 10), 391 => to_unsigned(518, 10), 392 => to_unsigned(804, 10), 393 => to_unsigned(587, 10), 394 => to_unsigned(997, 10), 395 => to_unsigned(561, 10), 396 => to_unsigned(83, 10), 397 => to_unsigned(352, 10), 398 => to_unsigned(122, 10), 399 => to_unsigned(396, 10), 400 => to_unsigned(453, 10), 401 => to_unsigned(415, 10), 402 => to_unsigned(377, 10), 403 => to_unsigned(794, 10), 404 => to_unsigned(961, 10), 405 => to_unsigned(813, 10), 406 => to_unsigned(539, 10), 407 => to_unsigned(384, 10), 408 => to_unsigned(632, 10), 409 => to_unsigned(412, 10), 410 => to_unsigned(667, 10), 411 => to_unsigned(308, 10), 412 => to_unsigned(565, 10), 413 => to_unsigned(487, 10), 414 => to_unsigned(763, 10), 415 => to_unsigned(195, 10), 416 => to_unsigned(935, 10), 417 => to_unsigned(649, 10), 418 => to_unsigned(234, 10), 419 => to_unsigned(1000, 10), 420 => to_unsigned(252, 10), 421 => to_unsigned(693, 10), 422 => to_unsigned(21, 10), 423 => to_unsigned(143, 10), 424 => to_unsigned(437, 10), 425 => to_unsigned(620, 10), 426 => to_unsigned(477, 10), 427 => to_unsigned(830, 10), 428 => to_unsigned(205, 10), 429 => to_unsigned(677, 10), 430 => to_unsigned(90, 10), 431 => to_unsigned(880, 10), 432 => to_unsigned(520, 10), 433 => to_unsigned(276, 10), 434 => to_unsigned(567, 10), 435 => to_unsigned(491, 10), 436 => to_unsigned(883, 10), 437 => to_unsigned(389, 10), 438 => to_unsigned(64, 10), 439 => to_unsigned(184, 10), 440 => to_unsigned(712, 10), 441 => to_unsigned(875, 10), 442 => to_unsigned(622, 10), 443 => to_unsigned(418, 10), 444 => to_unsigned(234, 10), 445 => to_unsigned(739, 10), 446 => to_unsigned(952, 10), 447 => to_unsigned(793, 10), 448 => to_unsigned(352, 10), 449 => to_unsigned(947, 10), 450 => to_unsigned(342, 10), 451 => to_unsigned(99, 10), 452 => to_unsigned(953, 10), 453 => to_unsigned(749, 10), 454 => to_unsigned(442, 10), 455 => to_unsigned(454, 10), 456 => to_unsigned(929, 10), 457 => to_unsigned(502, 10), 458 => to_unsigned(894, 10), 459 => to_unsigned(592, 10), 460 => to_unsigned(29, 10), 461 => to_unsigned(270, 10), 462 => to_unsigned(599, 10), 463 => to_unsigned(456, 10), 464 => to_unsigned(127, 10), 465 => to_unsigned(902, 10), 466 => to_unsigned(319, 10), 467 => to_unsigned(72, 10), 468 => to_unsigned(492, 10), 469 => to_unsigned(441, 10), 470 => to_unsigned(24, 10), 471 => to_unsigned(199, 10), 472 => to_unsigned(851, 10), 473 => to_unsigned(394, 10), 474 => to_unsigned(861, 10), 475 => to_unsigned(688, 10), 476 => to_unsigned(835, 10), 477 => to_unsigned(149, 10), 478 => to_unsigned(636, 10), 479 => to_unsigned(237, 10), 480 => to_unsigned(532, 10), 481 => to_unsigned(503, 10), 482 => to_unsigned(459, 10), 483 => to_unsigned(535, 10), 484 => to_unsigned(883, 10), 485 => to_unsigned(100, 10), 486 => to_unsigned(304, 10), 487 => to_unsigned(900, 10), 488 => to_unsigned(600, 10), 489 => to_unsigned(907, 10), 490 => to_unsigned(367, 10), 491 => to_unsigned(970, 10), 492 => to_unsigned(180, 10), 493 => to_unsigned(799, 10), 494 => to_unsigned(814, 10), 495 => to_unsigned(342, 10), 496 => to_unsigned(854, 10), 497 => to_unsigned(673, 10), 498 => to_unsigned(462, 10), 499 => to_unsigned(651, 10), 500 => to_unsigned(93, 10), 501 => to_unsigned(468, 10), 502 => to_unsigned(452, 10), 503 => to_unsigned(630, 10), 504 => to_unsigned(54, 10), 505 => to_unsigned(1000, 10), 506 => to_unsigned(452, 10), 507 => to_unsigned(707, 10), 508 => to_unsigned(437, 10), 509 => to_unsigned(931, 10), 510 => to_unsigned(411, 10), 511 => to_unsigned(219, 10), 512 => to_unsigned(403, 10), 513 => to_unsigned(140, 10), 514 => to_unsigned(74, 10), 515 => to_unsigned(26, 10), 516 => to_unsigned(612, 10), 517 => to_unsigned(871, 10), 518 => to_unsigned(872, 10), 519 => to_unsigned(198, 10), 520 => to_unsigned(405, 10), 521 => to_unsigned(999, 10), 522 => to_unsigned(623, 10), 523 => to_unsigned(29, 10), 524 => to_unsigned(806, 10), 525 => to_unsigned(121, 10), 526 => to_unsigned(436, 10), 527 => to_unsigned(625, 10), 528 => to_unsigned(142, 10), 529 => to_unsigned(331, 10), 530 => to_unsigned(451, 10), 531 => to_unsigned(318, 10), 532 => to_unsigned(128, 10), 533 => to_unsigned(38, 10), 534 => to_unsigned(991, 10), 535 => to_unsigned(42, 10), 536 => to_unsigned(642, 10), 537 => to_unsigned(804, 10), 538 => to_unsigned(110, 10), 539 => to_unsigned(385, 10), 540 => to_unsigned(846, 10), 541 => to_unsigned(713, 10), 542 => to_unsigned(49, 10), 543 => to_unsigned(88, 10), 544 => to_unsigned(317, 10), 545 => to_unsigned(864, 10), 546 => to_unsigned(12, 10), 547 => to_unsigned(403, 10), 548 => to_unsigned(752, 10), 549 => to_unsigned(198, 10), 550 => to_unsigned(534, 10), 551 => to_unsigned(75, 10), 552 => to_unsigned(682, 10), 553 => to_unsigned(977, 10), 554 => to_unsigned(454, 10), 555 => to_unsigned(488, 10), 556 => to_unsigned(458, 10), 557 => to_unsigned(514, 10), 558 => to_unsigned(80, 10), 559 => to_unsigned(351, 10), 560 => to_unsigned(263, 10), 561 => to_unsigned(973, 10), 562 => to_unsigned(789, 10), 563 => to_unsigned(603, 10), 564 => to_unsigned(49, 10), 565 => to_unsigned(333, 10), 566 => to_unsigned(137, 10), 567 => to_unsigned(955, 10), 568 => to_unsigned(425, 10), 569 => to_unsigned(382, 10), 570 => to_unsigned(222, 10), 571 => to_unsigned(585, 10), 572 => to_unsigned(62, 10), 573 => to_unsigned(811, 10), 574 => to_unsigned(803, 10), 575 => to_unsigned(118, 10), 576 => to_unsigned(373, 10), 577 => to_unsigned(10, 10), 578 => to_unsigned(629, 10), 579 => to_unsigned(296, 10), 580 => to_unsigned(73, 10), 581 => to_unsigned(58, 10), 582 => to_unsigned(995, 10), 583 => to_unsigned(752, 10), 584 => to_unsigned(484, 10), 585 => to_unsigned(280, 10), 586 => to_unsigned(812, 10), 587 => to_unsigned(815, 10), 588 => to_unsigned(838, 10), 589 => to_unsigned(39, 10), 590 => to_unsigned(387, 10), 591 => to_unsigned(1002, 10), 592 => to_unsigned(246, 10), 593 => to_unsigned(387, 10), 594 => to_unsigned(9, 10), 595 => to_unsigned(34, 10), 596 => to_unsigned(615, 10), 597 => to_unsigned(173, 10), 598 => to_unsigned(45, 10), 599 => to_unsigned(737, 10), 600 => to_unsigned(36, 10), 601 => to_unsigned(818, 10), 602 => to_unsigned(144, 10), 603 => to_unsigned(633, 10), 604 => to_unsigned(806, 10), 605 => to_unsigned(555, 10), 606 => to_unsigned(617, 10), 607 => to_unsigned(742, 10), 608 => to_unsigned(103, 10), 609 => to_unsigned(288, 10), 610 => to_unsigned(245, 10), 611 => to_unsigned(297, 10), 612 => to_unsigned(418, 10), 613 => to_unsigned(44, 10), 614 => to_unsigned(491, 10), 615 => to_unsigned(280, 10), 616 => to_unsigned(942, 10), 617 => to_unsigned(662, 10), 618 => to_unsigned(714, 10), 619 => to_unsigned(144, 10), 620 => to_unsigned(97, 10), 621 => to_unsigned(630, 10), 622 => to_unsigned(172, 10), 623 => to_unsigned(302, 10), 624 => to_unsigned(245, 10), 625 => to_unsigned(729, 10), 626 => to_unsigned(0, 10), 627 => to_unsigned(885, 10), 628 => to_unsigned(480, 10), 629 => to_unsigned(884, 10), 630 => to_unsigned(858, 10), 631 => to_unsigned(63, 10), 632 => to_unsigned(220, 10), 633 => to_unsigned(950, 10), 634 => to_unsigned(789, 10), 635 => to_unsigned(928, 10), 636 => to_unsigned(559, 10), 637 => to_unsigned(752, 10), 638 => to_unsigned(995, 10), 639 => to_unsigned(750, 10), 640 => to_unsigned(628, 10), 641 => to_unsigned(659, 10), 642 => to_unsigned(120, 10), 643 => to_unsigned(963, 10), 644 => to_unsigned(272, 10), 645 => to_unsigned(354, 10), 646 => to_unsigned(497, 10), 647 => to_unsigned(386, 10), 648 => to_unsigned(305, 10), 649 => to_unsigned(682, 10), 650 => to_unsigned(974, 10), 651 => to_unsigned(888, 10), 652 => to_unsigned(227, 10), 653 => to_unsigned(176, 10), 654 => to_unsigned(643, 10), 655 => to_unsigned(618, 10), 656 => to_unsigned(123, 10), 657 => to_unsigned(829, 10), 658 => to_unsigned(529, 10), 659 => to_unsigned(791, 10), 660 => to_unsigned(998, 10), 661 => to_unsigned(655, 10), 662 => to_unsigned(798, 10), 663 => to_unsigned(869, 10), 664 => to_unsigned(891, 10), 665 => to_unsigned(165, 10), 666 => to_unsigned(115, 10), 667 => to_unsigned(425, 10), 668 => to_unsigned(200, 10), 669 => to_unsigned(1003, 10), 670 => to_unsigned(979, 10), 671 => to_unsigned(221, 10), 672 => to_unsigned(333, 10), 673 => to_unsigned(444, 10), 674 => to_unsigned(984, 10), 675 => to_unsigned(821, 10), 676 => to_unsigned(29, 10), 677 => to_unsigned(382, 10), 678 => to_unsigned(330, 10), 679 => to_unsigned(471, 10), 680 => to_unsigned(456, 10), 681 => to_unsigned(263, 10), 682 => to_unsigned(647, 10), 683 => to_unsigned(976, 10), 684 => to_unsigned(924, 10), 685 => to_unsigned(609, 10), 686 => to_unsigned(17, 10), 687 => to_unsigned(792, 10), 688 => to_unsigned(64, 10), 689 => to_unsigned(930, 10), 690 => to_unsigned(159, 10), 691 => to_unsigned(188, 10), 692 => to_unsigned(735, 10), 693 => to_unsigned(586, 10), 694 => to_unsigned(855, 10), 695 => to_unsigned(629, 10), 696 => to_unsigned(812, 10), 697 => to_unsigned(535, 10), 698 => to_unsigned(585, 10), 699 => to_unsigned(589, 10), 700 => to_unsigned(624, 10), 701 => to_unsigned(261, 10), 702 => to_unsigned(297, 10), 703 => to_unsigned(782, 10), 704 => to_unsigned(394, 10), 705 => to_unsigned(692, 10), 706 => to_unsigned(925, 10), 707 => to_unsigned(630, 10), 708 => to_unsigned(987, 10), 709 => to_unsigned(548, 10), 710 => to_unsigned(527, 10), 711 => to_unsigned(977, 10), 712 => to_unsigned(1017, 10), 713 => to_unsigned(40, 10), 714 => to_unsigned(156, 10), 715 => to_unsigned(3, 10), 716 => to_unsigned(287, 10), 717 => to_unsigned(54, 10), 718 => to_unsigned(754, 10), 719 => to_unsigned(614, 10), 720 => to_unsigned(803, 10), 721 => to_unsigned(169, 10), 722 => to_unsigned(298, 10), 723 => to_unsigned(557, 10), 724 => to_unsigned(274, 10), 725 => to_unsigned(833, 10), 726 => to_unsigned(114, 10), 727 => to_unsigned(621, 10), 728 => to_unsigned(509, 10), 729 => to_unsigned(995, 10), 730 => to_unsigned(241, 10), 731 => to_unsigned(297, 10), 732 => to_unsigned(375, 10), 733 => to_unsigned(114, 10), 734 => to_unsigned(903, 10), 735 => to_unsigned(274, 10), 736 => to_unsigned(356, 10), 737 => to_unsigned(990, 10), 738 => to_unsigned(856, 10), 739 => to_unsigned(29, 10), 740 => to_unsigned(164, 10), 741 => to_unsigned(310, 10), 742 => to_unsigned(556, 10), 743 => to_unsigned(177, 10), 744 => to_unsigned(576, 10), 745 => to_unsigned(214, 10), 746 => to_unsigned(846, 10), 747 => to_unsigned(214, 10), 748 => to_unsigned(912, 10), 749 => to_unsigned(504, 10), 750 => to_unsigned(26, 10), 751 => to_unsigned(38, 10), 752 => to_unsigned(171, 10), 753 => to_unsigned(804, 10), 754 => to_unsigned(203, 10), 755 => to_unsigned(54, 10), 756 => to_unsigned(488, 10), 757 => to_unsigned(899, 10), 758 => to_unsigned(700, 10), 759 => to_unsigned(276, 10), 760 => to_unsigned(185, 10), 761 => to_unsigned(506, 10), 762 => to_unsigned(523, 10), 763 => to_unsigned(941, 10), 764 => to_unsigned(705, 10), 765 => to_unsigned(870, 10), 766 => to_unsigned(346, 10), 767 => to_unsigned(145, 10), 768 => to_unsigned(4, 10), 769 => to_unsigned(628, 10), 770 => to_unsigned(420, 10), 771 => to_unsigned(951, 10), 772 => to_unsigned(132, 10), 773 => to_unsigned(534, 10), 774 => to_unsigned(68, 10), 775 => to_unsigned(592, 10), 776 => to_unsigned(72, 10), 777 => to_unsigned(759, 10), 778 => to_unsigned(256, 10), 779 => to_unsigned(519, 10), 780 => to_unsigned(655, 10), 781 => to_unsigned(384, 10), 782 => to_unsigned(678, 10), 783 => to_unsigned(660, 10), 784 => to_unsigned(997, 10), 785 => to_unsigned(795, 10), 786 => to_unsigned(501, 10), 787 => to_unsigned(789, 10), 788 => to_unsigned(846, 10), 789 => to_unsigned(312, 10), 790 => to_unsigned(868, 10), 791 => to_unsigned(268, 10), 792 => to_unsigned(263, 10), 793 => to_unsigned(751, 10), 794 => to_unsigned(758, 10), 795 => to_unsigned(876, 10), 796 => to_unsigned(292, 10), 797 => to_unsigned(855, 10), 798 => to_unsigned(891, 10), 799 => to_unsigned(419, 10), 800 => to_unsigned(341, 10), 801 => to_unsigned(795, 10), 802 => to_unsigned(247, 10), 803 => to_unsigned(210, 10), 804 => to_unsigned(75, 10), 805 => to_unsigned(253, 10), 806 => to_unsigned(82, 10), 807 => to_unsigned(46, 10), 808 => to_unsigned(220, 10), 809 => to_unsigned(507, 10), 810 => to_unsigned(452, 10), 811 => to_unsigned(413, 10), 812 => to_unsigned(924, 10), 813 => to_unsigned(259, 10), 814 => to_unsigned(872, 10), 815 => to_unsigned(256, 10), 816 => to_unsigned(136, 10), 817 => to_unsigned(268, 10), 818 => to_unsigned(404, 10), 819 => to_unsigned(628, 10), 820 => to_unsigned(234, 10), 821 => to_unsigned(767, 10), 822 => to_unsigned(338, 10), 823 => to_unsigned(597, 10), 824 => to_unsigned(78, 10), 825 => to_unsigned(545, 10), 826 => to_unsigned(631, 10), 827 => to_unsigned(280, 10), 828 => to_unsigned(733, 10), 829 => to_unsigned(137, 10), 830 => to_unsigned(169, 10), 831 => to_unsigned(531, 10), 832 => to_unsigned(372, 10), 833 => to_unsigned(983, 10), 834 => to_unsigned(234, 10), 835 => to_unsigned(207, 10), 836 => to_unsigned(851, 10), 837 => to_unsigned(336, 10), 838 => to_unsigned(577, 10), 839 => to_unsigned(701, 10), 840 => to_unsigned(215, 10), 841 => to_unsigned(123, 10), 842 => to_unsigned(413, 10), 843 => to_unsigned(559, 10), 844 => to_unsigned(3, 10), 845 => to_unsigned(242, 10), 846 => to_unsigned(492, 10), 847 => to_unsigned(462, 10), 848 => to_unsigned(662, 10), 849 => to_unsigned(567, 10), 850 => to_unsigned(693, 10), 851 => to_unsigned(475, 10), 852 => to_unsigned(562, 10), 853 => to_unsigned(491, 10), 854 => to_unsigned(664, 10), 855 => to_unsigned(348, 10), 856 => to_unsigned(979, 10), 857 => to_unsigned(223, 10), 858 => to_unsigned(537, 10), 859 => to_unsigned(186, 10), 860 => to_unsigned(882, 10), 861 => to_unsigned(386, 10), 862 => to_unsigned(413, 10), 863 => to_unsigned(817, 10), 864 => to_unsigned(563, 10), 865 => to_unsigned(725, 10), 866 => to_unsigned(308, 10), 867 => to_unsigned(20, 10), 868 => to_unsigned(19, 10), 869 => to_unsigned(994, 10), 870 => to_unsigned(854, 10), 871 => to_unsigned(903, 10), 872 => to_unsigned(564, 10), 873 => to_unsigned(217, 10), 874 => to_unsigned(10, 10), 875 => to_unsigned(692, 10), 876 => to_unsigned(432, 10), 877 => to_unsigned(370, 10), 878 => to_unsigned(999, 10), 879 => to_unsigned(126, 10), 880 => to_unsigned(854, 10), 881 => to_unsigned(530, 10), 882 => to_unsigned(151, 10), 883 => to_unsigned(850, 10), 884 => to_unsigned(470, 10), 885 => to_unsigned(884, 10), 886 => to_unsigned(868, 10), 887 => to_unsigned(436, 10), 888 => to_unsigned(635, 10), 889 => to_unsigned(871, 10), 890 => to_unsigned(256, 10), 891 => to_unsigned(828, 10), 892 => to_unsigned(220, 10), 893 => to_unsigned(260, 10), 894 => to_unsigned(890, 10), 895 => to_unsigned(810, 10), 896 => to_unsigned(82, 10), 897 => to_unsigned(70, 10), 898 => to_unsigned(892, 10), 899 => to_unsigned(929, 10), 900 => to_unsigned(614, 10), 901 => to_unsigned(36, 10), 902 => to_unsigned(349, 10), 903 => to_unsigned(758, 10), 904 => to_unsigned(812, 10), 905 => to_unsigned(882, 10), 906 => to_unsigned(359, 10), 907 => to_unsigned(56, 10), 908 => to_unsigned(896, 10), 909 => to_unsigned(1016, 10), 910 => to_unsigned(688, 10), 911 => to_unsigned(877, 10), 912 => to_unsigned(536, 10), 913 => to_unsigned(793, 10), 914 => to_unsigned(817, 10), 915 => to_unsigned(917, 10), 916 => to_unsigned(316, 10), 917 => to_unsigned(129, 10), 918 => to_unsigned(608, 10), 919 => to_unsigned(62, 10), 920 => to_unsigned(828, 10), 921 => to_unsigned(904, 10), 922 => to_unsigned(633, 10), 923 => to_unsigned(253, 10), 924 => to_unsigned(8, 10), 925 => to_unsigned(699, 10), 926 => to_unsigned(887, 10), 927 => to_unsigned(288, 10), 928 => to_unsigned(223, 10), 929 => to_unsigned(56, 10), 930 => to_unsigned(855, 10), 931 => to_unsigned(279, 10), 932 => to_unsigned(441, 10), 933 => to_unsigned(399, 10), 934 => to_unsigned(511, 10), 935 => to_unsigned(166, 10), 936 => to_unsigned(549, 10), 937 => to_unsigned(310, 10), 938 => to_unsigned(480, 10), 939 => to_unsigned(822, 10), 940 => to_unsigned(96, 10), 941 => to_unsigned(681, 10), 942 => to_unsigned(110, 10), 943 => to_unsigned(285, 10), 944 => to_unsigned(380, 10), 945 => to_unsigned(557, 10), 946 => to_unsigned(255, 10), 947 => to_unsigned(897, 10), 948 => to_unsigned(671, 10), 949 => to_unsigned(638, 10), 950 => to_unsigned(798, 10), 951 => to_unsigned(217, 10), 952 => to_unsigned(547, 10), 953 => to_unsigned(786, 10), 954 => to_unsigned(31, 10), 955 => to_unsigned(708, 10), 956 => to_unsigned(6, 10), 957 => to_unsigned(969, 10), 958 => to_unsigned(114, 10), 959 => to_unsigned(711, 10), 960 => to_unsigned(133, 10), 961 => to_unsigned(939, 10), 962 => to_unsigned(702, 10), 963 => to_unsigned(633, 10), 964 => to_unsigned(354, 10), 965 => to_unsigned(731, 10), 966 => to_unsigned(969, 10), 967 => to_unsigned(739, 10), 968 => to_unsigned(176, 10), 969 => to_unsigned(238, 10), 970 => to_unsigned(598, 10), 971 => to_unsigned(356, 10), 972 => to_unsigned(375, 10), 973 => to_unsigned(515, 10), 974 => to_unsigned(467, 10), 975 => to_unsigned(187, 10), 976 => to_unsigned(276, 10), 977 => to_unsigned(912, 10), 978 => to_unsigned(293, 10), 979 => to_unsigned(685, 10), 980 => to_unsigned(259, 10), 981 => to_unsigned(895, 10), 982 => to_unsigned(536, 10), 983 => to_unsigned(876, 10), 984 => to_unsigned(575, 10), 985 => to_unsigned(288, 10), 986 => to_unsigned(72, 10), 987 => to_unsigned(853, 10), 988 => to_unsigned(792, 10), 989 => to_unsigned(964, 10), 990 => to_unsigned(7, 10), 991 => to_unsigned(924, 10), 992 => to_unsigned(359, 10), 993 => to_unsigned(49, 10), 994 => to_unsigned(478, 10), 995 => to_unsigned(610, 10), 996 => to_unsigned(230, 10), 997 => to_unsigned(612, 10), 998 => to_unsigned(448, 10), 999 => to_unsigned(835, 10), 1000 => to_unsigned(94, 10), 1001 => to_unsigned(613, 10), 1002 => to_unsigned(691, 10), 1003 => to_unsigned(818, 10), 1004 => to_unsigned(188, 10), 1005 => to_unsigned(970, 10), 1006 => to_unsigned(570, 10), 1007 => to_unsigned(464, 10), 1008 => to_unsigned(852, 10), 1009 => to_unsigned(652, 10), 1010 => to_unsigned(1022, 10), 1011 => to_unsigned(648, 10), 1012 => to_unsigned(579, 10), 1013 => to_unsigned(611, 10), 1014 => to_unsigned(635, 10), 1015 => to_unsigned(501, 10), 1016 => to_unsigned(425, 10), 1017 => to_unsigned(348, 10), 1018 => to_unsigned(801, 10), 1019 => to_unsigned(264, 10), 1020 => to_unsigned(227, 10), 1021 => to_unsigned(44, 10), 1022 => to_unsigned(272, 10), 1023 => to_unsigned(904, 10), 1024 => to_unsigned(13, 10), 1025 => to_unsigned(820, 10), 1026 => to_unsigned(650, 10), 1027 => to_unsigned(114, 10), 1028 => to_unsigned(374, 10), 1029 => to_unsigned(496, 10), 1030 => to_unsigned(192, 10), 1031 => to_unsigned(698, 10), 1032 => to_unsigned(16, 10), 1033 => to_unsigned(679, 10), 1034 => to_unsigned(972, 10), 1035 => to_unsigned(29, 10), 1036 => to_unsigned(20, 10), 1037 => to_unsigned(628, 10), 1038 => to_unsigned(416, 10), 1039 => to_unsigned(635, 10), 1040 => to_unsigned(87, 10), 1041 => to_unsigned(522, 10), 1042 => to_unsigned(18, 10), 1043 => to_unsigned(395, 10), 1044 => to_unsigned(42, 10), 1045 => to_unsigned(267, 10), 1046 => to_unsigned(455, 10), 1047 => to_unsigned(966, 10), 1048 => to_unsigned(407, 10), 1049 => to_unsigned(887, 10), 1050 => to_unsigned(192, 10), 1051 => to_unsigned(608, 10), 1052 => to_unsigned(392, 10), 1053 => to_unsigned(54, 10), 1054 => to_unsigned(387, 10), 1055 => to_unsigned(646, 10), 1056 => to_unsigned(622, 10), 1057 => to_unsigned(146, 10), 1058 => to_unsigned(452, 10), 1059 => to_unsigned(336, 10), 1060 => to_unsigned(476, 10), 1061 => to_unsigned(819, 10), 1062 => to_unsigned(72, 10), 1063 => to_unsigned(858, 10), 1064 => to_unsigned(179, 10), 1065 => to_unsigned(627, 10), 1066 => to_unsigned(132, 10), 1067 => to_unsigned(109, 10), 1068 => to_unsigned(243, 10), 1069 => to_unsigned(155, 10), 1070 => to_unsigned(768, 10), 1071 => to_unsigned(796, 10), 1072 => to_unsigned(606, 10), 1073 => to_unsigned(798, 10), 1074 => to_unsigned(45, 10), 1075 => to_unsigned(584, 10), 1076 => to_unsigned(60, 10), 1077 => to_unsigned(657, 10), 1078 => to_unsigned(210, 10), 1079 => to_unsigned(50, 10), 1080 => to_unsigned(250, 10), 1081 => to_unsigned(94, 10), 1082 => to_unsigned(974, 10), 1083 => to_unsigned(559, 10), 1084 => to_unsigned(534, 10), 1085 => to_unsigned(143, 10), 1086 => to_unsigned(983, 10), 1087 => to_unsigned(894, 10), 1088 => to_unsigned(539, 10), 1089 => to_unsigned(801, 10), 1090 => to_unsigned(245, 10), 1091 => to_unsigned(702, 10), 1092 => to_unsigned(965, 10), 1093 => to_unsigned(472, 10), 1094 => to_unsigned(956, 10), 1095 => to_unsigned(335, 10), 1096 => to_unsigned(315, 10), 1097 => to_unsigned(375, 10), 1098 => to_unsigned(130, 10), 1099 => to_unsigned(650, 10), 1100 => to_unsigned(142, 10), 1101 => to_unsigned(128, 10), 1102 => to_unsigned(487, 10), 1103 => to_unsigned(423, 10), 1104 => to_unsigned(15, 10), 1105 => to_unsigned(850, 10), 1106 => to_unsigned(240, 10), 1107 => to_unsigned(799, 10), 1108 => to_unsigned(713, 10), 1109 => to_unsigned(1001, 10), 1110 => to_unsigned(377, 10), 1111 => to_unsigned(810, 10), 1112 => to_unsigned(463, 10), 1113 => to_unsigned(633, 10), 1114 => to_unsigned(103, 10), 1115 => to_unsigned(888, 10), 1116 => to_unsigned(612, 10), 1117 => to_unsigned(835, 10), 1118 => to_unsigned(923, 10), 1119 => to_unsigned(944, 10), 1120 => to_unsigned(789, 10), 1121 => to_unsigned(164, 10), 1122 => to_unsigned(916, 10), 1123 => to_unsigned(871, 10), 1124 => to_unsigned(991, 10), 1125 => to_unsigned(1009, 10), 1126 => to_unsigned(395, 10), 1127 => to_unsigned(1018, 10), 1128 => to_unsigned(664, 10), 1129 => to_unsigned(977, 10), 1130 => to_unsigned(332, 10), 1131 => to_unsigned(962, 10), 1132 => to_unsigned(634, 10), 1133 => to_unsigned(193, 10), 1134 => to_unsigned(506, 10), 1135 => to_unsigned(913, 10), 1136 => to_unsigned(625, 10), 1137 => to_unsigned(588, 10), 1138 => to_unsigned(421, 10), 1139 => to_unsigned(436, 10), 1140 => to_unsigned(691, 10), 1141 => to_unsigned(46, 10), 1142 => to_unsigned(492, 10), 1143 => to_unsigned(101, 10), 1144 => to_unsigned(555, 10), 1145 => to_unsigned(772, 10), 1146 => to_unsigned(419, 10), 1147 => to_unsigned(175, 10), 1148 => to_unsigned(702, 10), 1149 => to_unsigned(534, 10), 1150 => to_unsigned(863, 10), 1151 => to_unsigned(384, 10), 1152 => to_unsigned(434, 10), 1153 => to_unsigned(456, 10), 1154 => to_unsigned(796, 10), 1155 => to_unsigned(312, 10), 1156 => to_unsigned(1009, 10), 1157 => to_unsigned(235, 10), 1158 => to_unsigned(503, 10), 1159 => to_unsigned(698, 10), 1160 => to_unsigned(781, 10), 1161 => to_unsigned(946, 10), 1162 => to_unsigned(364, 10), 1163 => to_unsigned(835, 10), 1164 => to_unsigned(632, 10), 1165 => to_unsigned(501, 10), 1166 => to_unsigned(807, 10), 1167 => to_unsigned(356, 10), 1168 => to_unsigned(697, 10), 1169 => to_unsigned(182, 10), 1170 => to_unsigned(263, 10), 1171 => to_unsigned(643, 10), 1172 => to_unsigned(566, 10), 1173 => to_unsigned(683, 10), 1174 => to_unsigned(1000, 10), 1175 => to_unsigned(70, 10), 1176 => to_unsigned(448, 10), 1177 => to_unsigned(662, 10), 1178 => to_unsigned(97, 10), 1179 => to_unsigned(222, 10), 1180 => to_unsigned(968, 10), 1181 => to_unsigned(462, 10), 1182 => to_unsigned(208, 10), 1183 => to_unsigned(974, 10), 1184 => to_unsigned(306, 10), 1185 => to_unsigned(897, 10), 1186 => to_unsigned(574, 10), 1187 => to_unsigned(387, 10), 1188 => to_unsigned(919, 10), 1189 => to_unsigned(26, 10), 1190 => to_unsigned(817, 10), 1191 => to_unsigned(791, 10), 1192 => to_unsigned(650, 10), 1193 => to_unsigned(783, 10), 1194 => to_unsigned(961, 10), 1195 => to_unsigned(508, 10), 1196 => to_unsigned(212, 10), 1197 => to_unsigned(215, 10), 1198 => to_unsigned(534, 10), 1199 => to_unsigned(1003, 10), 1200 => to_unsigned(1012, 10), 1201 => to_unsigned(142, 10), 1202 => to_unsigned(401, 10), 1203 => to_unsigned(942, 10), 1204 => to_unsigned(495, 10), 1205 => to_unsigned(589, 10), 1206 => to_unsigned(944, 10), 1207 => to_unsigned(701, 10), 1208 => to_unsigned(465, 10), 1209 => to_unsigned(433, 10), 1210 => to_unsigned(413, 10), 1211 => to_unsigned(124, 10), 1212 => to_unsigned(323, 10), 1213 => to_unsigned(140, 10), 1214 => to_unsigned(920, 10), 1215 => to_unsigned(536, 10), 1216 => to_unsigned(702, 10), 1217 => to_unsigned(933, 10), 1218 => to_unsigned(587, 10), 1219 => to_unsigned(357, 10), 1220 => to_unsigned(10, 10), 1221 => to_unsigned(198, 10), 1222 => to_unsigned(428, 10), 1223 => to_unsigned(898, 10), 1224 => to_unsigned(411, 10), 1225 => to_unsigned(569, 10), 1226 => to_unsigned(726, 10), 1227 => to_unsigned(125, 10), 1228 => to_unsigned(1009, 10), 1229 => to_unsigned(76, 10), 1230 => to_unsigned(127, 10), 1231 => to_unsigned(773, 10), 1232 => to_unsigned(655, 10), 1233 => to_unsigned(406, 10), 1234 => to_unsigned(61, 10), 1235 => to_unsigned(561, 10), 1236 => to_unsigned(690, 10), 1237 => to_unsigned(160, 10), 1238 => to_unsigned(338, 10), 1239 => to_unsigned(335, 10), 1240 => to_unsigned(178, 10), 1241 => to_unsigned(152, 10), 1242 => to_unsigned(57, 10), 1243 => to_unsigned(898, 10), 1244 => to_unsigned(148, 10), 1245 => to_unsigned(913, 10), 1246 => to_unsigned(741, 10), 1247 => to_unsigned(316, 10), 1248 => to_unsigned(470, 10), 1249 => to_unsigned(221, 10), 1250 => to_unsigned(500, 10), 1251 => to_unsigned(135, 10), 1252 => to_unsigned(664, 10), 1253 => to_unsigned(528, 10), 1254 => to_unsigned(707, 10), 1255 => to_unsigned(445, 10), 1256 => to_unsigned(237, 10), 1257 => to_unsigned(901, 10), 1258 => to_unsigned(497, 10), 1259 => to_unsigned(672, 10), 1260 => to_unsigned(688, 10), 1261 => to_unsigned(1006, 10), 1262 => to_unsigned(140, 10), 1263 => to_unsigned(769, 10), 1264 => to_unsigned(965, 10), 1265 => to_unsigned(171, 10), 1266 => to_unsigned(914, 10), 1267 => to_unsigned(841, 10), 1268 => to_unsigned(802, 10), 1269 => to_unsigned(696, 10), 1270 => to_unsigned(240, 10), 1271 => to_unsigned(746, 10), 1272 => to_unsigned(125, 10), 1273 => to_unsigned(616, 10), 1274 => to_unsigned(499, 10), 1275 => to_unsigned(213, 10), 1276 => to_unsigned(556, 10), 1277 => to_unsigned(889, 10), 1278 => to_unsigned(960, 10), 1279 => to_unsigned(761, 10), 1280 => to_unsigned(696, 10), 1281 => to_unsigned(970, 10), 1282 => to_unsigned(692, 10), 1283 => to_unsigned(121, 10), 1284 => to_unsigned(10, 10), 1285 => to_unsigned(92, 10), 1286 => to_unsigned(20, 10), 1287 => to_unsigned(918, 10), 1288 => to_unsigned(693, 10), 1289 => to_unsigned(98, 10), 1290 => to_unsigned(193, 10), 1291 => to_unsigned(902, 10), 1292 => to_unsigned(517, 10), 1293 => to_unsigned(352, 10), 1294 => to_unsigned(46, 10), 1295 => to_unsigned(713, 10), 1296 => to_unsigned(297, 10), 1297 => to_unsigned(216, 10), 1298 => to_unsigned(880, 10), 1299 => to_unsigned(115, 10), 1300 => to_unsigned(673, 10), 1301 => to_unsigned(804, 10), 1302 => to_unsigned(814, 10), 1303 => to_unsigned(363, 10), 1304 => to_unsigned(1012, 10), 1305 => to_unsigned(75, 10), 1306 => to_unsigned(364, 10), 1307 => to_unsigned(369, 10), 1308 => to_unsigned(448, 10), 1309 => to_unsigned(290, 10), 1310 => to_unsigned(188, 10), 1311 => to_unsigned(780, 10), 1312 => to_unsigned(697, 10), 1313 => to_unsigned(421, 10), 1314 => to_unsigned(448, 10), 1315 => to_unsigned(84, 10), 1316 => to_unsigned(555, 10), 1317 => to_unsigned(703, 10), 1318 => to_unsigned(197, 10), 1319 => to_unsigned(753, 10), 1320 => to_unsigned(977, 10), 1321 => to_unsigned(801, 10), 1322 => to_unsigned(161, 10), 1323 => to_unsigned(583, 10), 1324 => to_unsigned(243, 10), 1325 => to_unsigned(202, 10), 1326 => to_unsigned(583, 10), 1327 => to_unsigned(491, 10), 1328 => to_unsigned(642, 10), 1329 => to_unsigned(67, 10), 1330 => to_unsigned(780, 10), 1331 => to_unsigned(682, 10), 1332 => to_unsigned(526, 10), 1333 => to_unsigned(34, 10), 1334 => to_unsigned(355, 10), 1335 => to_unsigned(149, 10), 1336 => to_unsigned(919, 10), 1337 => to_unsigned(136, 10), 1338 => to_unsigned(1008, 10), 1339 => to_unsigned(665, 10), 1340 => to_unsigned(908, 10), 1341 => to_unsigned(809, 10), 1342 => to_unsigned(681, 10), 1343 => to_unsigned(998, 10), 1344 => to_unsigned(294, 10), 1345 => to_unsigned(638, 10), 1346 => to_unsigned(121, 10), 1347 => to_unsigned(687, 10), 1348 => to_unsigned(395, 10), 1349 => to_unsigned(518, 10), 1350 => to_unsigned(971, 10), 1351 => to_unsigned(911, 10), 1352 => to_unsigned(337, 10), 1353 => to_unsigned(1012, 10), 1354 => to_unsigned(146, 10), 1355 => to_unsigned(756, 10), 1356 => to_unsigned(517, 10), 1357 => to_unsigned(122, 10), 1358 => to_unsigned(399, 10), 1359 => to_unsigned(5, 10), 1360 => to_unsigned(843, 10), 1361 => to_unsigned(611, 10), 1362 => to_unsigned(963, 10), 1363 => to_unsigned(929, 10), 1364 => to_unsigned(41, 10), 1365 => to_unsigned(720, 10), 1366 => to_unsigned(655, 10), 1367 => to_unsigned(556, 10), 1368 => to_unsigned(254, 10), 1369 => to_unsigned(237, 10), 1370 => to_unsigned(792, 10), 1371 => to_unsigned(674, 10), 1372 => to_unsigned(446, 10), 1373 => to_unsigned(708, 10), 1374 => to_unsigned(392, 10), 1375 => to_unsigned(176, 10), 1376 => to_unsigned(179, 10), 1377 => to_unsigned(804, 10), 1378 => to_unsigned(602, 10), 1379 => to_unsigned(171, 10), 1380 => to_unsigned(321, 10), 1381 => to_unsigned(273, 10), 1382 => to_unsigned(696, 10), 1383 => to_unsigned(650, 10), 1384 => to_unsigned(263, 10), 1385 => to_unsigned(709, 10), 1386 => to_unsigned(922, 10), 1387 => to_unsigned(443, 10), 1388 => to_unsigned(10, 10), 1389 => to_unsigned(409, 10), 1390 => to_unsigned(166, 10), 1391 => to_unsigned(334, 10), 1392 => to_unsigned(942, 10), 1393 => to_unsigned(251, 10), 1394 => to_unsigned(985, 10), 1395 => to_unsigned(53, 10), 1396 => to_unsigned(236, 10), 1397 => to_unsigned(448, 10), 1398 => to_unsigned(630, 10), 1399 => to_unsigned(221, 10), 1400 => to_unsigned(507, 10), 1401 => to_unsigned(906, 10), 1402 => to_unsigned(725, 10), 1403 => to_unsigned(547, 10), 1404 => to_unsigned(437, 10), 1405 => to_unsigned(565, 10), 1406 => to_unsigned(956, 10), 1407 => to_unsigned(725, 10), 1408 => to_unsigned(988, 10), 1409 => to_unsigned(638, 10), 1410 => to_unsigned(25, 10), 1411 => to_unsigned(191, 10), 1412 => to_unsigned(644, 10), 1413 => to_unsigned(845, 10), 1414 => to_unsigned(719, 10), 1415 => to_unsigned(10, 10), 1416 => to_unsigned(279, 10), 1417 => to_unsigned(997, 10), 1418 => to_unsigned(872, 10), 1419 => to_unsigned(641, 10), 1420 => to_unsigned(954, 10), 1421 => to_unsigned(835, 10), 1422 => to_unsigned(540, 10), 1423 => to_unsigned(141, 10), 1424 => to_unsigned(717, 10), 1425 => to_unsigned(512, 10), 1426 => to_unsigned(318, 10), 1427 => to_unsigned(66, 10), 1428 => to_unsigned(183, 10), 1429 => to_unsigned(378, 10), 1430 => to_unsigned(318, 10), 1431 => to_unsigned(733, 10), 1432 => to_unsigned(872, 10), 1433 => to_unsigned(826, 10), 1434 => to_unsigned(716, 10), 1435 => to_unsigned(253, 10), 1436 => to_unsigned(478, 10), 1437 => to_unsigned(285, 10), 1438 => to_unsigned(664, 10), 1439 => to_unsigned(694, 10), 1440 => to_unsigned(253, 10), 1441 => to_unsigned(501, 10), 1442 => to_unsigned(246, 10), 1443 => to_unsigned(205, 10), 1444 => to_unsigned(1022, 10), 1445 => to_unsigned(778, 10), 1446 => to_unsigned(157, 10), 1447 => to_unsigned(450, 10), 1448 => to_unsigned(765, 10), 1449 => to_unsigned(199, 10), 1450 => to_unsigned(764, 10), 1451 => to_unsigned(67, 10), 1452 => to_unsigned(816, 10), 1453 => to_unsigned(860, 10), 1454 => to_unsigned(228, 10), 1455 => to_unsigned(623, 10), 1456 => to_unsigned(509, 10), 1457 => to_unsigned(160, 10), 1458 => to_unsigned(894, 10), 1459 => to_unsigned(618, 10), 1460 => to_unsigned(941, 10), 1461 => to_unsigned(951, 10), 1462 => to_unsigned(1005, 10), 1463 => to_unsigned(399, 10), 1464 => to_unsigned(630, 10), 1465 => to_unsigned(376, 10), 1466 => to_unsigned(448, 10), 1467 => to_unsigned(682, 10), 1468 => to_unsigned(159, 10), 1469 => to_unsigned(149, 10), 1470 => to_unsigned(137, 10), 1471 => to_unsigned(436, 10), 1472 => to_unsigned(432, 10), 1473 => to_unsigned(269, 10), 1474 => to_unsigned(375, 10), 1475 => to_unsigned(599, 10), 1476 => to_unsigned(308, 10), 1477 => to_unsigned(403, 10), 1478 => to_unsigned(985, 10), 1479 => to_unsigned(12, 10), 1480 => to_unsigned(869, 10), 1481 => to_unsigned(23, 10), 1482 => to_unsigned(757, 10), 1483 => to_unsigned(898, 10), 1484 => to_unsigned(70, 10), 1485 => to_unsigned(471, 10), 1486 => to_unsigned(92, 10), 1487 => to_unsigned(962, 10), 1488 => to_unsigned(759, 10), 1489 => to_unsigned(944, 10), 1490 => to_unsigned(596, 10), 1491 => to_unsigned(312, 10), 1492 => to_unsigned(225, 10), 1493 => to_unsigned(1008, 10), 1494 => to_unsigned(932, 10), 1495 => to_unsigned(290, 10), 1496 => to_unsigned(677, 10), 1497 => to_unsigned(107, 10), 1498 => to_unsigned(666, 10), 1499 => to_unsigned(930, 10), 1500 => to_unsigned(373, 10), 1501 => to_unsigned(869, 10), 1502 => to_unsigned(83, 10), 1503 => to_unsigned(119, 10), 1504 => to_unsigned(572, 10), 1505 => to_unsigned(926, 10), 1506 => to_unsigned(823, 10), 1507 => to_unsigned(401, 10), 1508 => to_unsigned(14, 10), 1509 => to_unsigned(396, 10), 1510 => to_unsigned(710, 10), 1511 => to_unsigned(549, 10), 1512 => to_unsigned(592, 10), 1513 => to_unsigned(664, 10), 1514 => to_unsigned(832, 10), 1515 => to_unsigned(990, 10), 1516 => to_unsigned(747, 10), 1517 => to_unsigned(719, 10), 1518 => to_unsigned(784, 10), 1519 => to_unsigned(91, 10), 1520 => to_unsigned(42, 10), 1521 => to_unsigned(260, 10), 1522 => to_unsigned(1020, 10), 1523 => to_unsigned(763, 10), 1524 => to_unsigned(37, 10), 1525 => to_unsigned(329, 10), 1526 => to_unsigned(70, 10), 1527 => to_unsigned(539, 10), 1528 => to_unsigned(800, 10), 1529 => to_unsigned(542, 10), 1530 => to_unsigned(630, 10), 1531 => to_unsigned(416, 10), 1532 => to_unsigned(420, 10), 1533 => to_unsigned(795, 10), 1534 => to_unsigned(614, 10), 1535 => to_unsigned(70, 10), 1536 => to_unsigned(583, 10), 1537 => to_unsigned(380, 10), 1538 => to_unsigned(545, 10), 1539 => to_unsigned(205, 10), 1540 => to_unsigned(692, 10), 1541 => to_unsigned(900, 10), 1542 => to_unsigned(70, 10), 1543 => to_unsigned(729, 10), 1544 => to_unsigned(617, 10), 1545 => to_unsigned(374, 10), 1546 => to_unsigned(984, 10), 1547 => to_unsigned(942, 10), 1548 => to_unsigned(319, 10), 1549 => to_unsigned(116, 10), 1550 => to_unsigned(178, 10), 1551 => to_unsigned(750, 10), 1552 => to_unsigned(657, 10), 1553 => to_unsigned(971, 10), 1554 => to_unsigned(125, 10), 1555 => to_unsigned(153, 10), 1556 => to_unsigned(626, 10), 1557 => to_unsigned(527, 10), 1558 => to_unsigned(595, 10), 1559 => to_unsigned(136, 10), 1560 => to_unsigned(143, 10), 1561 => to_unsigned(668, 10), 1562 => to_unsigned(283, 10), 1563 => to_unsigned(868, 10), 1564 => to_unsigned(765, 10), 1565 => to_unsigned(316, 10), 1566 => to_unsigned(756, 10), 1567 => to_unsigned(896, 10), 1568 => to_unsigned(404, 10), 1569 => to_unsigned(114, 10), 1570 => to_unsigned(707, 10), 1571 => to_unsigned(628, 10), 1572 => to_unsigned(532, 10), 1573 => to_unsigned(821, 10), 1574 => to_unsigned(600, 10), 1575 => to_unsigned(257, 10), 1576 => to_unsigned(830, 10), 1577 => to_unsigned(380, 10), 1578 => to_unsigned(482, 10), 1579 => to_unsigned(556, 10), 1580 => to_unsigned(95, 10), 1581 => to_unsigned(342, 10), 1582 => to_unsigned(547, 10), 1583 => to_unsigned(994, 10), 1584 => to_unsigned(446, 10), 1585 => to_unsigned(455, 10), 1586 => to_unsigned(402, 10), 1587 => to_unsigned(464, 10), 1588 => to_unsigned(543, 10), 1589 => to_unsigned(1020, 10), 1590 => to_unsigned(22, 10), 1591 => to_unsigned(973, 10), 1592 => to_unsigned(196, 10), 1593 => to_unsigned(583, 10), 1594 => to_unsigned(334, 10), 1595 => to_unsigned(258, 10), 1596 => to_unsigned(217, 10), 1597 => to_unsigned(602, 10), 1598 => to_unsigned(251, 10), 1599 => to_unsigned(173, 10), 1600 => to_unsigned(366, 10), 1601 => to_unsigned(839, 10), 1602 => to_unsigned(437, 10), 1603 => to_unsigned(654, 10), 1604 => to_unsigned(974, 10), 1605 => to_unsigned(436, 10), 1606 => to_unsigned(258, 10), 1607 => to_unsigned(972, 10), 1608 => to_unsigned(493, 10), 1609 => to_unsigned(129, 10), 1610 => to_unsigned(824, 10), 1611 => to_unsigned(98, 10), 1612 => to_unsigned(515, 10), 1613 => to_unsigned(333, 10), 1614 => to_unsigned(527, 10), 1615 => to_unsigned(515, 10), 1616 => to_unsigned(730, 10), 1617 => to_unsigned(158, 10), 1618 => to_unsigned(97, 10), 1619 => to_unsigned(939, 10), 1620 => to_unsigned(677, 10), 1621 => to_unsigned(899, 10), 1622 => to_unsigned(384, 10), 1623 => to_unsigned(509, 10), 1624 => to_unsigned(44, 10), 1625 => to_unsigned(159, 10), 1626 => to_unsigned(378, 10), 1627 => to_unsigned(216, 10), 1628 => to_unsigned(598, 10), 1629 => to_unsigned(288, 10), 1630 => to_unsigned(497, 10), 1631 => to_unsigned(834, 10), 1632 => to_unsigned(424, 10), 1633 => to_unsigned(457, 10), 1634 => to_unsigned(549, 10), 1635 => to_unsigned(738, 10), 1636 => to_unsigned(418, 10), 1637 => to_unsigned(1022, 10), 1638 => to_unsigned(588, 10), 1639 => to_unsigned(545, 10), 1640 => to_unsigned(79, 10), 1641 => to_unsigned(939, 10), 1642 => to_unsigned(856, 10), 1643 => to_unsigned(267, 10), 1644 => to_unsigned(615, 10), 1645 => to_unsigned(499, 10), 1646 => to_unsigned(972, 10), 1647 => to_unsigned(209, 10), 1648 => to_unsigned(699, 10), 1649 => to_unsigned(706, 10), 1650 => to_unsigned(1, 10), 1651 => to_unsigned(903, 10), 1652 => to_unsigned(922, 10), 1653 => to_unsigned(58, 10), 1654 => to_unsigned(791, 10), 1655 => to_unsigned(258, 10), 1656 => to_unsigned(37, 10), 1657 => to_unsigned(606, 10), 1658 => to_unsigned(479, 10), 1659 => to_unsigned(309, 10), 1660 => to_unsigned(653, 10), 1661 => to_unsigned(872, 10), 1662 => to_unsigned(460, 10), 1663 => to_unsigned(133, 10), 1664 => to_unsigned(55, 10), 1665 => to_unsigned(732, 10), 1666 => to_unsigned(11, 10), 1667 => to_unsigned(998, 10), 1668 => to_unsigned(656, 10), 1669 => to_unsigned(646, 10), 1670 => to_unsigned(963, 10), 1671 => to_unsigned(976, 10), 1672 => to_unsigned(766, 10), 1673 => to_unsigned(363, 10), 1674 => to_unsigned(622, 10), 1675 => to_unsigned(800, 10), 1676 => to_unsigned(471, 10), 1677 => to_unsigned(86, 10), 1678 => to_unsigned(193, 10), 1679 => to_unsigned(540, 10), 1680 => to_unsigned(259, 10), 1681 => to_unsigned(574, 10), 1682 => to_unsigned(496, 10), 1683 => to_unsigned(820, 10), 1684 => to_unsigned(368, 10), 1685 => to_unsigned(605, 10), 1686 => to_unsigned(947, 10), 1687 => to_unsigned(83, 10), 1688 => to_unsigned(21, 10), 1689 => to_unsigned(153, 10), 1690 => to_unsigned(815, 10), 1691 => to_unsigned(20, 10), 1692 => to_unsigned(533, 10), 1693 => to_unsigned(334, 10), 1694 => to_unsigned(754, 10), 1695 => to_unsigned(242, 10), 1696 => to_unsigned(815, 10), 1697 => to_unsigned(332, 10), 1698 => to_unsigned(129, 10), 1699 => to_unsigned(100, 10), 1700 => to_unsigned(950, 10), 1701 => to_unsigned(75, 10), 1702 => to_unsigned(283, 10), 1703 => to_unsigned(805, 10), 1704 => to_unsigned(869, 10), 1705 => to_unsigned(75, 10), 1706 => to_unsigned(956, 10), 1707 => to_unsigned(170, 10), 1708 => to_unsigned(511, 10), 1709 => to_unsigned(318, 10), 1710 => to_unsigned(46, 10), 1711 => to_unsigned(833, 10), 1712 => to_unsigned(484, 10), 1713 => to_unsigned(896, 10), 1714 => to_unsigned(835, 10), 1715 => to_unsigned(617, 10), 1716 => to_unsigned(222, 10), 1717 => to_unsigned(483, 10), 1718 => to_unsigned(55, 10), 1719 => to_unsigned(220, 10), 1720 => to_unsigned(842, 10), 1721 => to_unsigned(961, 10), 1722 => to_unsigned(1021, 10), 1723 => to_unsigned(674, 10), 1724 => to_unsigned(957, 10), 1725 => to_unsigned(22, 10), 1726 => to_unsigned(702, 10), 1727 => to_unsigned(131, 10), 1728 => to_unsigned(434, 10), 1729 => to_unsigned(415, 10), 1730 => to_unsigned(692, 10), 1731 => to_unsigned(269, 10), 1732 => to_unsigned(72, 10), 1733 => to_unsigned(79, 10), 1734 => to_unsigned(161, 10), 1735 => to_unsigned(286, 10), 1736 => to_unsigned(986, 10), 1737 => to_unsigned(372, 10), 1738 => to_unsigned(1015, 10), 1739 => to_unsigned(25, 10), 1740 => to_unsigned(839, 10), 1741 => to_unsigned(824, 10), 1742 => to_unsigned(888, 10), 1743 => to_unsigned(769, 10), 1744 => to_unsigned(660, 10), 1745 => to_unsigned(466, 10), 1746 => to_unsigned(900, 10), 1747 => to_unsigned(680, 10), 1748 => to_unsigned(133, 10), 1749 => to_unsigned(697, 10), 1750 => to_unsigned(593, 10), 1751 => to_unsigned(970, 10), 1752 => to_unsigned(544, 10), 1753 => to_unsigned(126, 10), 1754 => to_unsigned(586, 10), 1755 => to_unsigned(891, 10), 1756 => to_unsigned(511, 10), 1757 => to_unsigned(732, 10), 1758 => to_unsigned(835, 10), 1759 => to_unsigned(818, 10), 1760 => to_unsigned(634, 10), 1761 => to_unsigned(996, 10), 1762 => to_unsigned(443, 10), 1763 => to_unsigned(560, 10), 1764 => to_unsigned(826, 10), 1765 => to_unsigned(557, 10), 1766 => to_unsigned(177, 10), 1767 => to_unsigned(31, 10), 1768 => to_unsigned(41, 10), 1769 => to_unsigned(626, 10), 1770 => to_unsigned(231, 10), 1771 => to_unsigned(639, 10), 1772 => to_unsigned(206, 10), 1773 => to_unsigned(977, 10), 1774 => to_unsigned(591, 10), 1775 => to_unsigned(358, 10), 1776 => to_unsigned(573, 10), 1777 => to_unsigned(13, 10), 1778 => to_unsigned(592, 10), 1779 => to_unsigned(300, 10), 1780 => to_unsigned(747, 10), 1781 => to_unsigned(453, 10), 1782 => to_unsigned(991, 10), 1783 => to_unsigned(568, 10), 1784 => to_unsigned(977, 10), 1785 => to_unsigned(547, 10), 1786 => to_unsigned(477, 10), 1787 => to_unsigned(725, 10), 1788 => to_unsigned(803, 10), 1789 => to_unsigned(371, 10), 1790 => to_unsigned(826, 10), 1791 => to_unsigned(323, 10), 1792 => to_unsigned(791, 10), 1793 => to_unsigned(450, 10), 1794 => to_unsigned(92, 10), 1795 => to_unsigned(712, 10), 1796 => to_unsigned(518, 10), 1797 => to_unsigned(260, 10), 1798 => to_unsigned(1018, 10), 1799 => to_unsigned(230, 10), 1800 => to_unsigned(811, 10), 1801 => to_unsigned(698, 10), 1802 => to_unsigned(702, 10), 1803 => to_unsigned(924, 10), 1804 => to_unsigned(854, 10), 1805 => to_unsigned(1002, 10), 1806 => to_unsigned(256, 10), 1807 => to_unsigned(905, 10), 1808 => to_unsigned(324, 10), 1809 => to_unsigned(510, 10), 1810 => to_unsigned(884, 10), 1811 => to_unsigned(1020, 10), 1812 => to_unsigned(305, 10), 1813 => to_unsigned(289, 10), 1814 => to_unsigned(290, 10), 1815 => to_unsigned(349, 10), 1816 => to_unsigned(478, 10), 1817 => to_unsigned(649, 10), 1818 => to_unsigned(767, 10), 1819 => to_unsigned(316, 10), 1820 => to_unsigned(934, 10), 1821 => to_unsigned(669, 10), 1822 => to_unsigned(672, 10), 1823 => to_unsigned(487, 10), 1824 => to_unsigned(179, 10), 1825 => to_unsigned(445, 10), 1826 => to_unsigned(742, 10), 1827 => to_unsigned(65, 10), 1828 => to_unsigned(592, 10), 1829 => to_unsigned(851, 10), 1830 => to_unsigned(743, 10), 1831 => to_unsigned(29, 10), 1832 => to_unsigned(734, 10), 1833 => to_unsigned(601, 10), 1834 => to_unsigned(626, 10), 1835 => to_unsigned(832, 10), 1836 => to_unsigned(144, 10), 1837 => to_unsigned(608, 10), 1838 => to_unsigned(307, 10), 1839 => to_unsigned(642, 10), 1840 => to_unsigned(469, 10), 1841 => to_unsigned(1018, 10), 1842 => to_unsigned(605, 10), 1843 => to_unsigned(252, 10), 1844 => to_unsigned(985, 10), 1845 => to_unsigned(676, 10), 1846 => to_unsigned(189, 10), 1847 => to_unsigned(581, 10), 1848 => to_unsigned(74, 10), 1849 => to_unsigned(539, 10), 1850 => to_unsigned(748, 10), 1851 => to_unsigned(951, 10), 1852 => to_unsigned(276, 10), 1853 => to_unsigned(808, 10), 1854 => to_unsigned(433, 10), 1855 => to_unsigned(641, 10), 1856 => to_unsigned(84, 10), 1857 => to_unsigned(15, 10), 1858 => to_unsigned(358, 10), 1859 => to_unsigned(509, 10), 1860 => to_unsigned(138, 10), 1861 => to_unsigned(628, 10), 1862 => to_unsigned(862, 10), 1863 => to_unsigned(16, 10), 1864 => to_unsigned(960, 10), 1865 => to_unsigned(137, 10), 1866 => to_unsigned(411, 10), 1867 => to_unsigned(615, 10), 1868 => to_unsigned(275, 10), 1869 => to_unsigned(203, 10), 1870 => to_unsigned(405, 10), 1871 => to_unsigned(521, 10), 1872 => to_unsigned(369, 10), 1873 => to_unsigned(12, 10), 1874 => to_unsigned(1017, 10), 1875 => to_unsigned(138, 10), 1876 => to_unsigned(763, 10), 1877 => to_unsigned(205, 10), 1878 => to_unsigned(61, 10), 1879 => to_unsigned(555, 10), 1880 => to_unsigned(201, 10), 1881 => to_unsigned(520, 10), 1882 => to_unsigned(713, 10), 1883 => to_unsigned(242, 10), 1884 => to_unsigned(341, 10), 1885 => to_unsigned(9, 10), 1886 => to_unsigned(742, 10), 1887 => to_unsigned(415, 10), 1888 => to_unsigned(4, 10), 1889 => to_unsigned(886, 10), 1890 => to_unsigned(378, 10), 1891 => to_unsigned(960, 10), 1892 => to_unsigned(784, 10), 1893 => to_unsigned(800, 10), 1894 => to_unsigned(381, 10), 1895 => to_unsigned(447, 10), 1896 => to_unsigned(925, 10), 1897 => to_unsigned(804, 10), 1898 => to_unsigned(942, 10), 1899 => to_unsigned(649, 10), 1900 => to_unsigned(609, 10), 1901 => to_unsigned(735, 10), 1902 => to_unsigned(971, 10), 1903 => to_unsigned(429, 10), 1904 => to_unsigned(672, 10), 1905 => to_unsigned(594, 10), 1906 => to_unsigned(984, 10), 1907 => to_unsigned(152, 10), 1908 => to_unsigned(944, 10), 1909 => to_unsigned(827, 10), 1910 => to_unsigned(933, 10), 1911 => to_unsigned(851, 10), 1912 => to_unsigned(38, 10), 1913 => to_unsigned(656, 10), 1914 => to_unsigned(189, 10), 1915 => to_unsigned(274, 10), 1916 => to_unsigned(227, 10), 1917 => to_unsigned(624, 10), 1918 => to_unsigned(335, 10), 1919 => to_unsigned(202, 10), 1920 => to_unsigned(993, 10), 1921 => to_unsigned(91, 10), 1922 => to_unsigned(735, 10), 1923 => to_unsigned(347, 10), 1924 => to_unsigned(665, 10), 1925 => to_unsigned(137, 10), 1926 => to_unsigned(341, 10), 1927 => to_unsigned(949, 10), 1928 => to_unsigned(209, 10), 1929 => to_unsigned(645, 10), 1930 => to_unsigned(229, 10), 1931 => to_unsigned(825, 10), 1932 => to_unsigned(69, 10), 1933 => to_unsigned(197, 10), 1934 => to_unsigned(738, 10), 1935 => to_unsigned(944, 10), 1936 => to_unsigned(780, 10), 1937 => to_unsigned(977, 10), 1938 => to_unsigned(492, 10), 1939 => to_unsigned(598, 10), 1940 => to_unsigned(58, 10), 1941 => to_unsigned(149, 10), 1942 => to_unsigned(113, 10), 1943 => to_unsigned(866, 10), 1944 => to_unsigned(120, 10), 1945 => to_unsigned(546, 10), 1946 => to_unsigned(740, 10), 1947 => to_unsigned(369, 10), 1948 => to_unsigned(444, 10), 1949 => to_unsigned(809, 10), 1950 => to_unsigned(652, 10), 1951 => to_unsigned(155, 10), 1952 => to_unsigned(699, 10), 1953 => to_unsigned(27, 10), 1954 => to_unsigned(901, 10), 1955 => to_unsigned(396, 10), 1956 => to_unsigned(580, 10), 1957 => to_unsigned(759, 10), 1958 => to_unsigned(63, 10), 1959 => to_unsigned(500, 10), 1960 => to_unsigned(980, 10), 1961 => to_unsigned(703, 10), 1962 => to_unsigned(386, 10), 1963 => to_unsigned(536, 10), 1964 => to_unsigned(527, 10), 1965 => to_unsigned(209, 10), 1966 => to_unsigned(350, 10), 1967 => to_unsigned(525, 10), 1968 => to_unsigned(939, 10), 1969 => to_unsigned(345, 10), 1970 => to_unsigned(443, 10), 1971 => to_unsigned(860, 10), 1972 => to_unsigned(309, 10), 1973 => to_unsigned(399, 10), 1974 => to_unsigned(260, 10), 1975 => to_unsigned(64, 10), 1976 => to_unsigned(98, 10), 1977 => to_unsigned(505, 10), 1978 => to_unsigned(720, 10), 1979 => to_unsigned(162, 10), 1980 => to_unsigned(137, 10), 1981 => to_unsigned(709, 10), 1982 => to_unsigned(329, 10), 1983 => to_unsigned(262, 10), 1984 => to_unsigned(194, 10), 1985 => to_unsigned(896, 10), 1986 => to_unsigned(310, 10), 1987 => to_unsigned(801, 10), 1988 => to_unsigned(480, 10), 1989 => to_unsigned(89, 10), 1990 => to_unsigned(321, 10), 1991 => to_unsigned(692, 10), 1992 => to_unsigned(743, 10), 1993 => to_unsigned(550, 10), 1994 => to_unsigned(857, 10), 1995 => to_unsigned(768, 10), 1996 => to_unsigned(439, 10), 1997 => to_unsigned(377, 10), 1998 => to_unsigned(792, 10), 1999 => to_unsigned(732, 10), 2000 => to_unsigned(703, 10), 2001 => to_unsigned(254, 10), 2002 => to_unsigned(8, 10), 2003 => to_unsigned(283, 10), 2004 => to_unsigned(263, 10), 2005 => to_unsigned(188, 10), 2006 => to_unsigned(935, 10), 2007 => to_unsigned(643, 10), 2008 => to_unsigned(626, 10), 2009 => to_unsigned(356, 10), 2010 => to_unsigned(777, 10), 2011 => to_unsigned(318, 10), 2012 => to_unsigned(24, 10), 2013 => to_unsigned(959, 10), 2014 => to_unsigned(249, 10), 2015 => to_unsigned(749, 10), 2016 => to_unsigned(236, 10), 2017 => to_unsigned(998, 10), 2018 => to_unsigned(214, 10), 2019 => to_unsigned(707, 10), 2020 => to_unsigned(625, 10), 2021 => to_unsigned(1011, 10), 2022 => to_unsigned(584, 10), 2023 => to_unsigned(745, 10), 2024 => to_unsigned(689, 10), 2025 => to_unsigned(244, 10), 2026 => to_unsigned(148, 10), 2027 => to_unsigned(668, 10), 2028 => to_unsigned(716, 10), 2029 => to_unsigned(307, 10), 2030 => to_unsigned(174, 10), 2031 => to_unsigned(207, 10), 2032 => to_unsigned(729, 10), 2033 => to_unsigned(772, 10), 2034 => to_unsigned(556, 10), 2035 => to_unsigned(23, 10), 2036 => to_unsigned(948, 10), 2037 => to_unsigned(191, 10), 2038 => to_unsigned(27, 10), 2039 => to_unsigned(242, 10), 2040 => to_unsigned(696, 10), 2041 => to_unsigned(144, 10), 2042 => to_unsigned(127, 10), 2043 => to_unsigned(485, 10), 2044 => to_unsigned(979, 10), 2045 => to_unsigned(574, 10), 2046 => to_unsigned(309, 10), 2047 => to_unsigned(17, 10)),
            9 => (0 => to_unsigned(484, 10), 1 => to_unsigned(604, 10), 2 => to_unsigned(622, 10), 3 => to_unsigned(165, 10), 4 => to_unsigned(915, 10), 5 => to_unsigned(334, 10), 6 => to_unsigned(868, 10), 7 => to_unsigned(757, 10), 8 => to_unsigned(116, 10), 9 => to_unsigned(25, 10), 10 => to_unsigned(472, 10), 11 => to_unsigned(451, 10), 12 => to_unsigned(636, 10), 13 => to_unsigned(788, 10), 14 => to_unsigned(816, 10), 15 => to_unsigned(489, 10), 16 => to_unsigned(683, 10), 17 => to_unsigned(658, 10), 18 => to_unsigned(44, 10), 19 => to_unsigned(813, 10), 20 => to_unsigned(92, 10), 21 => to_unsigned(72, 10), 22 => to_unsigned(565, 10), 23 => to_unsigned(295, 10), 24 => to_unsigned(206, 10), 25 => to_unsigned(545, 10), 26 => to_unsigned(472, 10), 27 => to_unsigned(89, 10), 28 => to_unsigned(914, 10), 29 => to_unsigned(878, 10), 30 => to_unsigned(195, 10), 31 => to_unsigned(535, 10), 32 => to_unsigned(50, 10), 33 => to_unsigned(508, 10), 34 => to_unsigned(354, 10), 35 => to_unsigned(660, 10), 36 => to_unsigned(815, 10), 37 => to_unsigned(232, 10), 38 => to_unsigned(350, 10), 39 => to_unsigned(89, 10), 40 => to_unsigned(484, 10), 41 => to_unsigned(682, 10), 42 => to_unsigned(785, 10), 43 => to_unsigned(85, 10), 44 => to_unsigned(316, 10), 45 => to_unsigned(196, 10), 46 => to_unsigned(691, 10), 47 => to_unsigned(609, 10), 48 => to_unsigned(199, 10), 49 => to_unsigned(35, 10), 50 => to_unsigned(264, 10), 51 => to_unsigned(301, 10), 52 => to_unsigned(581, 10), 53 => to_unsigned(71, 10), 54 => to_unsigned(674, 10), 55 => to_unsigned(504, 10), 56 => to_unsigned(24, 10), 57 => to_unsigned(321, 10), 58 => to_unsigned(97, 10), 59 => to_unsigned(923, 10), 60 => to_unsigned(133, 10), 61 => to_unsigned(17, 10), 62 => to_unsigned(56, 10), 63 => to_unsigned(99, 10), 64 => to_unsigned(283, 10), 65 => to_unsigned(607, 10), 66 => to_unsigned(974, 10), 67 => to_unsigned(716, 10), 68 => to_unsigned(556, 10), 69 => to_unsigned(171, 10), 70 => to_unsigned(186, 10), 71 => to_unsigned(793, 10), 72 => to_unsigned(99, 10), 73 => to_unsigned(264, 10), 74 => to_unsigned(818, 10), 75 => to_unsigned(185, 10), 76 => to_unsigned(683, 10), 77 => to_unsigned(589, 10), 78 => to_unsigned(275, 10), 79 => to_unsigned(56, 10), 80 => to_unsigned(48, 10), 81 => to_unsigned(493, 10), 82 => to_unsigned(716, 10), 83 => to_unsigned(443, 10), 84 => to_unsigned(846, 10), 85 => to_unsigned(898, 10), 86 => to_unsigned(888, 10), 87 => to_unsigned(810, 10), 88 => to_unsigned(423, 10), 89 => to_unsigned(756, 10), 90 => to_unsigned(673, 10), 91 => to_unsigned(624, 10), 92 => to_unsigned(690, 10), 93 => to_unsigned(950, 10), 94 => to_unsigned(274, 10), 95 => to_unsigned(243, 10), 96 => to_unsigned(798, 10), 97 => to_unsigned(903, 10), 98 => to_unsigned(972, 10), 99 => to_unsigned(371, 10), 100 => to_unsigned(589, 10), 101 => to_unsigned(718, 10), 102 => to_unsigned(468, 10), 103 => to_unsigned(315, 10), 104 => to_unsigned(467, 10), 105 => to_unsigned(110, 10), 106 => to_unsigned(552, 10), 107 => to_unsigned(745, 10), 108 => to_unsigned(845, 10), 109 => to_unsigned(968, 10), 110 => to_unsigned(402, 10), 111 => to_unsigned(961, 10), 112 => to_unsigned(398, 10), 113 => to_unsigned(745, 10), 114 => to_unsigned(516, 10), 115 => to_unsigned(522, 10), 116 => to_unsigned(354, 10), 117 => to_unsigned(383, 10), 118 => to_unsigned(696, 10), 119 => to_unsigned(486, 10), 120 => to_unsigned(374, 10), 121 => to_unsigned(678, 10), 122 => to_unsigned(951, 10), 123 => to_unsigned(34, 10), 124 => to_unsigned(375, 10), 125 => to_unsigned(853, 10), 126 => to_unsigned(649, 10), 127 => to_unsigned(421, 10), 128 => to_unsigned(316, 10), 129 => to_unsigned(578, 10), 130 => to_unsigned(532, 10), 131 => to_unsigned(82, 10), 132 => to_unsigned(453, 10), 133 => to_unsigned(591, 10), 134 => to_unsigned(922, 10), 135 => to_unsigned(1006, 10), 136 => to_unsigned(210, 10), 137 => to_unsigned(48, 10), 138 => to_unsigned(1023, 10), 139 => to_unsigned(884, 10), 140 => to_unsigned(815, 10), 141 => to_unsigned(130, 10), 142 => to_unsigned(545, 10), 143 => to_unsigned(957, 10), 144 => to_unsigned(589, 10), 145 => to_unsigned(150, 10), 146 => to_unsigned(847, 10), 147 => to_unsigned(989, 10), 148 => to_unsigned(262, 10), 149 => to_unsigned(786, 10), 150 => to_unsigned(670, 10), 151 => to_unsigned(983, 10), 152 => to_unsigned(614, 10), 153 => to_unsigned(476, 10), 154 => to_unsigned(633, 10), 155 => to_unsigned(73, 10), 156 => to_unsigned(395, 10), 157 => to_unsigned(410, 10), 158 => to_unsigned(820, 10), 159 => to_unsigned(988, 10), 160 => to_unsigned(313, 10), 161 => to_unsigned(746, 10), 162 => to_unsigned(163, 10), 163 => to_unsigned(265, 10), 164 => to_unsigned(61, 10), 165 => to_unsigned(758, 10), 166 => to_unsigned(907, 10), 167 => to_unsigned(274, 10), 168 => to_unsigned(540, 10), 169 => to_unsigned(229, 10), 170 => to_unsigned(747, 10), 171 => to_unsigned(299, 10), 172 => to_unsigned(267, 10), 173 => to_unsigned(105, 10), 174 => to_unsigned(148, 10), 175 => to_unsigned(249, 10), 176 => to_unsigned(170, 10), 177 => to_unsigned(369, 10), 178 => to_unsigned(257, 10), 179 => to_unsigned(530, 10), 180 => to_unsigned(783, 10), 181 => to_unsigned(810, 10), 182 => to_unsigned(799, 10), 183 => to_unsigned(569, 10), 184 => to_unsigned(109, 10), 185 => to_unsigned(598, 10), 186 => to_unsigned(809, 10), 187 => to_unsigned(60, 10), 188 => to_unsigned(110, 10), 189 => to_unsigned(28, 10), 190 => to_unsigned(220, 10), 191 => to_unsigned(367, 10), 192 => to_unsigned(935, 10), 193 => to_unsigned(248, 10), 194 => to_unsigned(426, 10), 195 => to_unsigned(498, 10), 196 => to_unsigned(249, 10), 197 => to_unsigned(73, 10), 198 => to_unsigned(151, 10), 199 => to_unsigned(710, 10), 200 => to_unsigned(103, 10), 201 => to_unsigned(74, 10), 202 => to_unsigned(585, 10), 203 => to_unsigned(514, 10), 204 => to_unsigned(434, 10), 205 => to_unsigned(353, 10), 206 => to_unsigned(590, 10), 207 => to_unsigned(349, 10), 208 => to_unsigned(330, 10), 209 => to_unsigned(56, 10), 210 => to_unsigned(448, 10), 211 => to_unsigned(424, 10), 212 => to_unsigned(96, 10), 213 => to_unsigned(470, 10), 214 => to_unsigned(906, 10), 215 => to_unsigned(199, 10), 216 => to_unsigned(187, 10), 217 => to_unsigned(85, 10), 218 => to_unsigned(232, 10), 219 => to_unsigned(303, 10), 220 => to_unsigned(445, 10), 221 => to_unsigned(106, 10), 222 => to_unsigned(812, 10), 223 => to_unsigned(20, 10), 224 => to_unsigned(433, 10), 225 => to_unsigned(678, 10), 226 => to_unsigned(144, 10), 227 => to_unsigned(337, 10), 228 => to_unsigned(471, 10), 229 => to_unsigned(760, 10), 230 => to_unsigned(295, 10), 231 => to_unsigned(949, 10), 232 => to_unsigned(224, 10), 233 => to_unsigned(366, 10), 234 => to_unsigned(487, 10), 235 => to_unsigned(1022, 10), 236 => to_unsigned(241, 10), 237 => to_unsigned(320, 10), 238 => to_unsigned(462, 10), 239 => to_unsigned(451, 10), 240 => to_unsigned(325, 10), 241 => to_unsigned(630, 10), 242 => to_unsigned(549, 10), 243 => to_unsigned(11, 10), 244 => to_unsigned(65, 10), 245 => to_unsigned(3, 10), 246 => to_unsigned(251, 10), 247 => to_unsigned(70, 10), 248 => to_unsigned(290, 10), 249 => to_unsigned(699, 10), 250 => to_unsigned(489, 10), 251 => to_unsigned(347, 10), 252 => to_unsigned(786, 10), 253 => to_unsigned(9, 10), 254 => to_unsigned(873, 10), 255 => to_unsigned(1019, 10), 256 => to_unsigned(100, 10), 257 => to_unsigned(269, 10), 258 => to_unsigned(114, 10), 259 => to_unsigned(216, 10), 260 => to_unsigned(231, 10), 261 => to_unsigned(1006, 10), 262 => to_unsigned(583, 10), 263 => to_unsigned(89, 10), 264 => to_unsigned(845, 10), 265 => to_unsigned(798, 10), 266 => to_unsigned(838, 10), 267 => to_unsigned(946, 10), 268 => to_unsigned(136, 10), 269 => to_unsigned(233, 10), 270 => to_unsigned(819, 10), 271 => to_unsigned(794, 10), 272 => to_unsigned(650, 10), 273 => to_unsigned(290, 10), 274 => to_unsigned(821, 10), 275 => to_unsigned(537, 10), 276 => to_unsigned(68, 10), 277 => to_unsigned(879, 10), 278 => to_unsigned(394, 10), 279 => to_unsigned(589, 10), 280 => to_unsigned(94, 10), 281 => to_unsigned(830, 10), 282 => to_unsigned(767, 10), 283 => to_unsigned(95, 10), 284 => to_unsigned(162, 10), 285 => to_unsigned(102, 10), 286 => to_unsigned(471, 10), 287 => to_unsigned(817, 10), 288 => to_unsigned(318, 10), 289 => to_unsigned(492, 10), 290 => to_unsigned(226, 10), 291 => to_unsigned(888, 10), 292 => to_unsigned(336, 10), 293 => to_unsigned(534, 10), 294 => to_unsigned(153, 10), 295 => to_unsigned(203, 10), 296 => to_unsigned(519, 10), 297 => to_unsigned(1017, 10), 298 => to_unsigned(638, 10), 299 => to_unsigned(180, 10), 300 => to_unsigned(708, 10), 301 => to_unsigned(156, 10), 302 => to_unsigned(729, 10), 303 => to_unsigned(612, 10), 304 => to_unsigned(361, 10), 305 => to_unsigned(970, 10), 306 => to_unsigned(503, 10), 307 => to_unsigned(403, 10), 308 => to_unsigned(250, 10), 309 => to_unsigned(789, 10), 310 => to_unsigned(1014, 10), 311 => to_unsigned(407, 10), 312 => to_unsigned(31, 10), 313 => to_unsigned(93, 10), 314 => to_unsigned(237, 10), 315 => to_unsigned(181, 10), 316 => to_unsigned(864, 10), 317 => to_unsigned(555, 10), 318 => to_unsigned(20, 10), 319 => to_unsigned(382, 10), 320 => to_unsigned(848, 10), 321 => to_unsigned(1, 10), 322 => to_unsigned(260, 10), 323 => to_unsigned(629, 10), 324 => to_unsigned(158, 10), 325 => to_unsigned(605, 10), 326 => to_unsigned(494, 10), 327 => to_unsigned(40, 10), 328 => to_unsigned(905, 10), 329 => to_unsigned(61, 10), 330 => to_unsigned(865, 10), 331 => to_unsigned(1, 10), 332 => to_unsigned(281, 10), 333 => to_unsigned(976, 10), 334 => to_unsigned(26, 10), 335 => to_unsigned(609, 10), 336 => to_unsigned(329, 10), 337 => to_unsigned(39, 10), 338 => to_unsigned(923, 10), 339 => to_unsigned(316, 10), 340 => to_unsigned(966, 10), 341 => to_unsigned(488, 10), 342 => to_unsigned(858, 10), 343 => to_unsigned(924, 10), 344 => to_unsigned(833, 10), 345 => to_unsigned(725, 10), 346 => to_unsigned(336, 10), 347 => to_unsigned(337, 10), 348 => to_unsigned(198, 10), 349 => to_unsigned(41, 10), 350 => to_unsigned(61, 10), 351 => to_unsigned(941, 10), 352 => to_unsigned(81, 10), 353 => to_unsigned(489, 10), 354 => to_unsigned(133, 10), 355 => to_unsigned(225, 10), 356 => to_unsigned(836, 10), 357 => to_unsigned(492, 10), 358 => to_unsigned(105, 10), 359 => to_unsigned(543, 10), 360 => to_unsigned(681, 10), 361 => to_unsigned(183, 10), 362 => to_unsigned(229, 10), 363 => to_unsigned(942, 10), 364 => to_unsigned(366, 10), 365 => to_unsigned(403, 10), 366 => to_unsigned(932, 10), 367 => to_unsigned(487, 10), 368 => to_unsigned(774, 10), 369 => to_unsigned(894, 10), 370 => to_unsigned(116, 10), 371 => to_unsigned(553, 10), 372 => to_unsigned(77, 10), 373 => to_unsigned(961, 10), 374 => to_unsigned(454, 10), 375 => to_unsigned(666, 10), 376 => to_unsigned(680, 10), 377 => to_unsigned(642, 10), 378 => to_unsigned(332, 10), 379 => to_unsigned(343, 10), 380 => to_unsigned(686, 10), 381 => to_unsigned(84, 10), 382 => to_unsigned(562, 10), 383 => to_unsigned(489, 10), 384 => to_unsigned(241, 10), 385 => to_unsigned(195, 10), 386 => to_unsigned(259, 10), 387 => to_unsigned(101, 10), 388 => to_unsigned(274, 10), 389 => to_unsigned(63, 10), 390 => to_unsigned(644, 10), 391 => to_unsigned(752, 10), 392 => to_unsigned(236, 10), 393 => to_unsigned(135, 10), 394 => to_unsigned(401, 10), 395 => to_unsigned(305, 10), 396 => to_unsigned(667, 10), 397 => to_unsigned(49, 10), 398 => to_unsigned(96, 10), 399 => to_unsigned(474, 10), 400 => to_unsigned(206, 10), 401 => to_unsigned(497, 10), 402 => to_unsigned(589, 10), 403 => to_unsigned(778, 10), 404 => to_unsigned(167, 10), 405 => to_unsigned(985, 10), 406 => to_unsigned(863, 10), 407 => to_unsigned(299, 10), 408 => to_unsigned(789, 10), 409 => to_unsigned(297, 10), 410 => to_unsigned(125, 10), 411 => to_unsigned(650, 10), 412 => to_unsigned(682, 10), 413 => to_unsigned(489, 10), 414 => to_unsigned(579, 10), 415 => to_unsigned(966, 10), 416 => to_unsigned(938, 10), 417 => to_unsigned(464, 10), 418 => to_unsigned(31, 10), 419 => to_unsigned(190, 10), 420 => to_unsigned(65, 10), 421 => to_unsigned(214, 10), 422 => to_unsigned(938, 10), 423 => to_unsigned(225, 10), 424 => to_unsigned(135, 10), 425 => to_unsigned(312, 10), 426 => to_unsigned(2, 10), 427 => to_unsigned(159, 10), 428 => to_unsigned(665, 10), 429 => to_unsigned(691, 10), 430 => to_unsigned(73, 10), 431 => to_unsigned(299, 10), 432 => to_unsigned(225, 10), 433 => to_unsigned(549, 10), 434 => to_unsigned(869, 10), 435 => to_unsigned(130, 10), 436 => to_unsigned(696, 10), 437 => to_unsigned(357, 10), 438 => to_unsigned(363, 10), 439 => to_unsigned(51, 10), 440 => to_unsigned(499, 10), 441 => to_unsigned(67, 10), 442 => to_unsigned(484, 10), 443 => to_unsigned(983, 10), 444 => to_unsigned(38, 10), 445 => to_unsigned(712, 10), 446 => to_unsigned(435, 10), 447 => to_unsigned(515, 10), 448 => to_unsigned(356, 10), 449 => to_unsigned(795, 10), 450 => to_unsigned(461, 10), 451 => to_unsigned(462, 10), 452 => to_unsigned(285, 10), 453 => to_unsigned(115, 10), 454 => to_unsigned(823, 10), 455 => to_unsigned(668, 10), 456 => to_unsigned(112, 10), 457 => to_unsigned(318, 10), 458 => to_unsigned(362, 10), 459 => to_unsigned(578, 10), 460 => to_unsigned(412, 10), 461 => to_unsigned(465, 10), 462 => to_unsigned(294, 10), 463 => to_unsigned(513, 10), 464 => to_unsigned(603, 10), 465 => to_unsigned(358, 10), 466 => to_unsigned(287, 10), 467 => to_unsigned(910, 10), 468 => to_unsigned(167, 10), 469 => to_unsigned(702, 10), 470 => to_unsigned(359, 10), 471 => to_unsigned(378, 10), 472 => to_unsigned(956, 10), 473 => to_unsigned(885, 10), 474 => to_unsigned(634, 10), 475 => to_unsigned(611, 10), 476 => to_unsigned(988, 10), 477 => to_unsigned(456, 10), 478 => to_unsigned(902, 10), 479 => to_unsigned(197, 10), 480 => to_unsigned(1001, 10), 481 => to_unsigned(439, 10), 482 => to_unsigned(556, 10), 483 => to_unsigned(921, 10), 484 => to_unsigned(514, 10), 485 => to_unsigned(730, 10), 486 => to_unsigned(492, 10), 487 => to_unsigned(378, 10), 488 => to_unsigned(655, 10), 489 => to_unsigned(69, 10), 490 => to_unsigned(342, 10), 491 => to_unsigned(778, 10), 492 => to_unsigned(128, 10), 493 => to_unsigned(311, 10), 494 => to_unsigned(149, 10), 495 => to_unsigned(392, 10), 496 => to_unsigned(864, 10), 497 => to_unsigned(529, 10), 498 => to_unsigned(780, 10), 499 => to_unsigned(415, 10), 500 => to_unsigned(381, 10), 501 => to_unsigned(502, 10), 502 => to_unsigned(51, 10), 503 => to_unsigned(230, 10), 504 => to_unsigned(961, 10), 505 => to_unsigned(356, 10), 506 => to_unsigned(436, 10), 507 => to_unsigned(811, 10), 508 => to_unsigned(979, 10), 509 => to_unsigned(265, 10), 510 => to_unsigned(814, 10), 511 => to_unsigned(722, 10), 512 => to_unsigned(247, 10), 513 => to_unsigned(313, 10), 514 => to_unsigned(198, 10), 515 => to_unsigned(995, 10), 516 => to_unsigned(102, 10), 517 => to_unsigned(741, 10), 518 => to_unsigned(614, 10), 519 => to_unsigned(77, 10), 520 => to_unsigned(515, 10), 521 => to_unsigned(547, 10), 522 => to_unsigned(449, 10), 523 => to_unsigned(778, 10), 524 => to_unsigned(406, 10), 525 => to_unsigned(497, 10), 526 => to_unsigned(248, 10), 527 => to_unsigned(398, 10), 528 => to_unsigned(533, 10), 529 => to_unsigned(449, 10), 530 => to_unsigned(868, 10), 531 => to_unsigned(688, 10), 532 => to_unsigned(132, 10), 533 => to_unsigned(110, 10), 534 => to_unsigned(461, 10), 535 => to_unsigned(514, 10), 536 => to_unsigned(614, 10), 537 => to_unsigned(226, 10), 538 => to_unsigned(535, 10), 539 => to_unsigned(494, 10), 540 => to_unsigned(160, 10), 541 => to_unsigned(204, 10), 542 => to_unsigned(237, 10), 543 => to_unsigned(578, 10), 544 => to_unsigned(106, 10), 545 => to_unsigned(371, 10), 546 => to_unsigned(200, 10), 547 => to_unsigned(354, 10), 548 => to_unsigned(257, 10), 549 => to_unsigned(19, 10), 550 => to_unsigned(472, 10), 551 => to_unsigned(858, 10), 552 => to_unsigned(50, 10), 553 => to_unsigned(688, 10), 554 => to_unsigned(932, 10), 555 => to_unsigned(721, 10), 556 => to_unsigned(863, 10), 557 => to_unsigned(405, 10), 558 => to_unsigned(674, 10), 559 => to_unsigned(209, 10), 560 => to_unsigned(932, 10), 561 => to_unsigned(826, 10), 562 => to_unsigned(865, 10), 563 => to_unsigned(650, 10), 564 => to_unsigned(260, 10), 565 => to_unsigned(410, 10), 566 => to_unsigned(348, 10), 567 => to_unsigned(752, 10), 568 => to_unsigned(114, 10), 569 => to_unsigned(608, 10), 570 => to_unsigned(219, 10), 571 => to_unsigned(668, 10), 572 => to_unsigned(97, 10), 573 => to_unsigned(267, 10), 574 => to_unsigned(759, 10), 575 => to_unsigned(79, 10), 576 => to_unsigned(628, 10), 577 => to_unsigned(444, 10), 578 => to_unsigned(110, 10), 579 => to_unsigned(935, 10), 580 => to_unsigned(99, 10), 581 => to_unsigned(295, 10), 582 => to_unsigned(372, 10), 583 => to_unsigned(688, 10), 584 => to_unsigned(184, 10), 585 => to_unsigned(280, 10), 586 => to_unsigned(433, 10), 587 => to_unsigned(67, 10), 588 => to_unsigned(52, 10), 589 => to_unsigned(109, 10), 590 => to_unsigned(834, 10), 591 => to_unsigned(862, 10), 592 => to_unsigned(986, 10), 593 => to_unsigned(493, 10), 594 => to_unsigned(864, 10), 595 => to_unsigned(747, 10), 596 => to_unsigned(961, 10), 597 => to_unsigned(776, 10), 598 => to_unsigned(657, 10), 599 => to_unsigned(590, 10), 600 => to_unsigned(466, 10), 601 => to_unsigned(796, 10), 602 => to_unsigned(465, 10), 603 => to_unsigned(417, 10), 604 => to_unsigned(983, 10), 605 => to_unsigned(980, 10), 606 => to_unsigned(447, 10), 607 => to_unsigned(625, 10), 608 => to_unsigned(458, 10), 609 => to_unsigned(847, 10), 610 => to_unsigned(894, 10), 611 => to_unsigned(473, 10), 612 => to_unsigned(711, 10), 613 => to_unsigned(436, 10), 614 => to_unsigned(200, 10), 615 => to_unsigned(564, 10), 616 => to_unsigned(246, 10), 617 => to_unsigned(151, 10), 618 => to_unsigned(383, 10), 619 => to_unsigned(794, 10), 620 => to_unsigned(98, 10), 621 => to_unsigned(698, 10), 622 => to_unsigned(836, 10), 623 => to_unsigned(473, 10), 624 => to_unsigned(736, 10), 625 => to_unsigned(434, 10), 626 => to_unsigned(763, 10), 627 => to_unsigned(628, 10), 628 => to_unsigned(338, 10), 629 => to_unsigned(990, 10), 630 => to_unsigned(685, 10), 631 => to_unsigned(374, 10), 632 => to_unsigned(48, 10), 633 => to_unsigned(948, 10), 634 => to_unsigned(63, 10), 635 => to_unsigned(606, 10), 636 => to_unsigned(13, 10), 637 => to_unsigned(142, 10), 638 => to_unsigned(955, 10), 639 => to_unsigned(678, 10), 640 => to_unsigned(120, 10), 641 => to_unsigned(630, 10), 642 => to_unsigned(355, 10), 643 => to_unsigned(688, 10), 644 => to_unsigned(436, 10), 645 => to_unsigned(516, 10), 646 => to_unsigned(768, 10), 647 => to_unsigned(560, 10), 648 => to_unsigned(971, 10), 649 => to_unsigned(605, 10), 650 => to_unsigned(374, 10), 651 => to_unsigned(506, 10), 652 => to_unsigned(715, 10), 653 => to_unsigned(50, 10), 654 => to_unsigned(46, 10), 655 => to_unsigned(246, 10), 656 => to_unsigned(510, 10), 657 => to_unsigned(299, 10), 658 => to_unsigned(344, 10), 659 => to_unsigned(723, 10), 660 => to_unsigned(895, 10), 661 => to_unsigned(891, 10), 662 => to_unsigned(168, 10), 663 => to_unsigned(86, 10), 664 => to_unsigned(32, 10), 665 => to_unsigned(686, 10), 666 => to_unsigned(124, 10), 667 => to_unsigned(114, 10), 668 => to_unsigned(780, 10), 669 => to_unsigned(667, 10), 670 => to_unsigned(903, 10), 671 => to_unsigned(372, 10), 672 => to_unsigned(269, 10), 673 => to_unsigned(843, 10), 674 => to_unsigned(386, 10), 675 => to_unsigned(945, 10), 676 => to_unsigned(3, 10), 677 => to_unsigned(796, 10), 678 => to_unsigned(952, 10), 679 => to_unsigned(191, 10), 680 => to_unsigned(53, 10), 681 => to_unsigned(905, 10), 682 => to_unsigned(250, 10), 683 => to_unsigned(685, 10), 684 => to_unsigned(444, 10), 685 => to_unsigned(823, 10), 686 => to_unsigned(412, 10), 687 => to_unsigned(318, 10), 688 => to_unsigned(787, 10), 689 => to_unsigned(1015, 10), 690 => to_unsigned(436, 10), 691 => to_unsigned(727, 10), 692 => to_unsigned(691, 10), 693 => to_unsigned(475, 10), 694 => to_unsigned(869, 10), 695 => to_unsigned(838, 10), 696 => to_unsigned(660, 10), 697 => to_unsigned(79, 10), 698 => to_unsigned(730, 10), 699 => to_unsigned(213, 10), 700 => to_unsigned(764, 10), 701 => to_unsigned(725, 10), 702 => to_unsigned(400, 10), 703 => to_unsigned(515, 10), 704 => to_unsigned(220, 10), 705 => to_unsigned(499, 10), 706 => to_unsigned(884, 10), 707 => to_unsigned(838, 10), 708 => to_unsigned(86, 10), 709 => to_unsigned(27, 10), 710 => to_unsigned(658, 10), 711 => to_unsigned(215, 10), 712 => to_unsigned(90, 10), 713 => to_unsigned(908, 10), 714 => to_unsigned(187, 10), 715 => to_unsigned(124, 10), 716 => to_unsigned(135, 10), 717 => to_unsigned(73, 10), 718 => to_unsigned(771, 10), 719 => to_unsigned(222, 10), 720 => to_unsigned(655, 10), 721 => to_unsigned(263, 10), 722 => to_unsigned(1012, 10), 723 => to_unsigned(217, 10), 724 => to_unsigned(414, 10), 725 => to_unsigned(24, 10), 726 => to_unsigned(241, 10), 727 => to_unsigned(118, 10), 728 => to_unsigned(931, 10), 729 => to_unsigned(163, 10), 730 => to_unsigned(64, 10), 731 => to_unsigned(802, 10), 732 => to_unsigned(582, 10), 733 => to_unsigned(815, 10), 734 => to_unsigned(301, 10), 735 => to_unsigned(515, 10), 736 => to_unsigned(710, 10), 737 => to_unsigned(818, 10), 738 => to_unsigned(248, 10), 739 => to_unsigned(342, 10), 740 => to_unsigned(359, 10), 741 => to_unsigned(504, 10), 742 => to_unsigned(496, 10), 743 => to_unsigned(391, 10), 744 => to_unsigned(797, 10), 745 => to_unsigned(670, 10), 746 => to_unsigned(653, 10), 747 => to_unsigned(259, 10), 748 => to_unsigned(835, 10), 749 => to_unsigned(812, 10), 750 => to_unsigned(434, 10), 751 => to_unsigned(934, 10), 752 => to_unsigned(65, 10), 753 => to_unsigned(994, 10), 754 => to_unsigned(915, 10), 755 => to_unsigned(975, 10), 756 => to_unsigned(118, 10), 757 => to_unsigned(16, 10), 758 => to_unsigned(943, 10), 759 => to_unsigned(855, 10), 760 => to_unsigned(552, 10), 761 => to_unsigned(1015, 10), 762 => to_unsigned(119, 10), 763 => to_unsigned(98, 10), 764 => to_unsigned(15, 10), 765 => to_unsigned(817, 10), 766 => to_unsigned(573, 10), 767 => to_unsigned(226, 10), 768 => to_unsigned(55, 10), 769 => to_unsigned(879, 10), 770 => to_unsigned(715, 10), 771 => to_unsigned(762, 10), 772 => to_unsigned(68, 10), 773 => to_unsigned(413, 10), 774 => to_unsigned(136, 10), 775 => to_unsigned(971, 10), 776 => to_unsigned(976, 10), 777 => to_unsigned(321, 10), 778 => to_unsigned(47, 10), 779 => to_unsigned(209, 10), 780 => to_unsigned(365, 10), 781 => to_unsigned(863, 10), 782 => to_unsigned(616, 10), 783 => to_unsigned(749, 10), 784 => to_unsigned(506, 10), 785 => to_unsigned(117, 10), 786 => to_unsigned(509, 10), 787 => to_unsigned(14, 10), 788 => to_unsigned(766, 10), 789 => to_unsigned(686, 10), 790 => to_unsigned(824, 10), 791 => to_unsigned(1019, 10), 792 => to_unsigned(954, 10), 793 => to_unsigned(625, 10), 794 => to_unsigned(72, 10), 795 => to_unsigned(65, 10), 796 => to_unsigned(347, 10), 797 => to_unsigned(1003, 10), 798 => to_unsigned(713, 10), 799 => to_unsigned(577, 10), 800 => to_unsigned(899, 10), 801 => to_unsigned(688, 10), 802 => to_unsigned(509, 10), 803 => to_unsigned(575, 10), 804 => to_unsigned(686, 10), 805 => to_unsigned(929, 10), 806 => to_unsigned(1, 10), 807 => to_unsigned(291, 10), 808 => to_unsigned(248, 10), 809 => to_unsigned(449, 10), 810 => to_unsigned(737, 10), 811 => to_unsigned(452, 10), 812 => to_unsigned(511, 10), 813 => to_unsigned(922, 10), 814 => to_unsigned(690, 10), 815 => to_unsigned(27, 10), 816 => to_unsigned(370, 10), 817 => to_unsigned(943, 10), 818 => to_unsigned(778, 10), 819 => to_unsigned(660, 10), 820 => to_unsigned(373, 10), 821 => to_unsigned(38, 10), 822 => to_unsigned(472, 10), 823 => to_unsigned(68, 10), 824 => to_unsigned(973, 10), 825 => to_unsigned(858, 10), 826 => to_unsigned(235, 10), 827 => to_unsigned(445, 10), 828 => to_unsigned(165, 10), 829 => to_unsigned(255, 10), 830 => to_unsigned(178, 10), 831 => to_unsigned(586, 10), 832 => to_unsigned(299, 10), 833 => to_unsigned(28, 10), 834 => to_unsigned(427, 10), 835 => to_unsigned(10, 10), 836 => to_unsigned(727, 10), 837 => to_unsigned(574, 10), 838 => to_unsigned(996, 10), 839 => to_unsigned(519, 10), 840 => to_unsigned(879, 10), 841 => to_unsigned(625, 10), 842 => to_unsigned(81, 10), 843 => to_unsigned(692, 10), 844 => to_unsigned(832, 10), 845 => to_unsigned(0, 10), 846 => to_unsigned(330, 10), 847 => to_unsigned(758, 10), 848 => to_unsigned(283, 10), 849 => to_unsigned(769, 10), 850 => to_unsigned(500, 10), 851 => to_unsigned(459, 10), 852 => to_unsigned(506, 10), 853 => to_unsigned(990, 10), 854 => to_unsigned(38, 10), 855 => to_unsigned(123, 10), 856 => to_unsigned(176, 10), 857 => to_unsigned(66, 10), 858 => to_unsigned(799, 10), 859 => to_unsigned(318, 10), 860 => to_unsigned(270, 10), 861 => to_unsigned(75, 10), 862 => to_unsigned(443, 10), 863 => to_unsigned(725, 10), 864 => to_unsigned(694, 10), 865 => to_unsigned(765, 10), 866 => to_unsigned(839, 10), 867 => to_unsigned(588, 10), 868 => to_unsigned(756, 10), 869 => to_unsigned(816, 10), 870 => to_unsigned(683, 10), 871 => to_unsigned(369, 10), 872 => to_unsigned(752, 10), 873 => to_unsigned(5, 10), 874 => to_unsigned(189, 10), 875 => to_unsigned(961, 10), 876 => to_unsigned(161, 10), 877 => to_unsigned(229, 10), 878 => to_unsigned(704, 10), 879 => to_unsigned(44, 10), 880 => to_unsigned(815, 10), 881 => to_unsigned(193, 10), 882 => to_unsigned(530, 10), 883 => to_unsigned(859, 10), 884 => to_unsigned(895, 10), 885 => to_unsigned(626, 10), 886 => to_unsigned(904, 10), 887 => to_unsigned(557, 10), 888 => to_unsigned(755, 10), 889 => to_unsigned(334, 10), 890 => to_unsigned(792, 10), 891 => to_unsigned(1016, 10), 892 => to_unsigned(530, 10), 893 => to_unsigned(9, 10), 894 => to_unsigned(955, 10), 895 => to_unsigned(921, 10), 896 => to_unsigned(830, 10), 897 => to_unsigned(1019, 10), 898 => to_unsigned(153, 10), 899 => to_unsigned(935, 10), 900 => to_unsigned(536, 10), 901 => to_unsigned(756, 10), 902 => to_unsigned(488, 10), 903 => to_unsigned(44, 10), 904 => to_unsigned(513, 10), 905 => to_unsigned(518, 10), 906 => to_unsigned(302, 10), 907 => to_unsigned(299, 10), 908 => to_unsigned(419, 10), 909 => to_unsigned(606, 10), 910 => to_unsigned(497, 10), 911 => to_unsigned(1011, 10), 912 => to_unsigned(751, 10), 913 => to_unsigned(708, 10), 914 => to_unsigned(1004, 10), 915 => to_unsigned(209, 10), 916 => to_unsigned(648, 10), 917 => to_unsigned(628, 10), 918 => to_unsigned(680, 10), 919 => to_unsigned(67, 10), 920 => to_unsigned(870, 10), 921 => to_unsigned(103, 10), 922 => to_unsigned(885, 10), 923 => to_unsigned(1, 10), 924 => to_unsigned(0, 10), 925 => to_unsigned(732, 10), 926 => to_unsigned(815, 10), 927 => to_unsigned(116, 10), 928 => to_unsigned(674, 10), 929 => to_unsigned(145, 10), 930 => to_unsigned(66, 10), 931 => to_unsigned(154, 10), 932 => to_unsigned(548, 10), 933 => to_unsigned(23, 10), 934 => to_unsigned(192, 10), 935 => to_unsigned(222, 10), 936 => to_unsigned(833, 10), 937 => to_unsigned(836, 10), 938 => to_unsigned(982, 10), 939 => to_unsigned(731, 10), 940 => to_unsigned(390, 10), 941 => to_unsigned(381, 10), 942 => to_unsigned(765, 10), 943 => to_unsigned(216, 10), 944 => to_unsigned(981, 10), 945 => to_unsigned(810, 10), 946 => to_unsigned(254, 10), 947 => to_unsigned(747, 10), 948 => to_unsigned(122, 10), 949 => to_unsigned(311, 10), 950 => to_unsigned(756, 10), 951 => to_unsigned(516, 10), 952 => to_unsigned(419, 10), 953 => to_unsigned(935, 10), 954 => to_unsigned(355, 10), 955 => to_unsigned(897, 10), 956 => to_unsigned(1002, 10), 957 => to_unsigned(168, 10), 958 => to_unsigned(791, 10), 959 => to_unsigned(681, 10), 960 => to_unsigned(131, 10), 961 => to_unsigned(252, 10), 962 => to_unsigned(28, 10), 963 => to_unsigned(770, 10), 964 => to_unsigned(431, 10), 965 => to_unsigned(601, 10), 966 => to_unsigned(727, 10), 967 => to_unsigned(611, 10), 968 => to_unsigned(728, 10), 969 => to_unsigned(430, 10), 970 => to_unsigned(759, 10), 971 => to_unsigned(861, 10), 972 => to_unsigned(382, 10), 973 => to_unsigned(312, 10), 974 => to_unsigned(105, 10), 975 => to_unsigned(574, 10), 976 => to_unsigned(677, 10), 977 => to_unsigned(319, 10), 978 => to_unsigned(141, 10), 979 => to_unsigned(148, 10), 980 => to_unsigned(505, 10), 981 => to_unsigned(402, 10), 982 => to_unsigned(293, 10), 983 => to_unsigned(134, 10), 984 => to_unsigned(87, 10), 985 => to_unsigned(522, 10), 986 => to_unsigned(186, 10), 987 => to_unsigned(740, 10), 988 => to_unsigned(577, 10), 989 => to_unsigned(940, 10), 990 => to_unsigned(629, 10), 991 => to_unsigned(360, 10), 992 => to_unsigned(595, 10), 993 => to_unsigned(911, 10), 994 => to_unsigned(203, 10), 995 => to_unsigned(639, 10), 996 => to_unsigned(201, 10), 997 => to_unsigned(1004, 10), 998 => to_unsigned(465, 10), 999 => to_unsigned(554, 10), 1000 => to_unsigned(937, 10), 1001 => to_unsigned(793, 10), 1002 => to_unsigned(580, 10), 1003 => to_unsigned(975, 10), 1004 => to_unsigned(898, 10), 1005 => to_unsigned(255, 10), 1006 => to_unsigned(89, 10), 1007 => to_unsigned(519, 10), 1008 => to_unsigned(631, 10), 1009 => to_unsigned(575, 10), 1010 => to_unsigned(618, 10), 1011 => to_unsigned(17, 10), 1012 => to_unsigned(880, 10), 1013 => to_unsigned(380, 10), 1014 => to_unsigned(522, 10), 1015 => to_unsigned(675, 10), 1016 => to_unsigned(933, 10), 1017 => to_unsigned(766, 10), 1018 => to_unsigned(855, 10), 1019 => to_unsigned(809, 10), 1020 => to_unsigned(367, 10), 1021 => to_unsigned(477, 10), 1022 => to_unsigned(890, 10), 1023 => to_unsigned(815, 10), 1024 => to_unsigned(252, 10), 1025 => to_unsigned(174, 10), 1026 => to_unsigned(549, 10), 1027 => to_unsigned(681, 10), 1028 => to_unsigned(167, 10), 1029 => to_unsigned(934, 10), 1030 => to_unsigned(367, 10), 1031 => to_unsigned(889, 10), 1032 => to_unsigned(464, 10), 1033 => to_unsigned(436, 10), 1034 => to_unsigned(989, 10), 1035 => to_unsigned(18, 10), 1036 => to_unsigned(235, 10), 1037 => to_unsigned(48, 10), 1038 => to_unsigned(343, 10), 1039 => to_unsigned(645, 10), 1040 => to_unsigned(375, 10), 1041 => to_unsigned(504, 10), 1042 => to_unsigned(571, 10), 1043 => to_unsigned(182, 10), 1044 => to_unsigned(1014, 10), 1045 => to_unsigned(555, 10), 1046 => to_unsigned(877, 10), 1047 => to_unsigned(524, 10), 1048 => to_unsigned(27, 10), 1049 => to_unsigned(911, 10), 1050 => to_unsigned(411, 10), 1051 => to_unsigned(109, 10), 1052 => to_unsigned(912, 10), 1053 => to_unsigned(698, 10), 1054 => to_unsigned(817, 10), 1055 => to_unsigned(486, 10), 1056 => to_unsigned(442, 10), 1057 => to_unsigned(287, 10), 1058 => to_unsigned(434, 10), 1059 => to_unsigned(388, 10), 1060 => to_unsigned(408, 10), 1061 => to_unsigned(664, 10), 1062 => to_unsigned(972, 10), 1063 => to_unsigned(694, 10), 1064 => to_unsigned(110, 10), 1065 => to_unsigned(801, 10), 1066 => to_unsigned(379, 10), 1067 => to_unsigned(641, 10), 1068 => to_unsigned(76, 10), 1069 => to_unsigned(835, 10), 1070 => to_unsigned(89, 10), 1071 => to_unsigned(559, 10), 1072 => to_unsigned(402, 10), 1073 => to_unsigned(180, 10), 1074 => to_unsigned(147, 10), 1075 => to_unsigned(347, 10), 1076 => to_unsigned(593, 10), 1077 => to_unsigned(863, 10), 1078 => to_unsigned(795, 10), 1079 => to_unsigned(20, 10), 1080 => to_unsigned(885, 10), 1081 => to_unsigned(670, 10), 1082 => to_unsigned(1010, 10), 1083 => to_unsigned(429, 10), 1084 => to_unsigned(850, 10), 1085 => to_unsigned(498, 10), 1086 => to_unsigned(137, 10), 1087 => to_unsigned(209, 10), 1088 => to_unsigned(216, 10), 1089 => to_unsigned(96, 10), 1090 => to_unsigned(571, 10), 1091 => to_unsigned(527, 10), 1092 => to_unsigned(117, 10), 1093 => to_unsigned(726, 10), 1094 => to_unsigned(382, 10), 1095 => to_unsigned(652, 10), 1096 => to_unsigned(509, 10), 1097 => to_unsigned(294, 10), 1098 => to_unsigned(621, 10), 1099 => to_unsigned(97, 10), 1100 => to_unsigned(135, 10), 1101 => to_unsigned(259, 10), 1102 => to_unsigned(595, 10), 1103 => to_unsigned(816, 10), 1104 => to_unsigned(716, 10), 1105 => to_unsigned(677, 10), 1106 => to_unsigned(57, 10), 1107 => to_unsigned(747, 10), 1108 => to_unsigned(217, 10), 1109 => to_unsigned(440, 10), 1110 => to_unsigned(313, 10), 1111 => to_unsigned(908, 10), 1112 => to_unsigned(894, 10), 1113 => to_unsigned(312, 10), 1114 => to_unsigned(181, 10), 1115 => to_unsigned(239, 10), 1116 => to_unsigned(917, 10), 1117 => to_unsigned(496, 10), 1118 => to_unsigned(761, 10), 1119 => to_unsigned(307, 10), 1120 => to_unsigned(771, 10), 1121 => to_unsigned(605, 10), 1122 => to_unsigned(463, 10), 1123 => to_unsigned(969, 10), 1124 => to_unsigned(600, 10), 1125 => to_unsigned(508, 10), 1126 => to_unsigned(823, 10), 1127 => to_unsigned(386, 10), 1128 => to_unsigned(365, 10), 1129 => to_unsigned(339, 10), 1130 => to_unsigned(535, 10), 1131 => to_unsigned(277, 10), 1132 => to_unsigned(571, 10), 1133 => to_unsigned(602, 10), 1134 => to_unsigned(106, 10), 1135 => to_unsigned(49, 10), 1136 => to_unsigned(214, 10), 1137 => to_unsigned(490, 10), 1138 => to_unsigned(995, 10), 1139 => to_unsigned(843, 10), 1140 => to_unsigned(258, 10), 1141 => to_unsigned(945, 10), 1142 => to_unsigned(876, 10), 1143 => to_unsigned(724, 10), 1144 => to_unsigned(907, 10), 1145 => to_unsigned(819, 10), 1146 => to_unsigned(1003, 10), 1147 => to_unsigned(630, 10), 1148 => to_unsigned(165, 10), 1149 => to_unsigned(11, 10), 1150 => to_unsigned(411, 10), 1151 => to_unsigned(880, 10), 1152 => to_unsigned(500, 10), 1153 => to_unsigned(704, 10), 1154 => to_unsigned(754, 10), 1155 => to_unsigned(675, 10), 1156 => to_unsigned(192, 10), 1157 => to_unsigned(172, 10), 1158 => to_unsigned(995, 10), 1159 => to_unsigned(26, 10), 1160 => to_unsigned(747, 10), 1161 => to_unsigned(992, 10), 1162 => to_unsigned(492, 10), 1163 => to_unsigned(845, 10), 1164 => to_unsigned(253, 10), 1165 => to_unsigned(761, 10), 1166 => to_unsigned(200, 10), 1167 => to_unsigned(435, 10), 1168 => to_unsigned(179, 10), 1169 => to_unsigned(59, 10), 1170 => to_unsigned(144, 10), 1171 => to_unsigned(446, 10), 1172 => to_unsigned(135, 10), 1173 => to_unsigned(831, 10), 1174 => to_unsigned(691, 10), 1175 => to_unsigned(584, 10), 1176 => to_unsigned(384, 10), 1177 => to_unsigned(270, 10), 1178 => to_unsigned(953, 10), 1179 => to_unsigned(264, 10), 1180 => to_unsigned(426, 10), 1181 => to_unsigned(987, 10), 1182 => to_unsigned(871, 10), 1183 => to_unsigned(116, 10), 1184 => to_unsigned(20, 10), 1185 => to_unsigned(674, 10), 1186 => to_unsigned(152, 10), 1187 => to_unsigned(2, 10), 1188 => to_unsigned(193, 10), 1189 => to_unsigned(535, 10), 1190 => to_unsigned(95, 10), 1191 => to_unsigned(170, 10), 1192 => to_unsigned(28, 10), 1193 => to_unsigned(680, 10), 1194 => to_unsigned(855, 10), 1195 => to_unsigned(801, 10), 1196 => to_unsigned(500, 10), 1197 => to_unsigned(730, 10), 1198 => to_unsigned(716, 10), 1199 => to_unsigned(463, 10), 1200 => to_unsigned(20, 10), 1201 => to_unsigned(686, 10), 1202 => to_unsigned(991, 10), 1203 => to_unsigned(830, 10), 1204 => to_unsigned(762, 10), 1205 => to_unsigned(139, 10), 1206 => to_unsigned(355, 10), 1207 => to_unsigned(292, 10), 1208 => to_unsigned(460, 10), 1209 => to_unsigned(921, 10), 1210 => to_unsigned(20, 10), 1211 => to_unsigned(526, 10), 1212 => to_unsigned(893, 10), 1213 => to_unsigned(47, 10), 1214 => to_unsigned(413, 10), 1215 => to_unsigned(718, 10), 1216 => to_unsigned(735, 10), 1217 => to_unsigned(971, 10), 1218 => to_unsigned(623, 10), 1219 => to_unsigned(409, 10), 1220 => to_unsigned(347, 10), 1221 => to_unsigned(583, 10), 1222 => to_unsigned(204, 10), 1223 => to_unsigned(256, 10), 1224 => to_unsigned(733, 10), 1225 => to_unsigned(149, 10), 1226 => to_unsigned(646, 10), 1227 => to_unsigned(438, 10), 1228 => to_unsigned(761, 10), 1229 => to_unsigned(672, 10), 1230 => to_unsigned(559, 10), 1231 => to_unsigned(471, 10), 1232 => to_unsigned(326, 10), 1233 => to_unsigned(994, 10), 1234 => to_unsigned(852, 10), 1235 => to_unsigned(899, 10), 1236 => to_unsigned(929, 10), 1237 => to_unsigned(834, 10), 1238 => to_unsigned(681, 10), 1239 => to_unsigned(709, 10), 1240 => to_unsigned(964, 10), 1241 => to_unsigned(155, 10), 1242 => to_unsigned(908, 10), 1243 => to_unsigned(721, 10), 1244 => to_unsigned(791, 10), 1245 => to_unsigned(502, 10), 1246 => to_unsigned(714, 10), 1247 => to_unsigned(762, 10), 1248 => to_unsigned(695, 10), 1249 => to_unsigned(337, 10), 1250 => to_unsigned(762, 10), 1251 => to_unsigned(726, 10), 1252 => to_unsigned(164, 10), 1253 => to_unsigned(234, 10), 1254 => to_unsigned(32, 10), 1255 => to_unsigned(277, 10), 1256 => to_unsigned(760, 10), 1257 => to_unsigned(728, 10), 1258 => to_unsigned(804, 10), 1259 => to_unsigned(513, 10), 1260 => to_unsigned(119, 10), 1261 => to_unsigned(533, 10), 1262 => to_unsigned(334, 10), 1263 => to_unsigned(944, 10), 1264 => to_unsigned(876, 10), 1265 => to_unsigned(515, 10), 1266 => to_unsigned(403, 10), 1267 => to_unsigned(305, 10), 1268 => to_unsigned(398, 10), 1269 => to_unsigned(554, 10), 1270 => to_unsigned(570, 10), 1271 => to_unsigned(625, 10), 1272 => to_unsigned(759, 10), 1273 => to_unsigned(486, 10), 1274 => to_unsigned(910, 10), 1275 => to_unsigned(933, 10), 1276 => to_unsigned(711, 10), 1277 => to_unsigned(702, 10), 1278 => to_unsigned(565, 10), 1279 => to_unsigned(853, 10), 1280 => to_unsigned(804, 10), 1281 => to_unsigned(958, 10), 1282 => to_unsigned(134, 10), 1283 => to_unsigned(806, 10), 1284 => to_unsigned(274, 10), 1285 => to_unsigned(841, 10), 1286 => to_unsigned(357, 10), 1287 => to_unsigned(230, 10), 1288 => to_unsigned(59, 10), 1289 => to_unsigned(729, 10), 1290 => to_unsigned(951, 10), 1291 => to_unsigned(199, 10), 1292 => to_unsigned(602, 10), 1293 => to_unsigned(471, 10), 1294 => to_unsigned(147, 10), 1295 => to_unsigned(979, 10), 1296 => to_unsigned(773, 10), 1297 => to_unsigned(823, 10), 1298 => to_unsigned(308, 10), 1299 => to_unsigned(315, 10), 1300 => to_unsigned(508, 10), 1301 => to_unsigned(38, 10), 1302 => to_unsigned(427, 10), 1303 => to_unsigned(503, 10), 1304 => to_unsigned(281, 10), 1305 => to_unsigned(358, 10), 1306 => to_unsigned(53, 10), 1307 => to_unsigned(635, 10), 1308 => to_unsigned(642, 10), 1309 => to_unsigned(531, 10), 1310 => to_unsigned(47, 10), 1311 => to_unsigned(394, 10), 1312 => to_unsigned(238, 10), 1313 => to_unsigned(960, 10), 1314 => to_unsigned(987, 10), 1315 => to_unsigned(578, 10), 1316 => to_unsigned(181, 10), 1317 => to_unsigned(148, 10), 1318 => to_unsigned(764, 10), 1319 => to_unsigned(198, 10), 1320 => to_unsigned(428, 10), 1321 => to_unsigned(127, 10), 1322 => to_unsigned(811, 10), 1323 => to_unsigned(432, 10), 1324 => to_unsigned(747, 10), 1325 => to_unsigned(992, 10), 1326 => to_unsigned(365, 10), 1327 => to_unsigned(144, 10), 1328 => to_unsigned(383, 10), 1329 => to_unsigned(871, 10), 1330 => to_unsigned(617, 10), 1331 => to_unsigned(189, 10), 1332 => to_unsigned(196, 10), 1333 => to_unsigned(375, 10), 1334 => to_unsigned(403, 10), 1335 => to_unsigned(496, 10), 1336 => to_unsigned(904, 10), 1337 => to_unsigned(498, 10), 1338 => to_unsigned(976, 10), 1339 => to_unsigned(993, 10), 1340 => to_unsigned(437, 10), 1341 => to_unsigned(441, 10), 1342 => to_unsigned(656, 10), 1343 => to_unsigned(544, 10), 1344 => to_unsigned(354, 10), 1345 => to_unsigned(850, 10), 1346 => to_unsigned(669, 10), 1347 => to_unsigned(1004, 10), 1348 => to_unsigned(627, 10), 1349 => to_unsigned(279, 10), 1350 => to_unsigned(502, 10), 1351 => to_unsigned(702, 10), 1352 => to_unsigned(207, 10), 1353 => to_unsigned(230, 10), 1354 => to_unsigned(340, 10), 1355 => to_unsigned(798, 10), 1356 => to_unsigned(750, 10), 1357 => to_unsigned(442, 10), 1358 => to_unsigned(598, 10), 1359 => to_unsigned(1018, 10), 1360 => to_unsigned(732, 10), 1361 => to_unsigned(711, 10), 1362 => to_unsigned(741, 10), 1363 => to_unsigned(434, 10), 1364 => to_unsigned(117, 10), 1365 => to_unsigned(701, 10), 1366 => to_unsigned(813, 10), 1367 => to_unsigned(150, 10), 1368 => to_unsigned(568, 10), 1369 => to_unsigned(768, 10), 1370 => to_unsigned(512, 10), 1371 => to_unsigned(936, 10), 1372 => to_unsigned(680, 10), 1373 => to_unsigned(853, 10), 1374 => to_unsigned(220, 10), 1375 => to_unsigned(73, 10), 1376 => to_unsigned(267, 10), 1377 => to_unsigned(825, 10), 1378 => to_unsigned(990, 10), 1379 => to_unsigned(336, 10), 1380 => to_unsigned(448, 10), 1381 => to_unsigned(670, 10), 1382 => to_unsigned(173, 10), 1383 => to_unsigned(329, 10), 1384 => to_unsigned(450, 10), 1385 => to_unsigned(782, 10), 1386 => to_unsigned(140, 10), 1387 => to_unsigned(169, 10), 1388 => to_unsigned(14, 10), 1389 => to_unsigned(612, 10), 1390 => to_unsigned(811, 10), 1391 => to_unsigned(870, 10), 1392 => to_unsigned(201, 10), 1393 => to_unsigned(139, 10), 1394 => to_unsigned(382, 10), 1395 => to_unsigned(508, 10), 1396 => to_unsigned(858, 10), 1397 => to_unsigned(467, 10), 1398 => to_unsigned(54, 10), 1399 => to_unsigned(303, 10), 1400 => to_unsigned(555, 10), 1401 => to_unsigned(970, 10), 1402 => to_unsigned(148, 10), 1403 => to_unsigned(233, 10), 1404 => to_unsigned(1008, 10), 1405 => to_unsigned(52, 10), 1406 => to_unsigned(544, 10), 1407 => to_unsigned(915, 10), 1408 => to_unsigned(492, 10), 1409 => to_unsigned(873, 10), 1410 => to_unsigned(873, 10), 1411 => to_unsigned(350, 10), 1412 => to_unsigned(592, 10), 1413 => to_unsigned(410, 10), 1414 => to_unsigned(553, 10), 1415 => to_unsigned(1010, 10), 1416 => to_unsigned(822, 10), 1417 => to_unsigned(356, 10), 1418 => to_unsigned(592, 10), 1419 => to_unsigned(520, 10), 1420 => to_unsigned(886, 10), 1421 => to_unsigned(326, 10), 1422 => to_unsigned(21, 10), 1423 => to_unsigned(891, 10), 1424 => to_unsigned(727, 10), 1425 => to_unsigned(612, 10), 1426 => to_unsigned(156, 10), 1427 => to_unsigned(816, 10), 1428 => to_unsigned(329, 10), 1429 => to_unsigned(931, 10), 1430 => to_unsigned(382, 10), 1431 => to_unsigned(631, 10), 1432 => to_unsigned(285, 10), 1433 => to_unsigned(122, 10), 1434 => to_unsigned(686, 10), 1435 => to_unsigned(430, 10), 1436 => to_unsigned(815, 10), 1437 => to_unsigned(371, 10), 1438 => to_unsigned(991, 10), 1439 => to_unsigned(498, 10), 1440 => to_unsigned(712, 10), 1441 => to_unsigned(305, 10), 1442 => to_unsigned(481, 10), 1443 => to_unsigned(188, 10), 1444 => to_unsigned(774, 10), 1445 => to_unsigned(41, 10), 1446 => to_unsigned(999, 10), 1447 => to_unsigned(227, 10), 1448 => to_unsigned(738, 10), 1449 => to_unsigned(726, 10), 1450 => to_unsigned(878, 10), 1451 => to_unsigned(926, 10), 1452 => to_unsigned(768, 10), 1453 => to_unsigned(295, 10), 1454 => to_unsigned(121, 10), 1455 => to_unsigned(966, 10), 1456 => to_unsigned(78, 10), 1457 => to_unsigned(175, 10), 1458 => to_unsigned(727, 10), 1459 => to_unsigned(342, 10), 1460 => to_unsigned(615, 10), 1461 => to_unsigned(71, 10), 1462 => to_unsigned(683, 10), 1463 => to_unsigned(695, 10), 1464 => to_unsigned(26, 10), 1465 => to_unsigned(327, 10), 1466 => to_unsigned(632, 10), 1467 => to_unsigned(175, 10), 1468 => to_unsigned(6, 10), 1469 => to_unsigned(701, 10), 1470 => to_unsigned(552, 10), 1471 => to_unsigned(798, 10), 1472 => to_unsigned(740, 10), 1473 => to_unsigned(647, 10), 1474 => to_unsigned(139, 10), 1475 => to_unsigned(948, 10), 1476 => to_unsigned(539, 10), 1477 => to_unsigned(18, 10), 1478 => to_unsigned(849, 10), 1479 => to_unsigned(394, 10), 1480 => to_unsigned(404, 10), 1481 => to_unsigned(177, 10), 1482 => to_unsigned(705, 10), 1483 => to_unsigned(917, 10), 1484 => to_unsigned(318, 10), 1485 => to_unsigned(92, 10), 1486 => to_unsigned(233, 10), 1487 => to_unsigned(198, 10), 1488 => to_unsigned(956, 10), 1489 => to_unsigned(818, 10), 1490 => to_unsigned(412, 10), 1491 => to_unsigned(66, 10), 1492 => to_unsigned(1023, 10), 1493 => to_unsigned(842, 10), 1494 => to_unsigned(617, 10), 1495 => to_unsigned(886, 10), 1496 => to_unsigned(28, 10), 1497 => to_unsigned(592, 10), 1498 => to_unsigned(164, 10), 1499 => to_unsigned(638, 10), 1500 => to_unsigned(873, 10), 1501 => to_unsigned(432, 10), 1502 => to_unsigned(375, 10), 1503 => to_unsigned(349, 10), 1504 => to_unsigned(658, 10), 1505 => to_unsigned(641, 10), 1506 => to_unsigned(110, 10), 1507 => to_unsigned(210, 10), 1508 => to_unsigned(814, 10), 1509 => to_unsigned(826, 10), 1510 => to_unsigned(425, 10), 1511 => to_unsigned(976, 10), 1512 => to_unsigned(339, 10), 1513 => to_unsigned(966, 10), 1514 => to_unsigned(351, 10), 1515 => to_unsigned(10, 10), 1516 => to_unsigned(30, 10), 1517 => to_unsigned(500, 10), 1518 => to_unsigned(991, 10), 1519 => to_unsigned(227, 10), 1520 => to_unsigned(918, 10), 1521 => to_unsigned(138, 10), 1522 => to_unsigned(875, 10), 1523 => to_unsigned(141, 10), 1524 => to_unsigned(736, 10), 1525 => to_unsigned(654, 10), 1526 => to_unsigned(312, 10), 1527 => to_unsigned(269, 10), 1528 => to_unsigned(486, 10), 1529 => to_unsigned(160, 10), 1530 => to_unsigned(936, 10), 1531 => to_unsigned(803, 10), 1532 => to_unsigned(945, 10), 1533 => to_unsigned(411, 10), 1534 => to_unsigned(604, 10), 1535 => to_unsigned(1004, 10), 1536 => to_unsigned(986, 10), 1537 => to_unsigned(908, 10), 1538 => to_unsigned(223, 10), 1539 => to_unsigned(563, 10), 1540 => to_unsigned(33, 10), 1541 => to_unsigned(312, 10), 1542 => to_unsigned(814, 10), 1543 => to_unsigned(325, 10), 1544 => to_unsigned(1005, 10), 1545 => to_unsigned(635, 10), 1546 => to_unsigned(315, 10), 1547 => to_unsigned(724, 10), 1548 => to_unsigned(144, 10), 1549 => to_unsigned(295, 10), 1550 => to_unsigned(803, 10), 1551 => to_unsigned(408, 10), 1552 => to_unsigned(922, 10), 1553 => to_unsigned(775, 10), 1554 => to_unsigned(164, 10), 1555 => to_unsigned(613, 10), 1556 => to_unsigned(792, 10), 1557 => to_unsigned(466, 10), 1558 => to_unsigned(157, 10), 1559 => to_unsigned(154, 10), 1560 => to_unsigned(855, 10), 1561 => to_unsigned(942, 10), 1562 => to_unsigned(43, 10), 1563 => to_unsigned(150, 10), 1564 => to_unsigned(301, 10), 1565 => to_unsigned(427, 10), 1566 => to_unsigned(130, 10), 1567 => to_unsigned(209, 10), 1568 => to_unsigned(61, 10), 1569 => to_unsigned(448, 10), 1570 => to_unsigned(352, 10), 1571 => to_unsigned(555, 10), 1572 => to_unsigned(516, 10), 1573 => to_unsigned(422, 10), 1574 => to_unsigned(668, 10), 1575 => to_unsigned(58, 10), 1576 => to_unsigned(546, 10), 1577 => to_unsigned(157, 10), 1578 => to_unsigned(808, 10), 1579 => to_unsigned(492, 10), 1580 => to_unsigned(377, 10), 1581 => to_unsigned(144, 10), 1582 => to_unsigned(158, 10), 1583 => to_unsigned(255, 10), 1584 => to_unsigned(8, 10), 1585 => to_unsigned(812, 10), 1586 => to_unsigned(354, 10), 1587 => to_unsigned(833, 10), 1588 => to_unsigned(151, 10), 1589 => to_unsigned(635, 10), 1590 => to_unsigned(861, 10), 1591 => to_unsigned(852, 10), 1592 => to_unsigned(965, 10), 1593 => to_unsigned(925, 10), 1594 => to_unsigned(169, 10), 1595 => to_unsigned(957, 10), 1596 => to_unsigned(448, 10), 1597 => to_unsigned(807, 10), 1598 => to_unsigned(593, 10), 1599 => to_unsigned(23, 10), 1600 => to_unsigned(219, 10), 1601 => to_unsigned(908, 10), 1602 => to_unsigned(691, 10), 1603 => to_unsigned(727, 10), 1604 => to_unsigned(465, 10), 1605 => to_unsigned(347, 10), 1606 => to_unsigned(987, 10), 1607 => to_unsigned(876, 10), 1608 => to_unsigned(198, 10), 1609 => to_unsigned(820, 10), 1610 => to_unsigned(947, 10), 1611 => to_unsigned(202, 10), 1612 => to_unsigned(175, 10), 1613 => to_unsigned(9, 10), 1614 => to_unsigned(609, 10), 1615 => to_unsigned(49, 10), 1616 => to_unsigned(956, 10), 1617 => to_unsigned(331, 10), 1618 => to_unsigned(885, 10), 1619 => to_unsigned(796, 10), 1620 => to_unsigned(322, 10), 1621 => to_unsigned(697, 10), 1622 => to_unsigned(885, 10), 1623 => to_unsigned(134, 10), 1624 => to_unsigned(929, 10), 1625 => to_unsigned(139, 10), 1626 => to_unsigned(307, 10), 1627 => to_unsigned(475, 10), 1628 => to_unsigned(407, 10), 1629 => to_unsigned(719, 10), 1630 => to_unsigned(160, 10), 1631 => to_unsigned(196, 10), 1632 => to_unsigned(601, 10), 1633 => to_unsigned(743, 10), 1634 => to_unsigned(110, 10), 1635 => to_unsigned(952, 10), 1636 => to_unsigned(271, 10), 1637 => to_unsigned(472, 10), 1638 => to_unsigned(162, 10), 1639 => to_unsigned(674, 10), 1640 => to_unsigned(42, 10), 1641 => to_unsigned(24, 10), 1642 => to_unsigned(752, 10), 1643 => to_unsigned(539, 10), 1644 => to_unsigned(290, 10), 1645 => to_unsigned(922, 10), 1646 => to_unsigned(612, 10), 1647 => to_unsigned(602, 10), 1648 => to_unsigned(1018, 10), 1649 => to_unsigned(501, 10), 1650 => to_unsigned(638, 10), 1651 => to_unsigned(493, 10), 1652 => to_unsigned(427, 10), 1653 => to_unsigned(37, 10), 1654 => to_unsigned(120, 10), 1655 => to_unsigned(738, 10), 1656 => to_unsigned(612, 10), 1657 => to_unsigned(51, 10), 1658 => to_unsigned(55, 10), 1659 => to_unsigned(755, 10), 1660 => to_unsigned(235, 10), 1661 => to_unsigned(972, 10), 1662 => to_unsigned(296, 10), 1663 => to_unsigned(941, 10), 1664 => to_unsigned(275, 10), 1665 => to_unsigned(660, 10), 1666 => to_unsigned(970, 10), 1667 => to_unsigned(791, 10), 1668 => to_unsigned(470, 10), 1669 => to_unsigned(950, 10), 1670 => to_unsigned(450, 10), 1671 => to_unsigned(315, 10), 1672 => to_unsigned(127, 10), 1673 => to_unsigned(544, 10), 1674 => to_unsigned(691, 10), 1675 => to_unsigned(946, 10), 1676 => to_unsigned(992, 10), 1677 => to_unsigned(424, 10), 1678 => to_unsigned(362, 10), 1679 => to_unsigned(370, 10), 1680 => to_unsigned(888, 10), 1681 => to_unsigned(258, 10), 1682 => to_unsigned(82, 10), 1683 => to_unsigned(317, 10), 1684 => to_unsigned(84, 10), 1685 => to_unsigned(303, 10), 1686 => to_unsigned(250, 10), 1687 => to_unsigned(718, 10), 1688 => to_unsigned(727, 10), 1689 => to_unsigned(206, 10), 1690 => to_unsigned(1013, 10), 1691 => to_unsigned(823, 10), 1692 => to_unsigned(307, 10), 1693 => to_unsigned(821, 10), 1694 => to_unsigned(282, 10), 1695 => to_unsigned(831, 10), 1696 => to_unsigned(967, 10), 1697 => to_unsigned(319, 10), 1698 => to_unsigned(402, 10), 1699 => to_unsigned(233, 10), 1700 => to_unsigned(319, 10), 1701 => to_unsigned(150, 10), 1702 => to_unsigned(796, 10), 1703 => to_unsigned(443, 10), 1704 => to_unsigned(734, 10), 1705 => to_unsigned(516, 10), 1706 => to_unsigned(367, 10), 1707 => to_unsigned(632, 10), 1708 => to_unsigned(1003, 10), 1709 => to_unsigned(319, 10), 1710 => to_unsigned(364, 10), 1711 => to_unsigned(671, 10), 1712 => to_unsigned(105, 10), 1713 => to_unsigned(660, 10), 1714 => to_unsigned(689, 10), 1715 => to_unsigned(294, 10), 1716 => to_unsigned(731, 10), 1717 => to_unsigned(198, 10), 1718 => to_unsigned(105, 10), 1719 => to_unsigned(1022, 10), 1720 => to_unsigned(518, 10), 1721 => to_unsigned(418, 10), 1722 => to_unsigned(204, 10), 1723 => to_unsigned(971, 10), 1724 => to_unsigned(865, 10), 1725 => to_unsigned(310, 10), 1726 => to_unsigned(681, 10), 1727 => to_unsigned(324, 10), 1728 => to_unsigned(817, 10), 1729 => to_unsigned(791, 10), 1730 => to_unsigned(148, 10), 1731 => to_unsigned(897, 10), 1732 => to_unsigned(236, 10), 1733 => to_unsigned(654, 10), 1734 => to_unsigned(1022, 10), 1735 => to_unsigned(694, 10), 1736 => to_unsigned(136, 10), 1737 => to_unsigned(88, 10), 1738 => to_unsigned(252, 10), 1739 => to_unsigned(309, 10), 1740 => to_unsigned(464, 10), 1741 => to_unsigned(488, 10), 1742 => to_unsigned(994, 10), 1743 => to_unsigned(746, 10), 1744 => to_unsigned(537, 10), 1745 => to_unsigned(747, 10), 1746 => to_unsigned(699, 10), 1747 => to_unsigned(310, 10), 1748 => to_unsigned(500, 10), 1749 => to_unsigned(535, 10), 1750 => to_unsigned(0, 10), 1751 => to_unsigned(634, 10), 1752 => to_unsigned(180, 10), 1753 => to_unsigned(90, 10), 1754 => to_unsigned(8, 10), 1755 => to_unsigned(413, 10), 1756 => to_unsigned(794, 10), 1757 => to_unsigned(925, 10), 1758 => to_unsigned(552, 10), 1759 => to_unsigned(271, 10), 1760 => to_unsigned(257, 10), 1761 => to_unsigned(190, 10), 1762 => to_unsigned(585, 10), 1763 => to_unsigned(25, 10), 1764 => to_unsigned(379, 10), 1765 => to_unsigned(44, 10), 1766 => to_unsigned(283, 10), 1767 => to_unsigned(78, 10), 1768 => to_unsigned(881, 10), 1769 => to_unsigned(543, 10), 1770 => to_unsigned(241, 10), 1771 => to_unsigned(928, 10), 1772 => to_unsigned(767, 10), 1773 => to_unsigned(967, 10), 1774 => to_unsigned(39, 10), 1775 => to_unsigned(635, 10), 1776 => to_unsigned(10, 10), 1777 => to_unsigned(750, 10), 1778 => to_unsigned(937, 10), 1779 => to_unsigned(129, 10), 1780 => to_unsigned(542, 10), 1781 => to_unsigned(927, 10), 1782 => to_unsigned(42, 10), 1783 => to_unsigned(947, 10), 1784 => to_unsigned(375, 10), 1785 => to_unsigned(460, 10), 1786 => to_unsigned(709, 10), 1787 => to_unsigned(672, 10), 1788 => to_unsigned(481, 10), 1789 => to_unsigned(271, 10), 1790 => to_unsigned(814, 10), 1791 => to_unsigned(547, 10), 1792 => to_unsigned(313, 10), 1793 => to_unsigned(500, 10), 1794 => to_unsigned(230, 10), 1795 => to_unsigned(862, 10), 1796 => to_unsigned(581, 10), 1797 => to_unsigned(857, 10), 1798 => to_unsigned(677, 10), 1799 => to_unsigned(791, 10), 1800 => to_unsigned(949, 10), 1801 => to_unsigned(317, 10), 1802 => to_unsigned(920, 10), 1803 => to_unsigned(179, 10), 1804 => to_unsigned(662, 10), 1805 => to_unsigned(502, 10), 1806 => to_unsigned(838, 10), 1807 => to_unsigned(916, 10), 1808 => to_unsigned(209, 10), 1809 => to_unsigned(190, 10), 1810 => to_unsigned(88, 10), 1811 => to_unsigned(482, 10), 1812 => to_unsigned(65, 10), 1813 => to_unsigned(39, 10), 1814 => to_unsigned(171, 10), 1815 => to_unsigned(151, 10), 1816 => to_unsigned(795, 10), 1817 => to_unsigned(928, 10), 1818 => to_unsigned(985, 10), 1819 => to_unsigned(320, 10), 1820 => to_unsigned(499, 10), 1821 => to_unsigned(536, 10), 1822 => to_unsigned(869, 10), 1823 => to_unsigned(343, 10), 1824 => to_unsigned(241, 10), 1825 => to_unsigned(849, 10), 1826 => to_unsigned(254, 10), 1827 => to_unsigned(861, 10), 1828 => to_unsigned(436, 10), 1829 => to_unsigned(771, 10), 1830 => to_unsigned(757, 10), 1831 => to_unsigned(1010, 10), 1832 => to_unsigned(972, 10), 1833 => to_unsigned(483, 10), 1834 => to_unsigned(675, 10), 1835 => to_unsigned(810, 10), 1836 => to_unsigned(598, 10), 1837 => to_unsigned(124, 10), 1838 => to_unsigned(222, 10), 1839 => to_unsigned(582, 10), 1840 => to_unsigned(574, 10), 1841 => to_unsigned(57, 10), 1842 => to_unsigned(173, 10), 1843 => to_unsigned(200, 10), 1844 => to_unsigned(441, 10), 1845 => to_unsigned(239, 10), 1846 => to_unsigned(144, 10), 1847 => to_unsigned(198, 10), 1848 => to_unsigned(138, 10), 1849 => to_unsigned(332, 10), 1850 => to_unsigned(1018, 10), 1851 => to_unsigned(583, 10), 1852 => to_unsigned(968, 10), 1853 => to_unsigned(445, 10), 1854 => to_unsigned(93, 10), 1855 => to_unsigned(966, 10), 1856 => to_unsigned(775, 10), 1857 => to_unsigned(914, 10), 1858 => to_unsigned(832, 10), 1859 => to_unsigned(61, 10), 1860 => to_unsigned(250, 10), 1861 => to_unsigned(299, 10), 1862 => to_unsigned(143, 10), 1863 => to_unsigned(746, 10), 1864 => to_unsigned(474, 10), 1865 => to_unsigned(692, 10), 1866 => to_unsigned(230, 10), 1867 => to_unsigned(392, 10), 1868 => to_unsigned(274, 10), 1869 => to_unsigned(1004, 10), 1870 => to_unsigned(594, 10), 1871 => to_unsigned(334, 10), 1872 => to_unsigned(204, 10), 1873 => to_unsigned(92, 10), 1874 => to_unsigned(425, 10), 1875 => to_unsigned(720, 10), 1876 => to_unsigned(182, 10), 1877 => to_unsigned(254, 10), 1878 => to_unsigned(613, 10), 1879 => to_unsigned(226, 10), 1880 => to_unsigned(507, 10), 1881 => to_unsigned(685, 10), 1882 => to_unsigned(695, 10), 1883 => to_unsigned(347, 10), 1884 => to_unsigned(408, 10), 1885 => to_unsigned(320, 10), 1886 => to_unsigned(758, 10), 1887 => to_unsigned(9, 10), 1888 => to_unsigned(588, 10), 1889 => to_unsigned(354, 10), 1890 => to_unsigned(853, 10), 1891 => to_unsigned(14, 10), 1892 => to_unsigned(900, 10), 1893 => to_unsigned(393, 10), 1894 => to_unsigned(405, 10), 1895 => to_unsigned(659, 10), 1896 => to_unsigned(855, 10), 1897 => to_unsigned(283, 10), 1898 => to_unsigned(638, 10), 1899 => to_unsigned(1011, 10), 1900 => to_unsigned(593, 10), 1901 => to_unsigned(138, 10), 1902 => to_unsigned(798, 10), 1903 => to_unsigned(427, 10), 1904 => to_unsigned(928, 10), 1905 => to_unsigned(263, 10), 1906 => to_unsigned(36, 10), 1907 => to_unsigned(368, 10), 1908 => to_unsigned(443, 10), 1909 => to_unsigned(183, 10), 1910 => to_unsigned(590, 10), 1911 => to_unsigned(998, 10), 1912 => to_unsigned(640, 10), 1913 => to_unsigned(387, 10), 1914 => to_unsigned(475, 10), 1915 => to_unsigned(683, 10), 1916 => to_unsigned(26, 10), 1917 => to_unsigned(797, 10), 1918 => to_unsigned(839, 10), 1919 => to_unsigned(190, 10), 1920 => to_unsigned(856, 10), 1921 => to_unsigned(560, 10), 1922 => to_unsigned(853, 10), 1923 => to_unsigned(928, 10), 1924 => to_unsigned(903, 10), 1925 => to_unsigned(478, 10), 1926 => to_unsigned(199, 10), 1927 => to_unsigned(837, 10), 1928 => to_unsigned(464, 10), 1929 => to_unsigned(520, 10), 1930 => to_unsigned(952, 10), 1931 => to_unsigned(1021, 10), 1932 => to_unsigned(231, 10), 1933 => to_unsigned(472, 10), 1934 => to_unsigned(443, 10), 1935 => to_unsigned(75, 10), 1936 => to_unsigned(122, 10), 1937 => to_unsigned(982, 10), 1938 => to_unsigned(802, 10), 1939 => to_unsigned(312, 10), 1940 => to_unsigned(873, 10), 1941 => to_unsigned(675, 10), 1942 => to_unsigned(614, 10), 1943 => to_unsigned(426, 10), 1944 => to_unsigned(229, 10), 1945 => to_unsigned(901, 10), 1946 => to_unsigned(47, 10), 1947 => to_unsigned(986, 10), 1948 => to_unsigned(690, 10), 1949 => to_unsigned(749, 10), 1950 => to_unsigned(131, 10), 1951 => to_unsigned(409, 10), 1952 => to_unsigned(747, 10), 1953 => to_unsigned(193, 10), 1954 => to_unsigned(934, 10), 1955 => to_unsigned(242, 10), 1956 => to_unsigned(939, 10), 1957 => to_unsigned(599, 10), 1958 => to_unsigned(150, 10), 1959 => to_unsigned(621, 10), 1960 => to_unsigned(669, 10), 1961 => to_unsigned(291, 10), 1962 => to_unsigned(259, 10), 1963 => to_unsigned(979, 10), 1964 => to_unsigned(615, 10), 1965 => to_unsigned(701, 10), 1966 => to_unsigned(450, 10), 1967 => to_unsigned(276, 10), 1968 => to_unsigned(19, 10), 1969 => to_unsigned(1008, 10), 1970 => to_unsigned(837, 10), 1971 => to_unsigned(816, 10), 1972 => to_unsigned(892, 10), 1973 => to_unsigned(517, 10), 1974 => to_unsigned(559, 10), 1975 => to_unsigned(210, 10), 1976 => to_unsigned(420, 10), 1977 => to_unsigned(475, 10), 1978 => to_unsigned(74, 10), 1979 => to_unsigned(321, 10), 1980 => to_unsigned(639, 10), 1981 => to_unsigned(806, 10), 1982 => to_unsigned(129, 10), 1983 => to_unsigned(715, 10), 1984 => to_unsigned(687, 10), 1985 => to_unsigned(438, 10), 1986 => to_unsigned(79, 10), 1987 => to_unsigned(179, 10), 1988 => to_unsigned(41, 10), 1989 => to_unsigned(395, 10), 1990 => to_unsigned(775, 10), 1991 => to_unsigned(959, 10), 1992 => to_unsigned(123, 10), 1993 => to_unsigned(995, 10), 1994 => to_unsigned(918, 10), 1995 => to_unsigned(509, 10), 1996 => to_unsigned(294, 10), 1997 => to_unsigned(142, 10), 1998 => to_unsigned(718, 10), 1999 => to_unsigned(976, 10), 2000 => to_unsigned(495, 10), 2001 => to_unsigned(544, 10), 2002 => to_unsigned(361, 10), 2003 => to_unsigned(886, 10), 2004 => to_unsigned(489, 10), 2005 => to_unsigned(362, 10), 2006 => to_unsigned(651, 10), 2007 => to_unsigned(625, 10), 2008 => to_unsigned(1015, 10), 2009 => to_unsigned(801, 10), 2010 => to_unsigned(923, 10), 2011 => to_unsigned(228, 10), 2012 => to_unsigned(886, 10), 2013 => to_unsigned(734, 10), 2014 => to_unsigned(52, 10), 2015 => to_unsigned(97, 10), 2016 => to_unsigned(447, 10), 2017 => to_unsigned(918, 10), 2018 => to_unsigned(374, 10), 2019 => to_unsigned(640, 10), 2020 => to_unsigned(416, 10), 2021 => to_unsigned(160, 10), 2022 => to_unsigned(543, 10), 2023 => to_unsigned(191, 10), 2024 => to_unsigned(533, 10), 2025 => to_unsigned(738, 10), 2026 => to_unsigned(486, 10), 2027 => to_unsigned(441, 10), 2028 => to_unsigned(523, 10), 2029 => to_unsigned(988, 10), 2030 => to_unsigned(626, 10), 2031 => to_unsigned(725, 10), 2032 => to_unsigned(46, 10), 2033 => to_unsigned(166, 10), 2034 => to_unsigned(790, 10), 2035 => to_unsigned(399, 10), 2036 => to_unsigned(730, 10), 2037 => to_unsigned(811, 10), 2038 => to_unsigned(254, 10), 2039 => to_unsigned(164, 10), 2040 => to_unsigned(60, 10), 2041 => to_unsigned(372, 10), 2042 => to_unsigned(453, 10), 2043 => to_unsigned(677, 10), 2044 => to_unsigned(579, 10), 2045 => to_unsigned(470, 10), 2046 => to_unsigned(610, 10), 2047 => to_unsigned(439, 10))
        )
    );
    constant averages : averages_t := (
        0 => (0 => to_unsigned(681, 10), 1 => to_unsigned(572, 10), 2 => to_unsigned(579, 10), 3 => to_unsigned(297, 10), 4 => to_unsigned(367, 10), 5 => to_unsigned(327, 10), 6 => to_unsigned(554, 10), 7 => to_unsigned(510, 10), 8 => to_unsigned(470, 10), 9 => to_unsigned(532, 10), 10 => to_unsigned(358, 10), 11 => to_unsigned(724, 10), 12 => to_unsigned(507, 10), 13 => to_unsigned(508, 10), 14 => to_unsigned(314, 10), 15 => to_unsigned(489, 10), 16 => to_unsigned(377, 10), 17 => to_unsigned(601, 10), 18 => to_unsigned(547, 10), 19 => to_unsigned(419, 10), 20 => to_unsigned(532, 10), 21 => to_unsigned(538, 10), 22 => to_unsigned(418, 10), 23 => to_unsigned(505, 10), 24 => to_unsigned(511, 10), 25 => to_unsigned(590, 10), 26 => to_unsigned(680, 10), 27 => to_unsigned(499, 10), 28 => to_unsigned(480, 10), 29 => to_unsigned(443, 10), 30 => to_unsigned(593, 10), 31 => to_unsigned(544, 10), 32 => to_unsigned(423, 10), 33 => to_unsigned(693, 10), 34 => to_unsigned(550, 10), 35 => to_unsigned(469, 10), 36 => to_unsigned(449, 10), 37 => to_unsigned(462, 10), 38 => to_unsigned(375, 10), 39 => to_unsigned(593, 10), 40 => to_unsigned(452, 10), 41 => to_unsigned(515, 10), 42 => to_unsigned(499, 10), 43 => to_unsigned(229, 10), 44 => to_unsigned(447, 10), 45 => to_unsigned(468, 10), 46 => to_unsigned(622, 10), 47 => to_unsigned(483, 10), 48 => to_unsigned(503, 10), 49 => to_unsigned(553, 10), 50 => to_unsigned(461, 10), 51 => to_unsigned(618, 10), 52 => to_unsigned(591, 10), 53 => to_unsigned(508, 10), 54 => to_unsigned(459, 10), 55 => to_unsigned(521, 10), 56 => to_unsigned(373, 10), 57 => to_unsigned(517, 10), 58 => to_unsigned(401, 10), 59 => to_unsigned(472, 10), 60 => to_unsigned(637, 10), 61 => to_unsigned(537, 10), 62 => to_unsigned(333, 10), 63 => to_unsigned(507, 10), 64 => to_unsigned(440, 10), 65 => to_unsigned(422, 10), 66 => to_unsigned(487, 10), 67 => to_unsigned(551, 10), 68 => to_unsigned(555, 10), 69 => to_unsigned(497, 10), 70 => to_unsigned(525, 10), 71 => to_unsigned(525, 10), 72 => to_unsigned(387, 10), 73 => to_unsigned(571, 10), 74 => to_unsigned(618, 10), 75 => to_unsigned(530, 10), 76 => to_unsigned(570, 10), 77 => to_unsigned(417, 10), 78 => to_unsigned(483, 10), 79 => to_unsigned(694, 10), 80 => to_unsigned(467, 10), 81 => to_unsigned(557, 10), 82 => to_unsigned(574, 10), 83 => to_unsigned(412, 10), 84 => to_unsigned(455, 10), 85 => to_unsigned(565, 10), 86 => to_unsigned(555, 10), 87 => to_unsigned(505, 10), 88 => to_unsigned(430, 10), 89 => to_unsigned(477, 10), 90 => to_unsigned(462, 10), 91 => to_unsigned(623, 10), 92 => to_unsigned(399, 10), 93 => to_unsigned(393, 10), 94 => to_unsigned(401, 10), 95 => to_unsigned(597, 10), 96 => to_unsigned(614, 10), 97 => to_unsigned(419, 10), 98 => to_unsigned(467, 10), 99 => to_unsigned(637, 10), 100 => to_unsigned(662, 10), 101 => to_unsigned(470, 10), 102 => to_unsigned(556, 10), 103 => to_unsigned(324, 10), 104 => to_unsigned(639, 10), 105 => to_unsigned(561, 10), 106 => to_unsigned(541, 10), 107 => to_unsigned(488, 10), 108 => to_unsigned(532, 10), 109 => to_unsigned(478, 10), 110 => to_unsigned(496, 10), 111 => to_unsigned(541, 10), 112 => to_unsigned(626, 10), 113 => to_unsigned(384, 10), 114 => to_unsigned(595, 10), 115 => to_unsigned(565, 10), 116 => to_unsigned(478, 10), 117 => to_unsigned(399, 10), 118 => to_unsigned(482, 10), 119 => to_unsigned(605, 10), 120 => to_unsigned(565, 10), 121 => to_unsigned(580, 10), 122 => to_unsigned(514, 10), 123 => to_unsigned(252, 10), 124 => to_unsigned(437, 10), 125 => to_unsigned(595, 10), 126 => to_unsigned(452, 10), 127 => to_unsigned(584, 10), 128 => to_unsigned(411, 10), 129 => to_unsigned(401, 10), 130 => to_unsigned(592, 10), 131 => to_unsigned(581, 10), 132 => to_unsigned(404, 10), 133 => to_unsigned(629, 10), 134 => to_unsigned(561, 10), 135 => to_unsigned(628, 10), 136 => to_unsigned(618, 10), 137 => to_unsigned(479, 10), 138 => to_unsigned(614, 10), 139 => to_unsigned(584, 10), 140 => to_unsigned(502, 10), 141 => to_unsigned(382, 10), 142 => to_unsigned(526, 10), 143 => to_unsigned(531, 10), 144 => to_unsigned(590, 10), 145 => to_unsigned(500, 10), 146 => to_unsigned(445, 10), 147 => to_unsigned(570, 10), 148 => to_unsigned(483, 10), 149 => to_unsigned(582, 10), 150 => to_unsigned(415, 10), 151 => to_unsigned(488, 10), 152 => to_unsigned(501, 10), 153 => to_unsigned(632, 10), 154 => to_unsigned(713, 10), 155 => to_unsigned(335, 10), 156 => to_unsigned(422, 10), 157 => to_unsigned(507, 10), 158 => to_unsigned(379, 10), 159 => to_unsigned(473, 10), 160 => to_unsigned(434, 10), 161 => to_unsigned(566, 10), 162 => to_unsigned(550, 10), 163 => to_unsigned(306, 10), 164 => to_unsigned(597, 10), 165 => to_unsigned(402, 10), 166 => to_unsigned(538, 10), 167 => to_unsigned(632, 10), 168 => to_unsigned(483, 10), 169 => to_unsigned(384, 10), 170 => to_unsigned(486, 10), 171 => to_unsigned(580, 10), 172 => to_unsigned(597, 10), 173 => to_unsigned(477, 10), 174 => to_unsigned(548, 10), 175 => to_unsigned(369, 10), 176 => to_unsigned(514, 10), 177 => to_unsigned(473, 10), 178 => to_unsigned(602, 10), 179 => to_unsigned(567, 10), 180 => to_unsigned(226, 10), 181 => to_unsigned(563, 10), 182 => to_unsigned(470, 10), 183 => to_unsigned(690, 10), 184 => to_unsigned(581, 10), 185 => to_unsigned(416, 10), 186 => to_unsigned(440, 10), 187 => to_unsigned(402, 10), 188 => to_unsigned(303, 10), 189 => to_unsigned(609, 10), 190 => to_unsigned(419, 10), 191 => to_unsigned(541, 10), 192 => to_unsigned(483, 10), 193 => to_unsigned(322, 10), 194 => to_unsigned(426, 10), 195 => to_unsigned(690, 10), 196 => to_unsigned(378, 10), 197 => to_unsigned(529, 10), 198 => to_unsigned(474, 10), 199 => to_unsigned(510, 10), 200 => to_unsigned(616, 10), 201 => to_unsigned(546, 10), 202 => to_unsigned(546, 10), 203 => to_unsigned(407, 10), 204 => to_unsigned(509, 10), 205 => to_unsigned(502, 10), 206 => to_unsigned(466, 10), 207 => to_unsigned(640, 10), 208 => to_unsigned(457, 10), 209 => to_unsigned(403, 10), 210 => to_unsigned(295, 10), 211 => to_unsigned(573, 10), 212 => to_unsigned(666, 10), 213 => to_unsigned(543, 10), 214 => to_unsigned(379, 10), 215 => to_unsigned(510, 10), 216 => to_unsigned(411, 10), 217 => to_unsigned(540, 10), 218 => to_unsigned(632, 10), 219 => to_unsigned(691, 10), 220 => to_unsigned(690, 10), 221 => to_unsigned(564, 10), 222 => to_unsigned(427, 10), 223 => to_unsigned(766, 10), 224 => to_unsigned(550, 10), 225 => to_unsigned(481, 10), 226 => to_unsigned(476, 10), 227 => to_unsigned(571, 10), 228 => to_unsigned(326, 10), 229 => to_unsigned(569, 10), 230 => to_unsigned(562, 10), 231 => to_unsigned(502, 10), 232 => to_unsigned(494, 10), 233 => to_unsigned(403, 10), 234 => to_unsigned(358, 10), 235 => to_unsigned(758, 10), 236 => to_unsigned(496, 10), 237 => to_unsigned(579, 10), 238 => to_unsigned(538, 10), 239 => to_unsigned(567, 10), 240 => to_unsigned(685, 10), 241 => to_unsigned(522, 10), 242 => to_unsigned(648, 10), 243 => to_unsigned(515, 10), 244 => to_unsigned(522, 10), 245 => to_unsigned(496, 10), 246 => to_unsigned(591, 10), 247 => to_unsigned(442, 10), 248 => to_unsigned(537, 10), 249 => to_unsigned(596, 10), 250 => to_unsigned(541, 10), 251 => to_unsigned(409, 10), 252 => to_unsigned(509, 10), 253 => to_unsigned(449, 10), 254 => to_unsigned(563, 10), 255 => to_unsigned(509, 10), 256 => to_unsigned(494, 10), 257 => to_unsigned(685, 10), 258 => to_unsigned(556, 10), 259 => to_unsigned(419, 10), 260 => to_unsigned(551, 10), 261 => to_unsigned(421, 10), 262 => to_unsigned(557, 10), 263 => to_unsigned(584, 10), 264 => to_unsigned(503, 10), 265 => to_unsigned(503, 10), 266 => to_unsigned(524, 10), 267 => to_unsigned(448, 10), 268 => to_unsigned(335, 10), 269 => to_unsigned(577, 10), 270 => to_unsigned(593, 10), 271 => to_unsigned(555, 10), 272 => to_unsigned(468, 10), 273 => to_unsigned(571, 10), 274 => to_unsigned(477, 10), 275 => to_unsigned(405, 10), 276 => to_unsigned(652, 10), 277 => to_unsigned(484, 10), 278 => to_unsigned(381, 10), 279 => to_unsigned(503, 10), 280 => to_unsigned(715, 10), 281 => to_unsigned(537, 10), 282 => to_unsigned(608, 10), 283 => to_unsigned(609, 10), 284 => to_unsigned(561, 10), 285 => to_unsigned(460, 10), 286 => to_unsigned(468, 10), 287 => to_unsigned(483, 10), 288 => to_unsigned(536, 10), 289 => to_unsigned(437, 10), 290 => to_unsigned(488, 10), 291 => to_unsigned(480, 10), 292 => to_unsigned(521, 10), 293 => to_unsigned(383, 10), 294 => to_unsigned(611, 10), 295 => to_unsigned(587, 10), 296 => to_unsigned(487, 10), 297 => to_unsigned(506, 10), 298 => to_unsigned(441, 10), 299 => to_unsigned(590, 10), 300 => to_unsigned(327, 10), 301 => to_unsigned(469, 10), 302 => to_unsigned(498, 10), 303 => to_unsigned(411, 10), 304 => to_unsigned(708, 10), 305 => to_unsigned(430, 10), 306 => to_unsigned(770, 10), 307 => to_unsigned(472, 10), 308 => to_unsigned(408, 10), 309 => to_unsigned(504, 10), 310 => to_unsigned(345, 10), 311 => to_unsigned(575, 10), 312 => to_unsigned(532, 10), 313 => to_unsigned(502, 10), 314 => to_unsigned(463, 10), 315 => to_unsigned(672, 10), 316 => to_unsigned(524, 10), 317 => to_unsigned(542, 10), 318 => to_unsigned(512, 10), 319 => to_unsigned(446, 10), 320 => to_unsigned(461, 10), 321 => to_unsigned(461, 10), 322 => to_unsigned(380, 10), 323 => to_unsigned(429, 10), 324 => to_unsigned(537, 10), 325 => to_unsigned(574, 10), 326 => to_unsigned(534, 10), 327 => to_unsigned(514, 10), 328 => to_unsigned(630, 10), 329 => to_unsigned(588, 10), 330 => to_unsigned(425, 10), 331 => to_unsigned(498, 10), 332 => to_unsigned(588, 10), 333 => to_unsigned(547, 10), 334 => to_unsigned(431, 10), 335 => to_unsigned(465, 10), 336 => to_unsigned(329, 10), 337 => to_unsigned(660, 10), 338 => to_unsigned(534, 10), 339 => to_unsigned(597, 10), 340 => to_unsigned(513, 10), 341 => to_unsigned(672, 10), 342 => to_unsigned(515, 10), 343 => to_unsigned(566, 10), 344 => to_unsigned(390, 10), 345 => to_unsigned(636, 10), 346 => to_unsigned(339, 10), 347 => to_unsigned(596, 10), 348 => to_unsigned(556, 10), 349 => to_unsigned(387, 10), 350 => to_unsigned(308, 10), 351 => to_unsigned(549, 10), 352 => to_unsigned(558, 10), 353 => to_unsigned(385, 10), 354 => to_unsigned(401, 10), 355 => to_unsigned(406, 10), 356 => to_unsigned(402, 10), 357 => to_unsigned(479, 10), 358 => to_unsigned(417, 10), 359 => to_unsigned(497, 10), 360 => to_unsigned(372, 10), 361 => to_unsigned(453, 10), 362 => to_unsigned(638, 10), 363 => to_unsigned(386, 10), 364 => to_unsigned(543, 10), 365 => to_unsigned(708, 10), 366 => to_unsigned(564, 10), 367 => to_unsigned(355, 10), 368 => to_unsigned(630, 10), 369 => to_unsigned(405, 10), 370 => to_unsigned(657, 10), 371 => to_unsigned(471, 10), 372 => to_unsigned(515, 10), 373 => to_unsigned(484, 10), 374 => to_unsigned(503, 10), 375 => to_unsigned(583, 10), 376 => to_unsigned(646, 10), 377 => to_unsigned(391, 10), 378 => to_unsigned(589, 10), 379 => to_unsigned(524, 10), 380 => to_unsigned(568, 10), 381 => to_unsigned(462, 10), 382 => to_unsigned(740, 10), 383 => to_unsigned(548, 10), 384 => to_unsigned(435, 10), 385 => to_unsigned(336, 10), 386 => to_unsigned(507, 10), 387 => to_unsigned(491, 10), 388 => to_unsigned(630, 10), 389 => to_unsigned(610, 10), 390 => to_unsigned(584, 10), 391 => to_unsigned(585, 10), 392 => to_unsigned(590, 10), 393 => to_unsigned(625, 10), 394 => to_unsigned(561, 10), 395 => to_unsigned(482, 10), 396 => to_unsigned(560, 10), 397 => to_unsigned(549, 10), 398 => to_unsigned(432, 10), 399 => to_unsigned(506, 10), 400 => to_unsigned(473, 10), 401 => to_unsigned(795, 10), 402 => to_unsigned(362, 10), 403 => to_unsigned(354, 10), 404 => to_unsigned(454, 10), 405 => to_unsigned(447, 10), 406 => to_unsigned(379, 10), 407 => to_unsigned(600, 10), 408 => to_unsigned(320, 10), 409 => to_unsigned(507, 10), 410 => to_unsigned(418, 10), 411 => to_unsigned(613, 10), 412 => to_unsigned(711, 10), 413 => to_unsigned(620, 10), 414 => to_unsigned(337, 10), 415 => to_unsigned(670, 10), 416 => to_unsigned(388, 10), 417 => to_unsigned(508, 10), 418 => to_unsigned(626, 10), 419 => to_unsigned(490, 10), 420 => to_unsigned(438, 10), 421 => to_unsigned(502, 10), 422 => to_unsigned(609, 10), 423 => to_unsigned(550, 10), 424 => to_unsigned(427, 10), 425 => to_unsigned(316, 10), 426 => to_unsigned(338, 10), 427 => to_unsigned(637, 10), 428 => to_unsigned(463, 10), 429 => to_unsigned(557, 10), 430 => to_unsigned(411, 10), 431 => to_unsigned(434, 10), 432 => to_unsigned(410, 10), 433 => to_unsigned(408, 10), 434 => to_unsigned(601, 10), 435 => to_unsigned(537, 10), 436 => to_unsigned(526, 10), 437 => to_unsigned(601, 10), 438 => to_unsigned(572, 10), 439 => to_unsigned(490, 10), 440 => to_unsigned(393, 10), 441 => to_unsigned(419, 10), 442 => to_unsigned(533, 10), 443 => to_unsigned(487, 10), 444 => to_unsigned(422, 10), 445 => to_unsigned(515, 10), 446 => to_unsigned(355, 10), 447 => to_unsigned(439, 10), 448 => to_unsigned(546, 10), 449 => to_unsigned(584, 10), 450 => to_unsigned(690, 10), 451 => to_unsigned(635, 10), 452 => to_unsigned(593, 10), 453 => to_unsigned(435, 10), 454 => to_unsigned(476, 10), 455 => to_unsigned(593, 10), 456 => to_unsigned(554, 10), 457 => to_unsigned(483, 10), 458 => to_unsigned(437, 10), 459 => to_unsigned(472, 10), 460 => to_unsigned(398, 10), 461 => to_unsigned(532, 10), 462 => to_unsigned(382, 10), 463 => to_unsigned(386, 10), 464 => to_unsigned(467, 10), 465 => to_unsigned(407, 10), 466 => to_unsigned(478, 10), 467 => to_unsigned(647, 10), 468 => to_unsigned(576, 10), 469 => to_unsigned(534, 10), 470 => to_unsigned(554, 10), 471 => to_unsigned(358, 10), 472 => to_unsigned(548, 10), 473 => to_unsigned(506, 10), 474 => to_unsigned(740, 10), 475 => to_unsigned(529, 10), 476 => to_unsigned(582, 10), 477 => to_unsigned(490, 10), 478 => to_unsigned(536, 10), 479 => to_unsigned(521, 10), 480 => to_unsigned(315, 10), 481 => to_unsigned(626, 10), 482 => to_unsigned(495, 10), 483 => to_unsigned(437, 10), 484 => to_unsigned(446, 10), 485 => to_unsigned(692, 10), 486 => to_unsigned(618, 10), 487 => to_unsigned(343, 10), 488 => to_unsigned(531, 10), 489 => to_unsigned(327, 10), 490 => to_unsigned(517, 10), 491 => to_unsigned(424, 10), 492 => to_unsigned(496, 10), 493 => to_unsigned(481, 10), 494 => to_unsigned(477, 10), 495 => to_unsigned(538, 10), 496 => to_unsigned(511, 10), 497 => to_unsigned(519, 10), 498 => to_unsigned(383, 10), 499 => to_unsigned(496, 10), 500 => to_unsigned(568, 10), 501 => to_unsigned(723, 10), 502 => to_unsigned(529, 10), 503 => to_unsigned(567, 10), 504 => to_unsigned(593, 10), 505 => to_unsigned(756, 10), 506 => to_unsigned(510, 10), 507 => to_unsigned(628, 10), 508 => to_unsigned(520, 10), 509 => to_unsigned(520, 10), 510 => to_unsigned(412, 10), 511 => to_unsigned(393, 10), 512 => to_unsigned(592, 10), 513 => to_unsigned(554, 10), 514 => to_unsigned(420, 10), 515 => to_unsigned(600, 10), 516 => to_unsigned(411, 10), 517 => to_unsigned(475, 10), 518 => to_unsigned(643, 10), 519 => to_unsigned(519, 10), 520 => to_unsigned(281, 10), 521 => to_unsigned(457, 10), 522 => to_unsigned(544, 10), 523 => to_unsigned(502, 10), 524 => to_unsigned(475, 10), 525 => to_unsigned(533, 10), 526 => to_unsigned(572, 10), 527 => to_unsigned(607, 10), 528 => to_unsigned(408, 10), 529 => to_unsigned(456, 10), 530 => to_unsigned(437, 10), 531 => to_unsigned(540, 10), 532 => to_unsigned(749, 10), 533 => to_unsigned(419, 10), 534 => to_unsigned(479, 10), 535 => to_unsigned(786, 10), 536 => to_unsigned(368, 10), 537 => to_unsigned(504, 10), 538 => to_unsigned(589, 10), 539 => to_unsigned(547, 10), 540 => to_unsigned(515, 10), 541 => to_unsigned(456, 10), 542 => to_unsigned(573, 10), 543 => to_unsigned(447, 10), 544 => to_unsigned(595, 10), 545 => to_unsigned(460, 10), 546 => to_unsigned(462, 10), 547 => to_unsigned(269, 10), 548 => to_unsigned(449, 10), 549 => to_unsigned(587, 10), 550 => to_unsigned(462, 10), 551 => to_unsigned(402, 10), 552 => to_unsigned(515, 10), 553 => to_unsigned(408, 10), 554 => to_unsigned(603, 10), 555 => to_unsigned(595, 10), 556 => to_unsigned(544, 10), 557 => to_unsigned(576, 10), 558 => to_unsigned(537, 10), 559 => to_unsigned(645, 10), 560 => to_unsigned(411, 10), 561 => to_unsigned(502, 10), 562 => to_unsigned(452, 10), 563 => to_unsigned(657, 10), 564 => to_unsigned(403, 10), 565 => to_unsigned(439, 10), 566 => to_unsigned(498, 10), 567 => to_unsigned(450, 10), 568 => to_unsigned(524, 10), 569 => to_unsigned(471, 10), 570 => to_unsigned(411, 10), 571 => to_unsigned(532, 10), 572 => to_unsigned(546, 10), 573 => to_unsigned(446, 10), 574 => to_unsigned(427, 10), 575 => to_unsigned(486, 10), 576 => to_unsigned(479, 10), 577 => to_unsigned(535, 10), 578 => to_unsigned(328, 10), 579 => to_unsigned(350, 10), 580 => to_unsigned(550, 10), 581 => to_unsigned(466, 10), 582 => to_unsigned(354, 10), 583 => to_unsigned(662, 10), 584 => to_unsigned(539, 10), 585 => to_unsigned(524, 10), 586 => to_unsigned(676, 10), 587 => to_unsigned(629, 10), 588 => to_unsigned(447, 10), 589 => to_unsigned(462, 10), 590 => to_unsigned(634, 10), 591 => to_unsigned(567, 10), 592 => to_unsigned(442, 10), 593 => to_unsigned(623, 10), 594 => to_unsigned(463, 10), 595 => to_unsigned(519, 10), 596 => to_unsigned(361, 10), 597 => to_unsigned(570, 10), 598 => to_unsigned(449, 10), 599 => to_unsigned(316, 10), 600 => to_unsigned(576, 10), 601 => to_unsigned(665, 10), 602 => to_unsigned(595, 10), 603 => to_unsigned(379, 10), 604 => to_unsigned(585, 10), 605 => to_unsigned(529, 10), 606 => to_unsigned(609, 10), 607 => to_unsigned(607, 10), 608 => to_unsigned(555, 10), 609 => to_unsigned(616, 10), 610 => to_unsigned(621, 10), 611 => to_unsigned(416, 10), 612 => to_unsigned(427, 10), 613 => to_unsigned(502, 10), 614 => to_unsigned(436, 10), 615 => to_unsigned(514, 10), 616 => to_unsigned(510, 10), 617 => to_unsigned(685, 10), 618 => to_unsigned(465, 10), 619 => to_unsigned(429, 10), 620 => to_unsigned(523, 10), 621 => to_unsigned(524, 10), 622 => to_unsigned(703, 10), 623 => to_unsigned(606, 10), 624 => to_unsigned(602, 10), 625 => to_unsigned(654, 10), 626 => to_unsigned(653, 10), 627 => to_unsigned(501, 10), 628 => to_unsigned(583, 10), 629 => to_unsigned(420, 10), 630 => to_unsigned(439, 10), 631 => to_unsigned(524, 10), 632 => to_unsigned(518, 10), 633 => to_unsigned(525, 10), 634 => to_unsigned(511, 10), 635 => to_unsigned(410, 10), 636 => to_unsigned(479, 10), 637 => to_unsigned(449, 10), 638 => to_unsigned(405, 10), 639 => to_unsigned(453, 10), 640 => to_unsigned(507, 10), 641 => to_unsigned(523, 10), 642 => to_unsigned(619, 10), 643 => to_unsigned(445, 10), 644 => to_unsigned(484, 10), 645 => to_unsigned(542, 10), 646 => to_unsigned(592, 10), 647 => to_unsigned(645, 10), 648 => to_unsigned(502, 10), 649 => to_unsigned(420, 10), 650 => to_unsigned(515, 10), 651 => to_unsigned(566, 10), 652 => to_unsigned(551, 10), 653 => to_unsigned(533, 10), 654 => to_unsigned(652, 10), 655 => to_unsigned(358, 10), 656 => to_unsigned(366, 10), 657 => to_unsigned(549, 10), 658 => to_unsigned(481, 10), 659 => to_unsigned(594, 10), 660 => to_unsigned(449, 10), 661 => to_unsigned(439, 10), 662 => to_unsigned(587, 10), 663 => to_unsigned(448, 10), 664 => to_unsigned(609, 10), 665 => to_unsigned(453, 10), 666 => to_unsigned(526, 10), 667 => to_unsigned(507, 10), 668 => to_unsigned(579, 10), 669 => to_unsigned(362, 10), 670 => to_unsigned(609, 10), 671 => to_unsigned(722, 10), 672 => to_unsigned(355, 10), 673 => to_unsigned(593, 10), 674 => to_unsigned(442, 10), 675 => to_unsigned(506, 10), 676 => to_unsigned(350, 10), 677 => to_unsigned(555, 10), 678 => to_unsigned(300, 10), 679 => to_unsigned(385, 10), 680 => to_unsigned(380, 10), 681 => to_unsigned(441, 10), 682 => to_unsigned(516, 10), 683 => to_unsigned(506, 10), 684 => to_unsigned(489, 10), 685 => to_unsigned(547, 10), 686 => to_unsigned(480, 10), 687 => to_unsigned(416, 10), 688 => to_unsigned(336, 10), 689 => to_unsigned(526, 10), 690 => to_unsigned(454, 10), 691 => to_unsigned(510, 10), 692 => to_unsigned(418, 10), 693 => to_unsigned(510, 10), 694 => to_unsigned(471, 10), 695 => to_unsigned(383, 10), 696 => to_unsigned(448, 10), 697 => to_unsigned(461, 10), 698 => to_unsigned(556, 10), 699 => to_unsigned(315, 10), 700 => to_unsigned(540, 10), 701 => to_unsigned(420, 10), 702 => to_unsigned(631, 10), 703 => to_unsigned(476, 10), 704 => to_unsigned(706, 10), 705 => to_unsigned(488, 10), 706 => to_unsigned(563, 10), 707 => to_unsigned(425, 10), 708 => to_unsigned(576, 10), 709 => to_unsigned(439, 10), 710 => to_unsigned(359, 10), 711 => to_unsigned(512, 10), 712 => to_unsigned(460, 10), 713 => to_unsigned(584, 10), 714 => to_unsigned(290, 10), 715 => to_unsigned(539, 10), 716 => to_unsigned(491, 10), 717 => to_unsigned(541, 10), 718 => to_unsigned(539, 10), 719 => to_unsigned(579, 10), 720 => to_unsigned(450, 10), 721 => to_unsigned(486, 10), 722 => to_unsigned(569, 10), 723 => to_unsigned(544, 10), 724 => to_unsigned(560, 10), 725 => to_unsigned(604, 10), 726 => to_unsigned(449, 10), 727 => to_unsigned(610, 10), 728 => to_unsigned(510, 10), 729 => to_unsigned(469, 10), 730 => to_unsigned(361, 10), 731 => to_unsigned(526, 10), 732 => to_unsigned(460, 10), 733 => to_unsigned(725, 10), 734 => to_unsigned(577, 10), 735 => to_unsigned(588, 10), 736 => to_unsigned(572, 10), 737 => to_unsigned(505, 10), 738 => to_unsigned(503, 10), 739 => to_unsigned(574, 10), 740 => to_unsigned(484, 10), 741 => to_unsigned(275, 10), 742 => to_unsigned(619, 10), 743 => to_unsigned(649, 10), 744 => to_unsigned(595, 10), 745 => to_unsigned(532, 10), 746 => to_unsigned(432, 10), 747 => to_unsigned(477, 10), 748 => to_unsigned(580, 10), 749 => to_unsigned(547, 10), 750 => to_unsigned(632, 10), 751 => to_unsigned(682, 10), 752 => to_unsigned(557, 10), 753 => to_unsigned(600, 10), 754 => to_unsigned(497, 10), 755 => to_unsigned(489, 10), 756 => to_unsigned(460, 10), 757 => to_unsigned(498, 10), 758 => to_unsigned(489, 10), 759 => to_unsigned(521, 10), 760 => to_unsigned(511, 10), 761 => to_unsigned(586, 10), 762 => to_unsigned(391, 10), 763 => to_unsigned(431, 10), 764 => to_unsigned(506, 10), 765 => to_unsigned(674, 10), 766 => to_unsigned(639, 10), 767 => to_unsigned(553, 10), 768 => to_unsigned(566, 10), 769 => to_unsigned(476, 10), 770 => to_unsigned(635, 10), 771 => to_unsigned(319, 10), 772 => to_unsigned(612, 10), 773 => to_unsigned(436, 10), 774 => to_unsigned(624, 10), 775 => to_unsigned(354, 10), 776 => to_unsigned(533, 10), 777 => to_unsigned(547, 10), 778 => to_unsigned(566, 10), 779 => to_unsigned(586, 10), 780 => to_unsigned(404, 10), 781 => to_unsigned(480, 10), 782 => to_unsigned(580, 10), 783 => to_unsigned(423, 10), 784 => to_unsigned(562, 10), 785 => to_unsigned(684, 10), 786 => to_unsigned(446, 10), 787 => to_unsigned(442, 10), 788 => to_unsigned(503, 10), 789 => to_unsigned(652, 10), 790 => to_unsigned(531, 10), 791 => to_unsigned(458, 10), 792 => to_unsigned(620, 10), 793 => to_unsigned(708, 10), 794 => to_unsigned(376, 10), 795 => to_unsigned(578, 10), 796 => to_unsigned(662, 10), 797 => to_unsigned(385, 10), 798 => to_unsigned(604, 10), 799 => to_unsigned(478, 10), 800 => to_unsigned(508, 10), 801 => to_unsigned(572, 10), 802 => to_unsigned(499, 10), 803 => to_unsigned(548, 10), 804 => to_unsigned(410, 10), 805 => to_unsigned(450, 10), 806 => to_unsigned(474, 10), 807 => to_unsigned(524, 10), 808 => to_unsigned(542, 10), 809 => to_unsigned(428, 10), 810 => to_unsigned(430, 10), 811 => to_unsigned(510, 10), 812 => to_unsigned(535, 10), 813 => to_unsigned(497, 10), 814 => to_unsigned(567, 10), 815 => to_unsigned(546, 10), 816 => to_unsigned(493, 10), 817 => to_unsigned(519, 10), 818 => to_unsigned(571, 10), 819 => to_unsigned(601, 10), 820 => to_unsigned(473, 10), 821 => to_unsigned(671, 10), 822 => to_unsigned(523, 10), 823 => to_unsigned(411, 10), 824 => to_unsigned(499, 10), 825 => to_unsigned(702, 10), 826 => to_unsigned(526, 10), 827 => to_unsigned(478, 10), 828 => to_unsigned(485, 10), 829 => to_unsigned(565, 10), 830 => to_unsigned(662, 10), 831 => to_unsigned(530, 10), 832 => to_unsigned(549, 10), 833 => to_unsigned(469, 10), 834 => to_unsigned(686, 10), 835 => to_unsigned(411, 10), 836 => to_unsigned(408, 10), 837 => to_unsigned(539, 10), 838 => to_unsigned(416, 10), 839 => to_unsigned(510, 10), 840 => to_unsigned(417, 10), 841 => to_unsigned(355, 10), 842 => to_unsigned(522, 10), 843 => to_unsigned(600, 10), 844 => to_unsigned(433, 10), 845 => to_unsigned(706, 10), 846 => to_unsigned(438, 10), 847 => to_unsigned(533, 10), 848 => to_unsigned(651, 10), 849 => to_unsigned(400, 10), 850 => to_unsigned(697, 10), 851 => to_unsigned(347, 10), 852 => to_unsigned(502, 10), 853 => to_unsigned(377, 10), 854 => to_unsigned(492, 10), 855 => to_unsigned(490, 10), 856 => to_unsigned(530, 10), 857 => to_unsigned(553, 10), 858 => to_unsigned(810, 10), 859 => to_unsigned(615, 10), 860 => to_unsigned(651, 10), 861 => to_unsigned(629, 10), 862 => to_unsigned(488, 10), 863 => to_unsigned(436, 10), 864 => to_unsigned(587, 10), 865 => to_unsigned(408, 10), 866 => to_unsigned(470, 10), 867 => to_unsigned(678, 10), 868 => to_unsigned(403, 10), 869 => to_unsigned(495, 10), 870 => to_unsigned(332, 10), 871 => to_unsigned(542, 10), 872 => to_unsigned(496, 10), 873 => to_unsigned(372, 10), 874 => to_unsigned(523, 10), 875 => to_unsigned(442, 10), 876 => to_unsigned(355, 10), 877 => to_unsigned(366, 10), 878 => to_unsigned(530, 10), 879 => to_unsigned(343, 10), 880 => to_unsigned(491, 10), 881 => to_unsigned(692, 10), 882 => to_unsigned(454, 10), 883 => to_unsigned(521, 10), 884 => to_unsigned(519, 10), 885 => to_unsigned(582, 10), 886 => to_unsigned(454, 10), 887 => to_unsigned(432, 10), 888 => to_unsigned(415, 10), 889 => to_unsigned(559, 10), 890 => to_unsigned(306, 10), 891 => to_unsigned(503, 10), 892 => to_unsigned(506, 10), 893 => to_unsigned(542, 10), 894 => to_unsigned(543, 10), 895 => to_unsigned(587, 10), 896 => to_unsigned(440, 10), 897 => to_unsigned(535, 10), 898 => to_unsigned(446, 10), 899 => to_unsigned(449, 10), 900 => to_unsigned(291, 10), 901 => to_unsigned(599, 10), 902 => to_unsigned(271, 10), 903 => to_unsigned(593, 10), 904 => to_unsigned(518, 10), 905 => to_unsigned(430, 10), 906 => to_unsigned(387, 10), 907 => to_unsigned(743, 10), 908 => to_unsigned(481, 10), 909 => to_unsigned(482, 10), 910 => to_unsigned(408, 10), 911 => to_unsigned(563, 10), 912 => to_unsigned(555, 10), 913 => to_unsigned(464, 10), 914 => to_unsigned(375, 10), 915 => to_unsigned(560, 10), 916 => to_unsigned(515, 10), 917 => to_unsigned(634, 10), 918 => to_unsigned(531, 10), 919 => to_unsigned(561, 10), 920 => to_unsigned(505, 10), 921 => to_unsigned(456, 10), 922 => to_unsigned(631, 10), 923 => to_unsigned(433, 10), 924 => to_unsigned(643, 10), 925 => to_unsigned(535, 10), 926 => to_unsigned(467, 10), 927 => to_unsigned(474, 10), 928 => to_unsigned(532, 10), 929 => to_unsigned(539, 10), 930 => to_unsigned(320, 10), 931 => to_unsigned(511, 10), 932 => to_unsigned(410, 10), 933 => to_unsigned(629, 10), 934 => to_unsigned(469, 10), 935 => to_unsigned(469, 10), 936 => to_unsigned(584, 10), 937 => to_unsigned(568, 10), 938 => to_unsigned(550, 10), 939 => to_unsigned(392, 10), 940 => to_unsigned(488, 10), 941 => to_unsigned(545, 10), 942 => to_unsigned(346, 10), 943 => to_unsigned(408, 10), 944 => to_unsigned(646, 10), 945 => to_unsigned(718, 10), 946 => to_unsigned(553, 10), 947 => to_unsigned(685, 10), 948 => to_unsigned(639, 10), 949 => to_unsigned(522, 10), 950 => to_unsigned(490, 10), 951 => to_unsigned(432, 10), 952 => to_unsigned(431, 10), 953 => to_unsigned(424, 10), 954 => to_unsigned(404, 10), 955 => to_unsigned(462, 10), 956 => to_unsigned(426, 10), 957 => to_unsigned(336, 10), 958 => to_unsigned(579, 10), 959 => to_unsigned(429, 10), 960 => to_unsigned(536, 10), 961 => to_unsigned(597, 10), 962 => to_unsigned(481, 10), 963 => to_unsigned(518, 10), 964 => to_unsigned(559, 10), 965 => to_unsigned(424, 10), 966 => to_unsigned(479, 10), 967 => to_unsigned(389, 10), 968 => to_unsigned(263, 10), 969 => to_unsigned(620, 10), 970 => to_unsigned(476, 10), 971 => to_unsigned(543, 10), 972 => to_unsigned(574, 10), 973 => to_unsigned(368, 10), 974 => to_unsigned(526, 10), 975 => to_unsigned(572, 10), 976 => to_unsigned(540, 10), 977 => to_unsigned(647, 10), 978 => to_unsigned(430, 10), 979 => to_unsigned(482, 10), 980 => to_unsigned(524, 10), 981 => to_unsigned(608, 10), 982 => to_unsigned(632, 10), 983 => to_unsigned(493, 10), 984 => to_unsigned(478, 10), 985 => to_unsigned(528, 10), 986 => to_unsigned(477, 10), 987 => to_unsigned(520, 10), 988 => to_unsigned(490, 10), 989 => to_unsigned(504, 10), 990 => to_unsigned(480, 10), 991 => to_unsigned(441, 10), 992 => to_unsigned(534, 10), 993 => to_unsigned(580, 10), 994 => to_unsigned(582, 10), 995 => to_unsigned(429, 10), 996 => to_unsigned(485, 10), 997 => to_unsigned(612, 10), 998 => to_unsigned(553, 10), 999 => to_unsigned(715, 10), 1000 => to_unsigned(279, 10), 1001 => to_unsigned(361, 10), 1002 => to_unsigned(581, 10), 1003 => to_unsigned(560, 10), 1004 => to_unsigned(480, 10), 1005 => to_unsigned(585, 10), 1006 => to_unsigned(436, 10), 1007 => to_unsigned(487, 10), 1008 => to_unsigned(499, 10), 1009 => to_unsigned(463, 10), 1010 => to_unsigned(610, 10), 1011 => to_unsigned(403, 10), 1012 => to_unsigned(445, 10), 1013 => to_unsigned(514, 10), 1014 => to_unsigned(449, 10), 1015 => to_unsigned(495, 10), 1016 => to_unsigned(555, 10), 1017 => to_unsigned(544, 10), 1018 => to_unsigned(666, 10), 1019 => to_unsigned(687, 10), 1020 => to_unsigned(604, 10), 1021 => to_unsigned(462, 10), 1022 => to_unsigned(436, 10), 1023 => to_unsigned(496, 10), 1024 => to_unsigned(399, 10), 1025 => to_unsigned(510, 10), 1026 => to_unsigned(563, 10), 1027 => to_unsigned(454, 10), 1028 => to_unsigned(522, 10), 1029 => to_unsigned(634, 10), 1030 => to_unsigned(685, 10), 1031 => to_unsigned(436, 10), 1032 => to_unsigned(511, 10), 1033 => to_unsigned(413, 10), 1034 => to_unsigned(705, 10), 1035 => to_unsigned(566, 10), 1036 => to_unsigned(406, 10), 1037 => to_unsigned(390, 10), 1038 => to_unsigned(510, 10), 1039 => to_unsigned(507, 10), 1040 => to_unsigned(539, 10), 1041 => to_unsigned(607, 10), 1042 => to_unsigned(456, 10), 1043 => to_unsigned(414, 10), 1044 => to_unsigned(486, 10), 1045 => to_unsigned(361, 10), 1046 => to_unsigned(434, 10), 1047 => to_unsigned(319, 10), 1048 => to_unsigned(608, 10), 1049 => to_unsigned(546, 10), 1050 => to_unsigned(550, 10), 1051 => to_unsigned(339, 10), 1052 => to_unsigned(436, 10), 1053 => to_unsigned(548, 10), 1054 => to_unsigned(493, 10), 1055 => to_unsigned(417, 10), 1056 => to_unsigned(453, 10), 1057 => to_unsigned(604, 10), 1058 => to_unsigned(468, 10), 1059 => to_unsigned(555, 10), 1060 => to_unsigned(531, 10), 1061 => to_unsigned(526, 10), 1062 => to_unsigned(610, 10), 1063 => to_unsigned(470, 10), 1064 => to_unsigned(494, 10), 1065 => to_unsigned(532, 10), 1066 => to_unsigned(573, 10), 1067 => to_unsigned(466, 10), 1068 => to_unsigned(450, 10), 1069 => to_unsigned(310, 10), 1070 => to_unsigned(554, 10), 1071 => to_unsigned(538, 10), 1072 => to_unsigned(483, 10), 1073 => to_unsigned(453, 10), 1074 => to_unsigned(488, 10), 1075 => to_unsigned(438, 10), 1076 => to_unsigned(526, 10), 1077 => to_unsigned(509, 10), 1078 => to_unsigned(618, 10), 1079 => to_unsigned(397, 10), 1080 => to_unsigned(349, 10), 1081 => to_unsigned(449, 10), 1082 => to_unsigned(450, 10), 1083 => to_unsigned(571, 10), 1084 => to_unsigned(478, 10), 1085 => to_unsigned(598, 10), 1086 => to_unsigned(429, 10), 1087 => to_unsigned(502, 10), 1088 => to_unsigned(397, 10), 1089 => to_unsigned(433, 10), 1090 => to_unsigned(589, 10), 1091 => to_unsigned(512, 10), 1092 => to_unsigned(420, 10), 1093 => to_unsigned(350, 10), 1094 => to_unsigned(464, 10), 1095 => to_unsigned(566, 10), 1096 => to_unsigned(448, 10), 1097 => to_unsigned(537, 10), 1098 => to_unsigned(351, 10), 1099 => to_unsigned(459, 10), 1100 => to_unsigned(518, 10), 1101 => to_unsigned(522, 10), 1102 => to_unsigned(637, 10), 1103 => to_unsigned(561, 10), 1104 => to_unsigned(561, 10), 1105 => to_unsigned(597, 10), 1106 => to_unsigned(591, 10), 1107 => to_unsigned(579, 10), 1108 => to_unsigned(391, 10), 1109 => to_unsigned(389, 10), 1110 => to_unsigned(361, 10), 1111 => to_unsigned(534, 10), 1112 => to_unsigned(664, 10), 1113 => to_unsigned(476, 10), 1114 => to_unsigned(686, 10), 1115 => to_unsigned(523, 10), 1116 => to_unsigned(518, 10), 1117 => to_unsigned(655, 10), 1118 => to_unsigned(501, 10), 1119 => to_unsigned(534, 10), 1120 => to_unsigned(451, 10), 1121 => to_unsigned(765, 10), 1122 => to_unsigned(686, 10), 1123 => to_unsigned(524, 10), 1124 => to_unsigned(338, 10), 1125 => to_unsigned(483, 10), 1126 => to_unsigned(477, 10), 1127 => to_unsigned(582, 10), 1128 => to_unsigned(517, 10), 1129 => to_unsigned(487, 10), 1130 => to_unsigned(536, 10), 1131 => to_unsigned(310, 10), 1132 => to_unsigned(472, 10), 1133 => to_unsigned(469, 10), 1134 => to_unsigned(664, 10), 1135 => to_unsigned(291, 10), 1136 => to_unsigned(665, 10), 1137 => to_unsigned(631, 10), 1138 => to_unsigned(569, 10), 1139 => to_unsigned(457, 10), 1140 => to_unsigned(555, 10), 1141 => to_unsigned(458, 10), 1142 => to_unsigned(495, 10), 1143 => to_unsigned(512, 10), 1144 => to_unsigned(501, 10), 1145 => to_unsigned(562, 10), 1146 => to_unsigned(386, 10), 1147 => to_unsigned(509, 10), 1148 => to_unsigned(659, 10), 1149 => to_unsigned(669, 10), 1150 => to_unsigned(536, 10), 1151 => to_unsigned(378, 10), 1152 => to_unsigned(553, 10), 1153 => to_unsigned(629, 10), 1154 => to_unsigned(573, 10), 1155 => to_unsigned(504, 10), 1156 => to_unsigned(509, 10), 1157 => to_unsigned(456, 10), 1158 => to_unsigned(406, 10), 1159 => to_unsigned(594, 10), 1160 => to_unsigned(458, 10), 1161 => to_unsigned(643, 10), 1162 => to_unsigned(515, 10), 1163 => to_unsigned(408, 10), 1164 => to_unsigned(495, 10), 1165 => to_unsigned(424, 10), 1166 => to_unsigned(552, 10), 1167 => to_unsigned(468, 10), 1168 => to_unsigned(463, 10), 1169 => to_unsigned(635, 10), 1170 => to_unsigned(388, 10), 1171 => to_unsigned(519, 10), 1172 => to_unsigned(583, 10), 1173 => to_unsigned(538, 10), 1174 => to_unsigned(456, 10), 1175 => to_unsigned(412, 10), 1176 => to_unsigned(606, 10), 1177 => to_unsigned(596, 10), 1178 => to_unsigned(609, 10), 1179 => to_unsigned(496, 10), 1180 => to_unsigned(404, 10), 1181 => to_unsigned(457, 10), 1182 => to_unsigned(453, 10), 1183 => to_unsigned(454, 10), 1184 => to_unsigned(574, 10), 1185 => to_unsigned(459, 10), 1186 => to_unsigned(572, 10), 1187 => to_unsigned(488, 10), 1188 => to_unsigned(619, 10), 1189 => to_unsigned(404, 10), 1190 => to_unsigned(510, 10), 1191 => to_unsigned(585, 10), 1192 => to_unsigned(272, 10), 1193 => to_unsigned(372, 10), 1194 => to_unsigned(488, 10), 1195 => to_unsigned(694, 10), 1196 => to_unsigned(429, 10), 1197 => to_unsigned(599, 10), 1198 => to_unsigned(453, 10), 1199 => to_unsigned(393, 10), 1200 => to_unsigned(519, 10), 1201 => to_unsigned(590, 10), 1202 => to_unsigned(467, 10), 1203 => to_unsigned(497, 10), 1204 => to_unsigned(384, 10), 1205 => to_unsigned(674, 10), 1206 => to_unsigned(561, 10), 1207 => to_unsigned(484, 10), 1208 => to_unsigned(507, 10), 1209 => to_unsigned(633, 10), 1210 => to_unsigned(623, 10), 1211 => to_unsigned(493, 10), 1212 => to_unsigned(568, 10), 1213 => to_unsigned(464, 10), 1214 => to_unsigned(537, 10), 1215 => to_unsigned(580, 10), 1216 => to_unsigned(508, 10), 1217 => to_unsigned(481, 10), 1218 => to_unsigned(466, 10), 1219 => to_unsigned(650, 10), 1220 => to_unsigned(542, 10), 1221 => to_unsigned(464, 10), 1222 => to_unsigned(388, 10), 1223 => to_unsigned(561, 10), 1224 => to_unsigned(552, 10), 1225 => to_unsigned(449, 10), 1226 => to_unsigned(508, 10), 1227 => to_unsigned(364, 10), 1228 => to_unsigned(430, 10), 1229 => to_unsigned(650, 10), 1230 => to_unsigned(617, 10), 1231 => to_unsigned(495, 10), 1232 => to_unsigned(607, 10), 1233 => to_unsigned(558, 10), 1234 => to_unsigned(462, 10), 1235 => to_unsigned(492, 10), 1236 => to_unsigned(531, 10), 1237 => to_unsigned(470, 10), 1238 => to_unsigned(613, 10), 1239 => to_unsigned(514, 10), 1240 => to_unsigned(353, 10), 1241 => to_unsigned(469, 10), 1242 => to_unsigned(537, 10), 1243 => to_unsigned(592, 10), 1244 => to_unsigned(499, 10), 1245 => to_unsigned(655, 10), 1246 => to_unsigned(444, 10), 1247 => to_unsigned(490, 10), 1248 => to_unsigned(395, 10), 1249 => to_unsigned(577, 10), 1250 => to_unsigned(439, 10), 1251 => to_unsigned(557, 10), 1252 => to_unsigned(466, 10), 1253 => to_unsigned(501, 10), 1254 => to_unsigned(545, 10), 1255 => to_unsigned(503, 10), 1256 => to_unsigned(460, 10), 1257 => to_unsigned(424, 10), 1258 => to_unsigned(468, 10), 1259 => to_unsigned(578, 10), 1260 => to_unsigned(662, 10), 1261 => to_unsigned(384, 10), 1262 => to_unsigned(399, 10), 1263 => to_unsigned(455, 10), 1264 => to_unsigned(624, 10), 1265 => to_unsigned(487, 10), 1266 => to_unsigned(529, 10), 1267 => to_unsigned(469, 10), 1268 => to_unsigned(546, 10), 1269 => to_unsigned(530, 10), 1270 => to_unsigned(666, 10), 1271 => to_unsigned(477, 10), 1272 => to_unsigned(488, 10), 1273 => to_unsigned(360, 10), 1274 => to_unsigned(677, 10), 1275 => to_unsigned(369, 10), 1276 => to_unsigned(751, 10), 1277 => to_unsigned(525, 10), 1278 => to_unsigned(518, 10), 1279 => to_unsigned(493, 10), 1280 => to_unsigned(550, 10), 1281 => to_unsigned(514, 10), 1282 => to_unsigned(609, 10), 1283 => to_unsigned(519, 10), 1284 => to_unsigned(495, 10), 1285 => to_unsigned(412, 10), 1286 => to_unsigned(584, 10), 1287 => to_unsigned(520, 10), 1288 => to_unsigned(433, 10), 1289 => to_unsigned(462, 10), 1290 => to_unsigned(618, 10), 1291 => to_unsigned(596, 10), 1292 => to_unsigned(406, 10), 1293 => to_unsigned(533, 10), 1294 => to_unsigned(554, 10), 1295 => to_unsigned(520, 10), 1296 => to_unsigned(471, 10), 1297 => to_unsigned(470, 10), 1298 => to_unsigned(486, 10), 1299 => to_unsigned(640, 10), 1300 => to_unsigned(550, 10), 1301 => to_unsigned(410, 10), 1302 => to_unsigned(520, 10), 1303 => to_unsigned(444, 10), 1304 => to_unsigned(417, 10), 1305 => to_unsigned(496, 10), 1306 => to_unsigned(650, 10), 1307 => to_unsigned(476, 10), 1308 => to_unsigned(351, 10), 1309 => to_unsigned(454, 10), 1310 => to_unsigned(404, 10), 1311 => to_unsigned(538, 10), 1312 => to_unsigned(479, 10), 1313 => to_unsigned(555, 10), 1314 => to_unsigned(449, 10), 1315 => to_unsigned(428, 10), 1316 => to_unsigned(411, 10), 1317 => to_unsigned(574, 10), 1318 => to_unsigned(654, 10), 1319 => to_unsigned(394, 10), 1320 => to_unsigned(431, 10), 1321 => to_unsigned(504, 10), 1322 => to_unsigned(519, 10), 1323 => to_unsigned(344, 10), 1324 => to_unsigned(382, 10), 1325 => to_unsigned(642, 10), 1326 => to_unsigned(641, 10), 1327 => to_unsigned(424, 10), 1328 => to_unsigned(551, 10), 1329 => to_unsigned(499, 10), 1330 => to_unsigned(577, 10), 1331 => to_unsigned(653, 10), 1332 => to_unsigned(329, 10), 1333 => to_unsigned(490, 10), 1334 => to_unsigned(584, 10), 1335 => to_unsigned(642, 10), 1336 => to_unsigned(386, 10), 1337 => to_unsigned(582, 10), 1338 => to_unsigned(402, 10), 1339 => to_unsigned(502, 10), 1340 => to_unsigned(513, 10), 1341 => to_unsigned(408, 10), 1342 => to_unsigned(521, 10), 1343 => to_unsigned(743, 10), 1344 => to_unsigned(658, 10), 1345 => to_unsigned(522, 10), 1346 => to_unsigned(408, 10), 1347 => to_unsigned(483, 10), 1348 => to_unsigned(535, 10), 1349 => to_unsigned(488, 10), 1350 => to_unsigned(539, 10), 1351 => to_unsigned(489, 10), 1352 => to_unsigned(414, 10), 1353 => to_unsigned(643, 10), 1354 => to_unsigned(381, 10), 1355 => to_unsigned(405, 10), 1356 => to_unsigned(564, 10), 1357 => to_unsigned(555, 10), 1358 => to_unsigned(404, 10), 1359 => to_unsigned(504, 10), 1360 => to_unsigned(394, 10), 1361 => to_unsigned(366, 10), 1362 => to_unsigned(608, 10), 1363 => to_unsigned(543, 10), 1364 => to_unsigned(592, 10), 1365 => to_unsigned(537, 10), 1366 => to_unsigned(593, 10), 1367 => to_unsigned(523, 10), 1368 => to_unsigned(349, 10), 1369 => to_unsigned(446, 10), 1370 => to_unsigned(492, 10), 1371 => to_unsigned(440, 10), 1372 => to_unsigned(453, 10), 1373 => to_unsigned(555, 10), 1374 => to_unsigned(642, 10), 1375 => to_unsigned(540, 10), 1376 => to_unsigned(543, 10), 1377 => to_unsigned(362, 10), 1378 => to_unsigned(533, 10), 1379 => to_unsigned(308, 10), 1380 => to_unsigned(590, 10), 1381 => to_unsigned(426, 10), 1382 => to_unsigned(567, 10), 1383 => to_unsigned(560, 10), 1384 => to_unsigned(614, 10), 1385 => to_unsigned(396, 10), 1386 => to_unsigned(595, 10), 1387 => to_unsigned(540, 10), 1388 => to_unsigned(571, 10), 1389 => to_unsigned(433, 10), 1390 => to_unsigned(455, 10), 1391 => to_unsigned(423, 10), 1392 => to_unsigned(642, 10), 1393 => to_unsigned(533, 10), 1394 => to_unsigned(401, 10), 1395 => to_unsigned(485, 10), 1396 => to_unsigned(380, 10), 1397 => to_unsigned(546, 10), 1398 => to_unsigned(243, 10), 1399 => to_unsigned(605, 10), 1400 => to_unsigned(509, 10), 1401 => to_unsigned(663, 10), 1402 => to_unsigned(390, 10), 1403 => to_unsigned(516, 10), 1404 => to_unsigned(271, 10), 1405 => to_unsigned(540, 10), 1406 => to_unsigned(514, 10), 1407 => to_unsigned(557, 10), 1408 => to_unsigned(399, 10), 1409 => to_unsigned(584, 10), 1410 => to_unsigned(351, 10), 1411 => to_unsigned(484, 10), 1412 => to_unsigned(353, 10), 1413 => to_unsigned(497, 10), 1414 => to_unsigned(600, 10), 1415 => to_unsigned(365, 10), 1416 => to_unsigned(623, 10), 1417 => to_unsigned(405, 10), 1418 => to_unsigned(293, 10), 1419 => to_unsigned(375, 10), 1420 => to_unsigned(503, 10), 1421 => to_unsigned(510, 10), 1422 => to_unsigned(376, 10), 1423 => to_unsigned(653, 10), 1424 => to_unsigned(517, 10), 1425 => to_unsigned(497, 10), 1426 => to_unsigned(708, 10), 1427 => to_unsigned(700, 10), 1428 => to_unsigned(472, 10), 1429 => to_unsigned(561, 10), 1430 => to_unsigned(559, 10), 1431 => to_unsigned(471, 10), 1432 => to_unsigned(548, 10), 1433 => to_unsigned(606, 10), 1434 => to_unsigned(588, 10), 1435 => to_unsigned(469, 10), 1436 => to_unsigned(407, 10), 1437 => to_unsigned(402, 10), 1438 => to_unsigned(465, 10), 1439 => to_unsigned(440, 10), 1440 => to_unsigned(522, 10), 1441 => to_unsigned(407, 10), 1442 => to_unsigned(548, 10), 1443 => to_unsigned(517, 10), 1444 => to_unsigned(460, 10), 1445 => to_unsigned(571, 10), 1446 => to_unsigned(512, 10), 1447 => to_unsigned(563, 10), 1448 => to_unsigned(539, 10), 1449 => to_unsigned(518, 10), 1450 => to_unsigned(528, 10), 1451 => to_unsigned(567, 10), 1452 => to_unsigned(468, 10), 1453 => to_unsigned(431, 10), 1454 => to_unsigned(525, 10), 1455 => to_unsigned(619, 10), 1456 => to_unsigned(467, 10), 1457 => to_unsigned(691, 10), 1458 => to_unsigned(645, 10), 1459 => to_unsigned(453, 10), 1460 => to_unsigned(424, 10), 1461 => to_unsigned(532, 10), 1462 => to_unsigned(520, 10), 1463 => to_unsigned(486, 10), 1464 => to_unsigned(498, 10), 1465 => to_unsigned(465, 10), 1466 => to_unsigned(643, 10), 1467 => to_unsigned(321, 10), 1468 => to_unsigned(489, 10), 1469 => to_unsigned(538, 10), 1470 => to_unsigned(441, 10), 1471 => to_unsigned(400, 10), 1472 => to_unsigned(531, 10), 1473 => to_unsigned(583, 10), 1474 => to_unsigned(429, 10), 1475 => to_unsigned(488, 10), 1476 => to_unsigned(560, 10), 1477 => to_unsigned(531, 10), 1478 => to_unsigned(506, 10), 1479 => to_unsigned(422, 10), 1480 => to_unsigned(295, 10), 1481 => to_unsigned(432, 10), 1482 => to_unsigned(586, 10), 1483 => to_unsigned(556, 10), 1484 => to_unsigned(646, 10), 1485 => to_unsigned(459, 10), 1486 => to_unsigned(709, 10), 1487 => to_unsigned(376, 10), 1488 => to_unsigned(601, 10), 1489 => to_unsigned(622, 10), 1490 => to_unsigned(548, 10), 1491 => to_unsigned(502, 10), 1492 => to_unsigned(501, 10), 1493 => to_unsigned(597, 10), 1494 => to_unsigned(524, 10), 1495 => to_unsigned(589, 10), 1496 => to_unsigned(551, 10), 1497 => to_unsigned(521, 10), 1498 => to_unsigned(488, 10), 1499 => to_unsigned(581, 10), 1500 => to_unsigned(643, 10), 1501 => to_unsigned(401, 10), 1502 => to_unsigned(471, 10), 1503 => to_unsigned(390, 10), 1504 => to_unsigned(477, 10), 1505 => to_unsigned(382, 10), 1506 => to_unsigned(494, 10), 1507 => to_unsigned(701, 10), 1508 => to_unsigned(509, 10), 1509 => to_unsigned(505, 10), 1510 => to_unsigned(511, 10), 1511 => to_unsigned(480, 10), 1512 => to_unsigned(669, 10), 1513 => to_unsigned(612, 10), 1514 => to_unsigned(383, 10), 1515 => to_unsigned(444, 10), 1516 => to_unsigned(450, 10), 1517 => to_unsigned(553, 10), 1518 => to_unsigned(440, 10), 1519 => to_unsigned(595, 10), 1520 => to_unsigned(455, 10), 1521 => to_unsigned(392, 10), 1522 => to_unsigned(483, 10), 1523 => to_unsigned(554, 10), 1524 => to_unsigned(586, 10), 1525 => to_unsigned(434, 10), 1526 => to_unsigned(450, 10), 1527 => to_unsigned(435, 10), 1528 => to_unsigned(550, 10), 1529 => to_unsigned(476, 10), 1530 => to_unsigned(519, 10), 1531 => to_unsigned(678, 10), 1532 => to_unsigned(486, 10), 1533 => to_unsigned(357, 10), 1534 => to_unsigned(486, 10), 1535 => to_unsigned(488, 10), 1536 => to_unsigned(481, 10), 1537 => to_unsigned(669, 10), 1538 => to_unsigned(529, 10), 1539 => to_unsigned(571, 10), 1540 => to_unsigned(418, 10), 1541 => to_unsigned(606, 10), 1542 => to_unsigned(646, 10), 1543 => to_unsigned(409, 10), 1544 => to_unsigned(587, 10), 1545 => to_unsigned(392, 10), 1546 => to_unsigned(428, 10), 1547 => to_unsigned(605, 10), 1548 => to_unsigned(499, 10), 1549 => to_unsigned(498, 10), 1550 => to_unsigned(461, 10), 1551 => to_unsigned(437, 10), 1552 => to_unsigned(512, 10), 1553 => to_unsigned(617, 10), 1554 => to_unsigned(463, 10), 1555 => to_unsigned(364, 10), 1556 => to_unsigned(571, 10), 1557 => to_unsigned(564, 10), 1558 => to_unsigned(293, 10), 1559 => to_unsigned(548, 10), 1560 => to_unsigned(486, 10), 1561 => to_unsigned(591, 10), 1562 => to_unsigned(568, 10), 1563 => to_unsigned(404, 10), 1564 => to_unsigned(681, 10), 1565 => to_unsigned(364, 10), 1566 => to_unsigned(427, 10), 1567 => to_unsigned(504, 10), 1568 => to_unsigned(625, 10), 1569 => to_unsigned(396, 10), 1570 => to_unsigned(557, 10), 1571 => to_unsigned(568, 10), 1572 => to_unsigned(499, 10), 1573 => to_unsigned(625, 10), 1574 => to_unsigned(512, 10), 1575 => to_unsigned(707, 10), 1576 => to_unsigned(583, 10), 1577 => to_unsigned(563, 10), 1578 => to_unsigned(420, 10), 1579 => to_unsigned(405, 10), 1580 => to_unsigned(306, 10), 1581 => to_unsigned(475, 10), 1582 => to_unsigned(467, 10), 1583 => to_unsigned(664, 10), 1584 => to_unsigned(483, 10), 1585 => to_unsigned(394, 10), 1586 => to_unsigned(580, 10), 1587 => to_unsigned(517, 10), 1588 => to_unsigned(514, 10), 1589 => to_unsigned(334, 10), 1590 => to_unsigned(494, 10), 1591 => to_unsigned(502, 10), 1592 => to_unsigned(543, 10), 1593 => to_unsigned(510, 10), 1594 => to_unsigned(554, 10), 1595 => to_unsigned(613, 10), 1596 => to_unsigned(455, 10), 1597 => to_unsigned(531, 10), 1598 => to_unsigned(438, 10), 1599 => to_unsigned(685, 10), 1600 => to_unsigned(547, 10), 1601 => to_unsigned(496, 10), 1602 => to_unsigned(611, 10), 1603 => to_unsigned(414, 10), 1604 => to_unsigned(497, 10), 1605 => to_unsigned(610, 10), 1606 => to_unsigned(542, 10), 1607 => to_unsigned(380, 10), 1608 => to_unsigned(643, 10), 1609 => to_unsigned(660, 10), 1610 => to_unsigned(603, 10), 1611 => to_unsigned(462, 10), 1612 => to_unsigned(510, 10), 1613 => to_unsigned(429, 10), 1614 => to_unsigned(611, 10), 1615 => to_unsigned(686, 10), 1616 => to_unsigned(375, 10), 1617 => to_unsigned(422, 10), 1618 => to_unsigned(591, 10), 1619 => to_unsigned(563, 10), 1620 => to_unsigned(432, 10), 1621 => to_unsigned(497, 10), 1622 => to_unsigned(653, 10), 1623 => to_unsigned(299, 10), 1624 => to_unsigned(489, 10), 1625 => to_unsigned(484, 10), 1626 => to_unsigned(445, 10), 1627 => to_unsigned(582, 10), 1628 => to_unsigned(567, 10), 1629 => to_unsigned(621, 10), 1630 => to_unsigned(469, 10), 1631 => to_unsigned(571, 10), 1632 => to_unsigned(428, 10), 1633 => to_unsigned(632, 10), 1634 => to_unsigned(617, 10), 1635 => to_unsigned(512, 10), 1636 => to_unsigned(588, 10), 1637 => to_unsigned(527, 10), 1638 => to_unsigned(333, 10), 1639 => to_unsigned(660, 10), 1640 => to_unsigned(429, 10), 1641 => to_unsigned(636, 10), 1642 => to_unsigned(508, 10), 1643 => to_unsigned(616, 10), 1644 => to_unsigned(398, 10), 1645 => to_unsigned(468, 10), 1646 => to_unsigned(477, 10), 1647 => to_unsigned(595, 10), 1648 => to_unsigned(514, 10), 1649 => to_unsigned(414, 10), 1650 => to_unsigned(673, 10), 1651 => to_unsigned(588, 10), 1652 => to_unsigned(408, 10), 1653 => to_unsigned(446, 10), 1654 => to_unsigned(626, 10), 1655 => to_unsigned(431, 10), 1656 => to_unsigned(432, 10), 1657 => to_unsigned(369, 10), 1658 => to_unsigned(544, 10), 1659 => to_unsigned(524, 10), 1660 => to_unsigned(495, 10), 1661 => to_unsigned(516, 10), 1662 => to_unsigned(421, 10), 1663 => to_unsigned(309, 10), 1664 => to_unsigned(378, 10), 1665 => to_unsigned(363, 10), 1666 => to_unsigned(565, 10), 1667 => to_unsigned(762, 10), 1668 => to_unsigned(438, 10), 1669 => to_unsigned(478, 10), 1670 => to_unsigned(675, 10), 1671 => to_unsigned(502, 10), 1672 => to_unsigned(583, 10), 1673 => to_unsigned(525, 10), 1674 => to_unsigned(573, 10), 1675 => to_unsigned(633, 10), 1676 => to_unsigned(439, 10), 1677 => to_unsigned(632, 10), 1678 => to_unsigned(617, 10), 1679 => to_unsigned(530, 10), 1680 => to_unsigned(498, 10), 1681 => to_unsigned(537, 10), 1682 => to_unsigned(559, 10), 1683 => to_unsigned(507, 10), 1684 => to_unsigned(342, 10), 1685 => to_unsigned(399, 10), 1686 => to_unsigned(703, 10), 1687 => to_unsigned(530, 10), 1688 => to_unsigned(340, 10), 1689 => to_unsigned(378, 10), 1690 => to_unsigned(477, 10), 1691 => to_unsigned(551, 10), 1692 => to_unsigned(401, 10), 1693 => to_unsigned(506, 10), 1694 => to_unsigned(400, 10), 1695 => to_unsigned(410, 10), 1696 => to_unsigned(435, 10), 1697 => to_unsigned(523, 10), 1698 => to_unsigned(649, 10), 1699 => to_unsigned(434, 10), 1700 => to_unsigned(540, 10), 1701 => to_unsigned(517, 10), 1702 => to_unsigned(442, 10), 1703 => to_unsigned(676, 10), 1704 => to_unsigned(489, 10), 1705 => to_unsigned(406, 10), 1706 => to_unsigned(293, 10), 1707 => to_unsigned(439, 10), 1708 => to_unsigned(723, 10), 1709 => to_unsigned(456, 10), 1710 => to_unsigned(506, 10), 1711 => to_unsigned(622, 10), 1712 => to_unsigned(485, 10), 1713 => to_unsigned(534, 10), 1714 => to_unsigned(560, 10), 1715 => to_unsigned(580, 10), 1716 => to_unsigned(510, 10), 1717 => to_unsigned(669, 10), 1718 => to_unsigned(484, 10), 1719 => to_unsigned(598, 10), 1720 => to_unsigned(646, 10), 1721 => to_unsigned(451, 10), 1722 => to_unsigned(527, 10), 1723 => to_unsigned(596, 10), 1724 => to_unsigned(617, 10), 1725 => to_unsigned(404, 10), 1726 => to_unsigned(506, 10), 1727 => to_unsigned(523, 10), 1728 => to_unsigned(417, 10), 1729 => to_unsigned(419, 10), 1730 => to_unsigned(461, 10), 1731 => to_unsigned(575, 10), 1732 => to_unsigned(490, 10), 1733 => to_unsigned(293, 10), 1734 => to_unsigned(525, 10), 1735 => to_unsigned(532, 10), 1736 => to_unsigned(446, 10), 1737 => to_unsigned(646, 10), 1738 => to_unsigned(582, 10), 1739 => to_unsigned(626, 10), 1740 => to_unsigned(413, 10), 1741 => to_unsigned(654, 10), 1742 => to_unsigned(565, 10), 1743 => to_unsigned(554, 10), 1744 => to_unsigned(473, 10), 1745 => to_unsigned(671, 10), 1746 => to_unsigned(472, 10), 1747 => to_unsigned(627, 10), 1748 => to_unsigned(486, 10), 1749 => to_unsigned(564, 10), 1750 => to_unsigned(525, 10), 1751 => to_unsigned(510, 10), 1752 => to_unsigned(462, 10), 1753 => to_unsigned(628, 10), 1754 => to_unsigned(562, 10), 1755 => to_unsigned(592, 10), 1756 => to_unsigned(457, 10), 1757 => to_unsigned(554, 10), 1758 => to_unsigned(534, 10), 1759 => to_unsigned(619, 10), 1760 => to_unsigned(324, 10), 1761 => to_unsigned(390, 10), 1762 => to_unsigned(541, 10), 1763 => to_unsigned(447, 10), 1764 => to_unsigned(466, 10), 1765 => to_unsigned(587, 10), 1766 => to_unsigned(494, 10), 1767 => to_unsigned(522, 10), 1768 => to_unsigned(464, 10), 1769 => to_unsigned(507, 10), 1770 => to_unsigned(410, 10), 1771 => to_unsigned(398, 10), 1772 => to_unsigned(677, 10), 1773 => to_unsigned(502, 10), 1774 => to_unsigned(449, 10), 1775 => to_unsigned(181, 10), 1776 => to_unsigned(509, 10), 1777 => to_unsigned(523, 10), 1778 => to_unsigned(555, 10), 1779 => to_unsigned(608, 10), 1780 => to_unsigned(586, 10), 1781 => to_unsigned(520, 10), 1782 => to_unsigned(641, 10), 1783 => to_unsigned(471, 10), 1784 => to_unsigned(428, 10), 1785 => to_unsigned(579, 10), 1786 => to_unsigned(603, 10), 1787 => to_unsigned(486, 10), 1788 => to_unsigned(521, 10), 1789 => to_unsigned(611, 10), 1790 => to_unsigned(564, 10), 1791 => to_unsigned(486, 10), 1792 => to_unsigned(496, 10), 1793 => to_unsigned(428, 10), 1794 => to_unsigned(533, 10), 1795 => to_unsigned(395, 10), 1796 => to_unsigned(472, 10), 1797 => to_unsigned(484, 10), 1798 => to_unsigned(501, 10), 1799 => to_unsigned(473, 10), 1800 => to_unsigned(597, 10), 1801 => to_unsigned(576, 10), 1802 => to_unsigned(468, 10), 1803 => to_unsigned(382, 10), 1804 => to_unsigned(594, 10), 1805 => to_unsigned(597, 10), 1806 => to_unsigned(602, 10), 1807 => to_unsigned(493, 10), 1808 => to_unsigned(395, 10), 1809 => to_unsigned(418, 10), 1810 => to_unsigned(572, 10), 1811 => to_unsigned(471, 10), 1812 => to_unsigned(560, 10), 1813 => to_unsigned(521, 10), 1814 => to_unsigned(491, 10), 1815 => to_unsigned(566, 10), 1816 => to_unsigned(594, 10), 1817 => to_unsigned(732, 10), 1818 => to_unsigned(482, 10), 1819 => to_unsigned(505, 10), 1820 => to_unsigned(409, 10), 1821 => to_unsigned(549, 10), 1822 => to_unsigned(625, 10), 1823 => to_unsigned(603, 10), 1824 => to_unsigned(637, 10), 1825 => to_unsigned(530, 10), 1826 => to_unsigned(364, 10), 1827 => to_unsigned(615, 10), 1828 => to_unsigned(423, 10), 1829 => to_unsigned(456, 10), 1830 => to_unsigned(543, 10), 1831 => to_unsigned(609, 10), 1832 => to_unsigned(555, 10), 1833 => to_unsigned(670, 10), 1834 => to_unsigned(470, 10), 1835 => to_unsigned(454, 10), 1836 => to_unsigned(621, 10), 1837 => to_unsigned(613, 10), 1838 => to_unsigned(484, 10), 1839 => to_unsigned(434, 10), 1840 => to_unsigned(531, 10), 1841 => to_unsigned(467, 10), 1842 => to_unsigned(508, 10), 1843 => to_unsigned(353, 10), 1844 => to_unsigned(520, 10), 1845 => to_unsigned(698, 10), 1846 => to_unsigned(634, 10), 1847 => to_unsigned(608, 10), 1848 => to_unsigned(466, 10), 1849 => to_unsigned(297, 10), 1850 => to_unsigned(493, 10), 1851 => to_unsigned(430, 10), 1852 => to_unsigned(560, 10), 1853 => to_unsigned(679, 10), 1854 => to_unsigned(566, 10), 1855 => to_unsigned(601, 10), 1856 => to_unsigned(518, 10), 1857 => to_unsigned(751, 10), 1858 => to_unsigned(550, 10), 1859 => to_unsigned(524, 10), 1860 => to_unsigned(569, 10), 1861 => to_unsigned(604, 10), 1862 => to_unsigned(390, 10), 1863 => to_unsigned(478, 10), 1864 => to_unsigned(434, 10), 1865 => to_unsigned(596, 10), 1866 => to_unsigned(484, 10), 1867 => to_unsigned(554, 10), 1868 => to_unsigned(486, 10), 1869 => to_unsigned(706, 10), 1870 => to_unsigned(447, 10), 1871 => to_unsigned(471, 10), 1872 => to_unsigned(405, 10), 1873 => to_unsigned(586, 10), 1874 => to_unsigned(666, 10), 1875 => to_unsigned(472, 10), 1876 => to_unsigned(484, 10), 1877 => to_unsigned(721, 10), 1878 => to_unsigned(572, 10), 1879 => to_unsigned(608, 10), 1880 => to_unsigned(544, 10), 1881 => to_unsigned(555, 10), 1882 => to_unsigned(551, 10), 1883 => to_unsigned(320, 10), 1884 => to_unsigned(521, 10), 1885 => to_unsigned(516, 10), 1886 => to_unsigned(546, 10), 1887 => to_unsigned(308, 10), 1888 => to_unsigned(603, 10), 1889 => to_unsigned(556, 10), 1890 => to_unsigned(435, 10), 1891 => to_unsigned(454, 10), 1892 => to_unsigned(547, 10), 1893 => to_unsigned(461, 10), 1894 => to_unsigned(472, 10), 1895 => to_unsigned(380, 10), 1896 => to_unsigned(406, 10), 1897 => to_unsigned(416, 10), 1898 => to_unsigned(459, 10), 1899 => to_unsigned(567, 10), 1900 => to_unsigned(478, 10), 1901 => to_unsigned(585, 10), 1902 => to_unsigned(578, 10), 1903 => to_unsigned(550, 10), 1904 => to_unsigned(607, 10), 1905 => to_unsigned(448, 10), 1906 => to_unsigned(478, 10), 1907 => to_unsigned(412, 10), 1908 => to_unsigned(418, 10), 1909 => to_unsigned(432, 10), 1910 => to_unsigned(658, 10), 1911 => to_unsigned(502, 10), 1912 => to_unsigned(615, 10), 1913 => to_unsigned(366, 10), 1914 => to_unsigned(436, 10), 1915 => to_unsigned(500, 10), 1916 => to_unsigned(587, 10), 1917 => to_unsigned(468, 10), 1918 => to_unsigned(320, 10), 1919 => to_unsigned(471, 10), 1920 => to_unsigned(375, 10), 1921 => to_unsigned(522, 10), 1922 => to_unsigned(385, 10), 1923 => to_unsigned(515, 10), 1924 => to_unsigned(520, 10), 1925 => to_unsigned(468, 10), 1926 => to_unsigned(406, 10), 1927 => to_unsigned(613, 10), 1928 => to_unsigned(734, 10), 1929 => to_unsigned(577, 10), 1930 => to_unsigned(439, 10), 1931 => to_unsigned(582, 10), 1932 => to_unsigned(301, 10), 1933 => to_unsigned(576, 10), 1934 => to_unsigned(537, 10), 1935 => to_unsigned(717, 10), 1936 => to_unsigned(457, 10), 1937 => to_unsigned(343, 10), 1938 => to_unsigned(397, 10), 1939 => to_unsigned(538, 10), 1940 => to_unsigned(451, 10), 1941 => to_unsigned(565, 10), 1942 => to_unsigned(648, 10), 1943 => to_unsigned(493, 10), 1944 => to_unsigned(569, 10), 1945 => to_unsigned(732, 10), 1946 => to_unsigned(274, 10), 1947 => to_unsigned(653, 10), 1948 => to_unsigned(573, 10), 1949 => to_unsigned(651, 10), 1950 => to_unsigned(370, 10), 1951 => to_unsigned(330, 10), 1952 => to_unsigned(551, 10), 1953 => to_unsigned(434, 10), 1954 => to_unsigned(672, 10), 1955 => to_unsigned(661, 10), 1956 => to_unsigned(344, 10), 1957 => to_unsigned(369, 10), 1958 => to_unsigned(523, 10), 1959 => to_unsigned(575, 10), 1960 => to_unsigned(575, 10), 1961 => to_unsigned(725, 10), 1962 => to_unsigned(502, 10), 1963 => to_unsigned(474, 10), 1964 => to_unsigned(367, 10), 1965 => to_unsigned(461, 10), 1966 => to_unsigned(700, 10), 1967 => to_unsigned(564, 10), 1968 => to_unsigned(508, 10), 1969 => to_unsigned(579, 10), 1970 => to_unsigned(489, 10), 1971 => to_unsigned(413, 10), 1972 => to_unsigned(551, 10), 1973 => to_unsigned(591, 10), 1974 => to_unsigned(464, 10), 1975 => to_unsigned(389, 10), 1976 => to_unsigned(410, 10), 1977 => to_unsigned(495, 10), 1978 => to_unsigned(490, 10), 1979 => to_unsigned(656, 10), 1980 => to_unsigned(524, 10), 1981 => to_unsigned(483, 10), 1982 => to_unsigned(521, 10), 1983 => to_unsigned(469, 10), 1984 => to_unsigned(617, 10), 1985 => to_unsigned(459, 10), 1986 => to_unsigned(406, 10), 1987 => to_unsigned(444, 10), 1988 => to_unsigned(462, 10), 1989 => to_unsigned(590, 10), 1990 => to_unsigned(532, 10), 1991 => to_unsigned(528, 10), 1992 => to_unsigned(452, 10), 1993 => to_unsigned(421, 10), 1994 => to_unsigned(506, 10), 1995 => to_unsigned(620, 10), 1996 => to_unsigned(403, 10), 1997 => to_unsigned(590, 10), 1998 => to_unsigned(433, 10), 1999 => to_unsigned(526, 10), 2000 => to_unsigned(348, 10), 2001 => to_unsigned(451, 10), 2002 => to_unsigned(421, 10), 2003 => to_unsigned(541, 10), 2004 => to_unsigned(362, 10), 2005 => to_unsigned(389, 10), 2006 => to_unsigned(532, 10), 2007 => to_unsigned(574, 10), 2008 => to_unsigned(496, 10), 2009 => to_unsigned(597, 10), 2010 => to_unsigned(388, 10), 2011 => to_unsigned(439, 10), 2012 => to_unsigned(354, 10), 2013 => to_unsigned(533, 10), 2014 => to_unsigned(513, 10), 2015 => to_unsigned(585, 10), 2016 => to_unsigned(515, 10), 2017 => to_unsigned(616, 10), 2018 => to_unsigned(441, 10), 2019 => to_unsigned(412, 10), 2020 => to_unsigned(436, 10), 2021 => to_unsigned(469, 10), 2022 => to_unsigned(550, 10), 2023 => to_unsigned(388, 10), 2024 => to_unsigned(412, 10), 2025 => to_unsigned(424, 10), 2026 => to_unsigned(681, 10), 2027 => to_unsigned(547, 10), 2028 => to_unsigned(636, 10), 2029 => to_unsigned(516, 10), 2030 => to_unsigned(642, 10), 2031 => to_unsigned(608, 10), 2032 => to_unsigned(584, 10), 2033 => to_unsigned(456, 10), 2034 => to_unsigned(356, 10), 2035 => to_unsigned(459, 10), 2036 => to_unsigned(498, 10), 2037 => to_unsigned(517, 10), 2038 => to_unsigned(402, 10), 2039 => to_unsigned(521, 10), 2040 => to_unsigned(433, 10), 2041 => to_unsigned(570, 10), 2042 => to_unsigned(589, 10), 2043 => to_unsigned(464, 10), 2044 => to_unsigned(374, 10), 2045 => to_unsigned(508, 10), 2046 => to_unsigned(322, 10), 2047 => to_unsigned(499, 10)),
        1 => (0 => to_unsigned(405, 10), 1 => to_unsigned(361, 10), 2 => to_unsigned(493, 10), 3 => to_unsigned(501, 10), 4 => to_unsigned(567, 10), 5 => to_unsigned(532, 10), 6 => to_unsigned(492, 10), 7 => to_unsigned(376, 10), 8 => to_unsigned(633, 10), 9 => to_unsigned(598, 10), 10 => to_unsigned(336, 10), 11 => to_unsigned(543, 10), 12 => to_unsigned(442, 10), 13 => to_unsigned(415, 10), 14 => to_unsigned(443, 10), 15 => to_unsigned(549, 10), 16 => to_unsigned(643, 10), 17 => to_unsigned(560, 10), 18 => to_unsigned(599, 10), 19 => to_unsigned(579, 10), 20 => to_unsigned(617, 10), 21 => to_unsigned(599, 10), 22 => to_unsigned(496, 10), 23 => to_unsigned(591, 10), 24 => to_unsigned(578, 10), 25 => to_unsigned(379, 10), 26 => to_unsigned(638, 10), 27 => to_unsigned(459, 10), 28 => to_unsigned(620, 10), 29 => to_unsigned(376, 10), 30 => to_unsigned(543, 10), 31 => to_unsigned(513, 10), 32 => to_unsigned(474, 10), 33 => to_unsigned(306, 10), 34 => to_unsigned(464, 10), 35 => to_unsigned(618, 10), 36 => to_unsigned(542, 10), 37 => to_unsigned(422, 10), 38 => to_unsigned(589, 10), 39 => to_unsigned(496, 10), 40 => to_unsigned(603, 10), 41 => to_unsigned(424, 10), 42 => to_unsigned(458, 10), 43 => to_unsigned(653, 10), 44 => to_unsigned(618, 10), 45 => to_unsigned(527, 10), 46 => to_unsigned(543, 10), 47 => to_unsigned(472, 10), 48 => to_unsigned(526, 10), 49 => to_unsigned(490, 10), 50 => to_unsigned(540, 10), 51 => to_unsigned(545, 10), 52 => to_unsigned(409, 10), 53 => to_unsigned(597, 10), 54 => to_unsigned(470, 10), 55 => to_unsigned(603, 10), 56 => to_unsigned(518, 10), 57 => to_unsigned(443, 10), 58 => to_unsigned(468, 10), 59 => to_unsigned(466, 10), 60 => to_unsigned(427, 10), 61 => to_unsigned(543, 10), 62 => to_unsigned(564, 10), 63 => to_unsigned(609, 10), 64 => to_unsigned(582, 10), 65 => to_unsigned(455, 10), 66 => to_unsigned(495, 10), 67 => to_unsigned(253, 10), 68 => to_unsigned(413, 10), 69 => to_unsigned(561, 10), 70 => to_unsigned(451, 10), 71 => to_unsigned(500, 10), 72 => to_unsigned(433, 10), 73 => to_unsigned(349, 10), 74 => to_unsigned(471, 10), 75 => to_unsigned(630, 10), 76 => to_unsigned(488, 10), 77 => to_unsigned(427, 10), 78 => to_unsigned(511, 10), 79 => to_unsigned(498, 10), 80 => to_unsigned(533, 10), 81 => to_unsigned(585, 10), 82 => to_unsigned(527, 10), 83 => to_unsigned(545, 10), 84 => to_unsigned(678, 10), 85 => to_unsigned(530, 10), 86 => to_unsigned(523, 10), 87 => to_unsigned(501, 10), 88 => to_unsigned(629, 10), 89 => to_unsigned(569, 10), 90 => to_unsigned(633, 10), 91 => to_unsigned(371, 10), 92 => to_unsigned(496, 10), 93 => to_unsigned(515, 10), 94 => to_unsigned(500, 10), 95 => to_unsigned(712, 10), 96 => to_unsigned(501, 10), 97 => to_unsigned(548, 10), 98 => to_unsigned(501, 10), 99 => to_unsigned(488, 10), 100 => to_unsigned(530, 10), 101 => to_unsigned(652, 10), 102 => to_unsigned(376, 10), 103 => to_unsigned(580, 10), 104 => to_unsigned(401, 10), 105 => to_unsigned(432, 10), 106 => to_unsigned(453, 10), 107 => to_unsigned(358, 10), 108 => to_unsigned(567, 10), 109 => to_unsigned(574, 10), 110 => to_unsigned(388, 10), 111 => to_unsigned(545, 10), 112 => to_unsigned(360, 10), 113 => to_unsigned(632, 10), 114 => to_unsigned(465, 10), 115 => to_unsigned(426, 10), 116 => to_unsigned(491, 10), 117 => to_unsigned(658, 10), 118 => to_unsigned(538, 10), 119 => to_unsigned(669, 10), 120 => to_unsigned(458, 10), 121 => to_unsigned(383, 10), 122 => to_unsigned(429, 10), 123 => to_unsigned(509, 10), 124 => to_unsigned(654, 10), 125 => to_unsigned(535, 10), 126 => to_unsigned(539, 10), 127 => to_unsigned(497, 10), 128 => to_unsigned(535, 10), 129 => to_unsigned(491, 10), 130 => to_unsigned(560, 10), 131 => to_unsigned(542, 10), 132 => to_unsigned(593, 10), 133 => to_unsigned(474, 10), 134 => to_unsigned(751, 10), 135 => to_unsigned(451, 10), 136 => to_unsigned(593, 10), 137 => to_unsigned(425, 10), 138 => to_unsigned(463, 10), 139 => to_unsigned(539, 10), 140 => to_unsigned(542, 10), 141 => to_unsigned(629, 10), 142 => to_unsigned(564, 10), 143 => to_unsigned(487, 10), 144 => to_unsigned(684, 10), 145 => to_unsigned(342, 10), 146 => to_unsigned(623, 10), 147 => to_unsigned(498, 10), 148 => to_unsigned(495, 10), 149 => to_unsigned(517, 10), 150 => to_unsigned(579, 10), 151 => to_unsigned(318, 10), 152 => to_unsigned(323, 10), 153 => to_unsigned(515, 10), 154 => to_unsigned(357, 10), 155 => to_unsigned(458, 10), 156 => to_unsigned(316, 10), 157 => to_unsigned(615, 10), 158 => to_unsigned(687, 10), 159 => to_unsigned(452, 10), 160 => to_unsigned(576, 10), 161 => to_unsigned(527, 10), 162 => to_unsigned(592, 10), 163 => to_unsigned(472, 10), 164 => to_unsigned(589, 10), 165 => to_unsigned(496, 10), 166 => to_unsigned(626, 10), 167 => to_unsigned(408, 10), 168 => to_unsigned(443, 10), 169 => to_unsigned(551, 10), 170 => to_unsigned(508, 10), 171 => to_unsigned(567, 10), 172 => to_unsigned(612, 10), 173 => to_unsigned(453, 10), 174 => to_unsigned(584, 10), 175 => to_unsigned(541, 10), 176 => to_unsigned(620, 10), 177 => to_unsigned(289, 10), 178 => to_unsigned(612, 10), 179 => to_unsigned(732, 10), 180 => to_unsigned(532, 10), 181 => to_unsigned(626, 10), 182 => to_unsigned(640, 10), 183 => to_unsigned(523, 10), 184 => to_unsigned(460, 10), 185 => to_unsigned(635, 10), 186 => to_unsigned(319, 10), 187 => to_unsigned(682, 10), 188 => to_unsigned(557, 10), 189 => to_unsigned(510, 10), 190 => to_unsigned(562, 10), 191 => to_unsigned(644, 10), 192 => to_unsigned(570, 10), 193 => to_unsigned(487, 10), 194 => to_unsigned(407, 10), 195 => to_unsigned(500, 10), 196 => to_unsigned(651, 10), 197 => to_unsigned(373, 10), 198 => to_unsigned(635, 10), 199 => to_unsigned(484, 10), 200 => to_unsigned(377, 10), 201 => to_unsigned(361, 10), 202 => to_unsigned(484, 10), 203 => to_unsigned(451, 10), 204 => to_unsigned(691, 10), 205 => to_unsigned(491, 10), 206 => to_unsigned(589, 10), 207 => to_unsigned(239, 10), 208 => to_unsigned(516, 10), 209 => to_unsigned(480, 10), 210 => to_unsigned(428, 10), 211 => to_unsigned(456, 10), 212 => to_unsigned(389, 10), 213 => to_unsigned(484, 10), 214 => to_unsigned(410, 10), 215 => to_unsigned(477, 10), 216 => to_unsigned(373, 10), 217 => to_unsigned(635, 10), 218 => to_unsigned(439, 10), 219 => to_unsigned(605, 10), 220 => to_unsigned(556, 10), 221 => to_unsigned(520, 10), 222 => to_unsigned(616, 10), 223 => to_unsigned(338, 10), 224 => to_unsigned(521, 10), 225 => to_unsigned(677, 10), 226 => to_unsigned(406, 10), 227 => to_unsigned(367, 10), 228 => to_unsigned(560, 10), 229 => to_unsigned(666, 10), 230 => to_unsigned(360, 10), 231 => to_unsigned(396, 10), 232 => to_unsigned(469, 10), 233 => to_unsigned(447, 10), 234 => to_unsigned(506, 10), 235 => to_unsigned(371, 10), 236 => to_unsigned(491, 10), 237 => to_unsigned(523, 10), 238 => to_unsigned(594, 10), 239 => to_unsigned(400, 10), 240 => to_unsigned(616, 10), 241 => to_unsigned(576, 10), 242 => to_unsigned(481, 10), 243 => to_unsigned(576, 10), 244 => to_unsigned(581, 10), 245 => to_unsigned(525, 10), 246 => to_unsigned(401, 10), 247 => to_unsigned(618, 10), 248 => to_unsigned(392, 10), 249 => to_unsigned(364, 10), 250 => to_unsigned(526, 10), 251 => to_unsigned(524, 10), 252 => to_unsigned(489, 10), 253 => to_unsigned(596, 10), 254 => to_unsigned(505, 10), 255 => to_unsigned(497, 10), 256 => to_unsigned(439, 10), 257 => to_unsigned(529, 10), 258 => to_unsigned(618, 10), 259 => to_unsigned(505, 10), 260 => to_unsigned(466, 10), 261 => to_unsigned(595, 10), 262 => to_unsigned(554, 10), 263 => to_unsigned(340, 10), 264 => to_unsigned(574, 10), 265 => to_unsigned(504, 10), 266 => to_unsigned(577, 10), 267 => to_unsigned(453, 10), 268 => to_unsigned(595, 10), 269 => to_unsigned(428, 10), 270 => to_unsigned(464, 10), 271 => to_unsigned(423, 10), 272 => to_unsigned(487, 10), 273 => to_unsigned(359, 10), 274 => to_unsigned(510, 10), 275 => to_unsigned(377, 10), 276 => to_unsigned(566, 10), 277 => to_unsigned(514, 10), 278 => to_unsigned(689, 10), 279 => to_unsigned(468, 10), 280 => to_unsigned(545, 10), 281 => to_unsigned(342, 10), 282 => to_unsigned(518, 10), 283 => to_unsigned(407, 10), 284 => to_unsigned(626, 10), 285 => to_unsigned(646, 10), 286 => to_unsigned(349, 10), 287 => to_unsigned(498, 10), 288 => to_unsigned(531, 10), 289 => to_unsigned(568, 10), 290 => to_unsigned(603, 10), 291 => to_unsigned(441, 10), 292 => to_unsigned(502, 10), 293 => to_unsigned(536, 10), 294 => to_unsigned(511, 10), 295 => to_unsigned(477, 10), 296 => to_unsigned(351, 10), 297 => to_unsigned(644, 10), 298 => to_unsigned(596, 10), 299 => to_unsigned(582, 10), 300 => to_unsigned(462, 10), 301 => to_unsigned(442, 10), 302 => to_unsigned(387, 10), 303 => to_unsigned(536, 10), 304 => to_unsigned(433, 10), 305 => to_unsigned(416, 10), 306 => to_unsigned(479, 10), 307 => to_unsigned(623, 10), 308 => to_unsigned(549, 10), 309 => to_unsigned(471, 10), 310 => to_unsigned(372, 10), 311 => to_unsigned(523, 10), 312 => to_unsigned(332, 10), 313 => to_unsigned(398, 10), 314 => to_unsigned(463, 10), 315 => to_unsigned(459, 10), 316 => to_unsigned(508, 10), 317 => to_unsigned(391, 10), 318 => to_unsigned(421, 10), 319 => to_unsigned(568, 10), 320 => to_unsigned(455, 10), 321 => to_unsigned(445, 10), 322 => to_unsigned(383, 10), 323 => to_unsigned(764, 10), 324 => to_unsigned(623, 10), 325 => to_unsigned(503, 10), 326 => to_unsigned(499, 10), 327 => to_unsigned(679, 10), 328 => to_unsigned(512, 10), 329 => to_unsigned(597, 10), 330 => to_unsigned(557, 10), 331 => to_unsigned(488, 10), 332 => to_unsigned(542, 10), 333 => to_unsigned(599, 10), 334 => to_unsigned(579, 10), 335 => to_unsigned(754, 10), 336 => to_unsigned(576, 10), 337 => to_unsigned(637, 10), 338 => to_unsigned(574, 10), 339 => to_unsigned(643, 10), 340 => to_unsigned(750, 10), 341 => to_unsigned(347, 10), 342 => to_unsigned(693, 10), 343 => to_unsigned(441, 10), 344 => to_unsigned(476, 10), 345 => to_unsigned(405, 10), 346 => to_unsigned(463, 10), 347 => to_unsigned(546, 10), 348 => to_unsigned(627, 10), 349 => to_unsigned(507, 10), 350 => to_unsigned(411, 10), 351 => to_unsigned(490, 10), 352 => to_unsigned(533, 10), 353 => to_unsigned(434, 10), 354 => to_unsigned(517, 10), 355 => to_unsigned(515, 10), 356 => to_unsigned(481, 10), 357 => to_unsigned(550, 10), 358 => to_unsigned(471, 10), 359 => to_unsigned(626, 10), 360 => to_unsigned(585, 10), 361 => to_unsigned(665, 10), 362 => to_unsigned(717, 10), 363 => to_unsigned(599, 10), 364 => to_unsigned(476, 10), 365 => to_unsigned(737, 10), 366 => to_unsigned(654, 10), 367 => to_unsigned(553, 10), 368 => to_unsigned(590, 10), 369 => to_unsigned(631, 10), 370 => to_unsigned(744, 10), 371 => to_unsigned(413, 10), 372 => to_unsigned(510, 10), 373 => to_unsigned(509, 10), 374 => to_unsigned(460, 10), 375 => to_unsigned(380, 10), 376 => to_unsigned(604, 10), 377 => to_unsigned(587, 10), 378 => to_unsigned(262, 10), 379 => to_unsigned(532, 10), 380 => to_unsigned(486, 10), 381 => to_unsigned(440, 10), 382 => to_unsigned(424, 10), 383 => to_unsigned(504, 10), 384 => to_unsigned(526, 10), 385 => to_unsigned(337, 10), 386 => to_unsigned(468, 10), 387 => to_unsigned(682, 10), 388 => to_unsigned(362, 10), 389 => to_unsigned(475, 10), 390 => to_unsigned(595, 10), 391 => to_unsigned(469, 10), 392 => to_unsigned(524, 10), 393 => to_unsigned(410, 10), 394 => to_unsigned(454, 10), 395 => to_unsigned(528, 10), 396 => to_unsigned(475, 10), 397 => to_unsigned(455, 10), 398 => to_unsigned(373, 10), 399 => to_unsigned(376, 10), 400 => to_unsigned(662, 10), 401 => to_unsigned(667, 10), 402 => to_unsigned(406, 10), 403 => to_unsigned(625, 10), 404 => to_unsigned(617, 10), 405 => to_unsigned(565, 10), 406 => to_unsigned(531, 10), 407 => to_unsigned(534, 10), 408 => to_unsigned(438, 10), 409 => to_unsigned(531, 10), 410 => to_unsigned(563, 10), 411 => to_unsigned(342, 10), 412 => to_unsigned(395, 10), 413 => to_unsigned(519, 10), 414 => to_unsigned(417, 10), 415 => to_unsigned(525, 10), 416 => to_unsigned(358, 10), 417 => to_unsigned(527, 10), 418 => to_unsigned(494, 10), 419 => to_unsigned(363, 10), 420 => to_unsigned(591, 10), 421 => to_unsigned(440, 10), 422 => to_unsigned(408, 10), 423 => to_unsigned(468, 10), 424 => to_unsigned(534, 10), 425 => to_unsigned(519, 10), 426 => to_unsigned(584, 10), 427 => to_unsigned(539, 10), 428 => to_unsigned(488, 10), 429 => to_unsigned(706, 10), 430 => to_unsigned(420, 10), 431 => to_unsigned(317, 10), 432 => to_unsigned(558, 10), 433 => to_unsigned(399, 10), 434 => to_unsigned(574, 10), 435 => to_unsigned(562, 10), 436 => to_unsigned(438, 10), 437 => to_unsigned(552, 10), 438 => to_unsigned(550, 10), 439 => to_unsigned(413, 10), 440 => to_unsigned(521, 10), 441 => to_unsigned(537, 10), 442 => to_unsigned(548, 10), 443 => to_unsigned(476, 10), 444 => to_unsigned(527, 10), 445 => to_unsigned(422, 10), 446 => to_unsigned(359, 10), 447 => to_unsigned(610, 10), 448 => to_unsigned(699, 10), 449 => to_unsigned(431, 10), 450 => to_unsigned(522, 10), 451 => to_unsigned(417, 10), 452 => to_unsigned(560, 10), 453 => to_unsigned(442, 10), 454 => to_unsigned(452, 10), 455 => to_unsigned(471, 10), 456 => to_unsigned(337, 10), 457 => to_unsigned(435, 10), 458 => to_unsigned(403, 10), 459 => to_unsigned(726, 10), 460 => to_unsigned(629, 10), 461 => to_unsigned(480, 10), 462 => to_unsigned(572, 10), 463 => to_unsigned(463, 10), 464 => to_unsigned(598, 10), 465 => to_unsigned(650, 10), 466 => to_unsigned(323, 10), 467 => to_unsigned(590, 10), 468 => to_unsigned(394, 10), 469 => to_unsigned(467, 10), 470 => to_unsigned(528, 10), 471 => to_unsigned(491, 10), 472 => to_unsigned(388, 10), 473 => to_unsigned(473, 10), 474 => to_unsigned(594, 10), 475 => to_unsigned(567, 10), 476 => to_unsigned(628, 10), 477 => to_unsigned(667, 10), 478 => to_unsigned(491, 10), 479 => to_unsigned(386, 10), 480 => to_unsigned(579, 10), 481 => to_unsigned(369, 10), 482 => to_unsigned(514, 10), 483 => to_unsigned(475, 10), 484 => to_unsigned(571, 10), 485 => to_unsigned(652, 10), 486 => to_unsigned(488, 10), 487 => to_unsigned(619, 10), 488 => to_unsigned(552, 10), 489 => to_unsigned(467, 10), 490 => to_unsigned(612, 10), 491 => to_unsigned(486, 10), 492 => to_unsigned(571, 10), 493 => to_unsigned(593, 10), 494 => to_unsigned(396, 10), 495 => to_unsigned(370, 10), 496 => to_unsigned(479, 10), 497 => to_unsigned(616, 10), 498 => to_unsigned(605, 10), 499 => to_unsigned(449, 10), 500 => to_unsigned(425, 10), 501 => to_unsigned(411, 10), 502 => to_unsigned(585, 10), 503 => to_unsigned(452, 10), 504 => to_unsigned(519, 10), 505 => to_unsigned(496, 10), 506 => to_unsigned(743, 10), 507 => to_unsigned(636, 10), 508 => to_unsigned(676, 10), 509 => to_unsigned(429, 10), 510 => to_unsigned(558, 10), 511 => to_unsigned(561, 10), 512 => to_unsigned(606, 10), 513 => to_unsigned(627, 10), 514 => to_unsigned(602, 10), 515 => to_unsigned(507, 10), 516 => to_unsigned(420, 10), 517 => to_unsigned(486, 10), 518 => to_unsigned(429, 10), 519 => to_unsigned(620, 10), 520 => to_unsigned(474, 10), 521 => to_unsigned(529, 10), 522 => to_unsigned(443, 10), 523 => to_unsigned(498, 10), 524 => to_unsigned(537, 10), 525 => to_unsigned(530, 10), 526 => to_unsigned(386, 10), 527 => to_unsigned(623, 10), 528 => to_unsigned(575, 10), 529 => to_unsigned(515, 10), 530 => to_unsigned(442, 10), 531 => to_unsigned(744, 10), 532 => to_unsigned(567, 10), 533 => to_unsigned(552, 10), 534 => to_unsigned(473, 10), 535 => to_unsigned(411, 10), 536 => to_unsigned(375, 10), 537 => to_unsigned(619, 10), 538 => to_unsigned(515, 10), 539 => to_unsigned(585, 10), 540 => to_unsigned(374, 10), 541 => to_unsigned(288, 10), 542 => to_unsigned(616, 10), 543 => to_unsigned(397, 10), 544 => to_unsigned(525, 10), 545 => to_unsigned(579, 10), 546 => to_unsigned(766, 10), 547 => to_unsigned(571, 10), 548 => to_unsigned(462, 10), 549 => to_unsigned(478, 10), 550 => to_unsigned(436, 10), 551 => to_unsigned(630, 10), 552 => to_unsigned(320, 10), 553 => to_unsigned(482, 10), 554 => to_unsigned(659, 10), 555 => to_unsigned(486, 10), 556 => to_unsigned(526, 10), 557 => to_unsigned(521, 10), 558 => to_unsigned(434, 10), 559 => to_unsigned(514, 10), 560 => to_unsigned(485, 10), 561 => to_unsigned(485, 10), 562 => to_unsigned(478, 10), 563 => to_unsigned(478, 10), 564 => to_unsigned(470, 10), 565 => to_unsigned(456, 10), 566 => to_unsigned(530, 10), 567 => to_unsigned(507, 10), 568 => to_unsigned(415, 10), 569 => to_unsigned(575, 10), 570 => to_unsigned(524, 10), 571 => to_unsigned(575, 10), 572 => to_unsigned(370, 10), 573 => to_unsigned(422, 10), 574 => to_unsigned(508, 10), 575 => to_unsigned(437, 10), 576 => to_unsigned(356, 10), 577 => to_unsigned(569, 10), 578 => to_unsigned(575, 10), 579 => to_unsigned(480, 10), 580 => to_unsigned(547, 10), 581 => to_unsigned(371, 10), 582 => to_unsigned(416, 10), 583 => to_unsigned(616, 10), 584 => to_unsigned(364, 10), 585 => to_unsigned(567, 10), 586 => to_unsigned(575, 10), 587 => to_unsigned(562, 10), 588 => to_unsigned(546, 10), 589 => to_unsigned(649, 10), 590 => to_unsigned(402, 10), 591 => to_unsigned(534, 10), 592 => to_unsigned(472, 10), 593 => to_unsigned(514, 10), 594 => to_unsigned(688, 10), 595 => to_unsigned(568, 10), 596 => to_unsigned(468, 10), 597 => to_unsigned(349, 10), 598 => to_unsigned(498, 10), 599 => to_unsigned(497, 10), 600 => to_unsigned(438, 10), 601 => to_unsigned(649, 10), 602 => to_unsigned(644, 10), 603 => to_unsigned(317, 10), 604 => to_unsigned(657, 10), 605 => to_unsigned(420, 10), 606 => to_unsigned(561, 10), 607 => to_unsigned(492, 10), 608 => to_unsigned(341, 10), 609 => to_unsigned(570, 10), 610 => to_unsigned(482, 10), 611 => to_unsigned(684, 10), 612 => to_unsigned(589, 10), 613 => to_unsigned(547, 10), 614 => to_unsigned(397, 10), 615 => to_unsigned(635, 10), 616 => to_unsigned(595, 10), 617 => to_unsigned(555, 10), 618 => to_unsigned(472, 10), 619 => to_unsigned(499, 10), 620 => to_unsigned(534, 10), 621 => to_unsigned(557, 10), 622 => to_unsigned(537, 10), 623 => to_unsigned(461, 10), 624 => to_unsigned(392, 10), 625 => to_unsigned(589, 10), 626 => to_unsigned(379, 10), 627 => to_unsigned(563, 10), 628 => to_unsigned(450, 10), 629 => to_unsigned(627, 10), 630 => to_unsigned(533, 10), 631 => to_unsigned(629, 10), 632 => to_unsigned(641, 10), 633 => to_unsigned(554, 10), 634 => to_unsigned(658, 10), 635 => to_unsigned(622, 10), 636 => to_unsigned(375, 10), 637 => to_unsigned(664, 10), 638 => to_unsigned(501, 10), 639 => to_unsigned(511, 10), 640 => to_unsigned(547, 10), 641 => to_unsigned(405, 10), 642 => to_unsigned(622, 10), 643 => to_unsigned(592, 10), 644 => to_unsigned(594, 10), 645 => to_unsigned(438, 10), 646 => to_unsigned(553, 10), 647 => to_unsigned(633, 10), 648 => to_unsigned(566, 10), 649 => to_unsigned(563, 10), 650 => to_unsigned(464, 10), 651 => to_unsigned(463, 10), 652 => to_unsigned(387, 10), 653 => to_unsigned(547, 10), 654 => to_unsigned(391, 10), 655 => to_unsigned(355, 10), 656 => to_unsigned(549, 10), 657 => to_unsigned(426, 10), 658 => to_unsigned(561, 10), 659 => to_unsigned(526, 10), 660 => to_unsigned(562, 10), 661 => to_unsigned(472, 10), 662 => to_unsigned(463, 10), 663 => to_unsigned(368, 10), 664 => to_unsigned(416, 10), 665 => to_unsigned(552, 10), 666 => to_unsigned(384, 10), 667 => to_unsigned(381, 10), 668 => to_unsigned(497, 10), 669 => to_unsigned(481, 10), 670 => to_unsigned(538, 10), 671 => to_unsigned(594, 10), 672 => to_unsigned(362, 10), 673 => to_unsigned(671, 10), 674 => to_unsigned(451, 10), 675 => to_unsigned(443, 10), 676 => to_unsigned(517, 10), 677 => to_unsigned(470, 10), 678 => to_unsigned(438, 10), 679 => to_unsigned(476, 10), 680 => to_unsigned(613, 10), 681 => to_unsigned(567, 10), 682 => to_unsigned(445, 10), 683 => to_unsigned(419, 10), 684 => to_unsigned(585, 10), 685 => to_unsigned(507, 10), 686 => to_unsigned(676, 10), 687 => to_unsigned(492, 10), 688 => to_unsigned(490, 10), 689 => to_unsigned(608, 10), 690 => to_unsigned(566, 10), 691 => to_unsigned(475, 10), 692 => to_unsigned(645, 10), 693 => to_unsigned(480, 10), 694 => to_unsigned(540, 10), 695 => to_unsigned(488, 10), 696 => to_unsigned(435, 10), 697 => to_unsigned(383, 10), 698 => to_unsigned(671, 10), 699 => to_unsigned(452, 10), 700 => to_unsigned(406, 10), 701 => to_unsigned(589, 10), 702 => to_unsigned(438, 10), 703 => to_unsigned(484, 10), 704 => to_unsigned(449, 10), 705 => to_unsigned(404, 10), 706 => to_unsigned(653, 10), 707 => to_unsigned(714, 10), 708 => to_unsigned(349, 10), 709 => to_unsigned(521, 10), 710 => to_unsigned(674, 10), 711 => to_unsigned(401, 10), 712 => to_unsigned(437, 10), 713 => to_unsigned(467, 10), 714 => to_unsigned(508, 10), 715 => to_unsigned(473, 10), 716 => to_unsigned(743, 10), 717 => to_unsigned(590, 10), 718 => to_unsigned(606, 10), 719 => to_unsigned(507, 10), 720 => to_unsigned(557, 10), 721 => to_unsigned(643, 10), 722 => to_unsigned(614, 10), 723 => to_unsigned(721, 10), 724 => to_unsigned(487, 10), 725 => to_unsigned(472, 10), 726 => to_unsigned(636, 10), 727 => to_unsigned(407, 10), 728 => to_unsigned(484, 10), 729 => to_unsigned(603, 10), 730 => to_unsigned(643, 10), 731 => to_unsigned(522, 10), 732 => to_unsigned(545, 10), 733 => to_unsigned(362, 10), 734 => to_unsigned(488, 10), 735 => to_unsigned(630, 10), 736 => to_unsigned(511, 10), 737 => to_unsigned(438, 10), 738 => to_unsigned(559, 10), 739 => to_unsigned(342, 10), 740 => to_unsigned(504, 10), 741 => to_unsigned(645, 10), 742 => to_unsigned(682, 10), 743 => to_unsigned(541, 10), 744 => to_unsigned(570, 10), 745 => to_unsigned(485, 10), 746 => to_unsigned(544, 10), 747 => to_unsigned(530, 10), 748 => to_unsigned(546, 10), 749 => to_unsigned(629, 10), 750 => to_unsigned(441, 10), 751 => to_unsigned(496, 10), 752 => to_unsigned(550, 10), 753 => to_unsigned(490, 10), 754 => to_unsigned(548, 10), 755 => to_unsigned(588, 10), 756 => to_unsigned(428, 10), 757 => to_unsigned(519, 10), 758 => to_unsigned(445, 10), 759 => to_unsigned(348, 10), 760 => to_unsigned(524, 10), 761 => to_unsigned(719, 10), 762 => to_unsigned(398, 10), 763 => to_unsigned(516, 10), 764 => to_unsigned(571, 10), 765 => to_unsigned(497, 10), 766 => to_unsigned(528, 10), 767 => to_unsigned(497, 10), 768 => to_unsigned(343, 10), 769 => to_unsigned(535, 10), 770 => to_unsigned(432, 10), 771 => to_unsigned(521, 10), 772 => to_unsigned(519, 10), 773 => to_unsigned(381, 10), 774 => to_unsigned(621, 10), 775 => to_unsigned(462, 10), 776 => to_unsigned(718, 10), 777 => to_unsigned(586, 10), 778 => to_unsigned(598, 10), 779 => to_unsigned(545, 10), 780 => to_unsigned(477, 10), 781 => to_unsigned(576, 10), 782 => to_unsigned(588, 10), 783 => to_unsigned(559, 10), 784 => to_unsigned(373, 10), 785 => to_unsigned(490, 10), 786 => to_unsigned(462, 10), 787 => to_unsigned(541, 10), 788 => to_unsigned(640, 10), 789 => to_unsigned(548, 10), 790 => to_unsigned(717, 10), 791 => to_unsigned(650, 10), 792 => to_unsigned(325, 10), 793 => to_unsigned(428, 10), 794 => to_unsigned(459, 10), 795 => to_unsigned(575, 10), 796 => to_unsigned(486, 10), 797 => to_unsigned(546, 10), 798 => to_unsigned(713, 10), 799 => to_unsigned(651, 10), 800 => to_unsigned(522, 10), 801 => to_unsigned(491, 10), 802 => to_unsigned(565, 10), 803 => to_unsigned(580, 10), 804 => to_unsigned(557, 10), 805 => to_unsigned(384, 10), 806 => to_unsigned(501, 10), 807 => to_unsigned(590, 10), 808 => to_unsigned(668, 10), 809 => to_unsigned(530, 10), 810 => to_unsigned(390, 10), 811 => to_unsigned(662, 10), 812 => to_unsigned(571, 10), 813 => to_unsigned(552, 10), 814 => to_unsigned(460, 10), 815 => to_unsigned(523, 10), 816 => to_unsigned(596, 10), 817 => to_unsigned(591, 10), 818 => to_unsigned(501, 10), 819 => to_unsigned(511, 10), 820 => to_unsigned(496, 10), 821 => to_unsigned(313, 10), 822 => to_unsigned(374, 10), 823 => to_unsigned(596, 10), 824 => to_unsigned(659, 10), 825 => to_unsigned(522, 10), 826 => to_unsigned(491, 10), 827 => to_unsigned(230, 10), 828 => to_unsigned(487, 10), 829 => to_unsigned(626, 10), 830 => to_unsigned(463, 10), 831 => to_unsigned(463, 10), 832 => to_unsigned(635, 10), 833 => to_unsigned(558, 10), 834 => to_unsigned(510, 10), 835 => to_unsigned(383, 10), 836 => to_unsigned(531, 10), 837 => to_unsigned(575, 10), 838 => to_unsigned(386, 10), 839 => to_unsigned(568, 10), 840 => to_unsigned(482, 10), 841 => to_unsigned(475, 10), 842 => to_unsigned(444, 10), 843 => to_unsigned(486, 10), 844 => to_unsigned(598, 10), 845 => to_unsigned(704, 10), 846 => to_unsigned(641, 10), 847 => to_unsigned(468, 10), 848 => to_unsigned(278, 10), 849 => to_unsigned(559, 10), 850 => to_unsigned(591, 10), 851 => to_unsigned(353, 10), 852 => to_unsigned(595, 10), 853 => to_unsigned(559, 10), 854 => to_unsigned(506, 10), 855 => to_unsigned(431, 10), 856 => to_unsigned(519, 10), 857 => to_unsigned(432, 10), 858 => to_unsigned(668, 10), 859 => to_unsigned(424, 10), 860 => to_unsigned(400, 10), 861 => to_unsigned(524, 10), 862 => to_unsigned(421, 10), 863 => to_unsigned(512, 10), 864 => to_unsigned(648, 10), 865 => to_unsigned(520, 10), 866 => to_unsigned(373, 10), 867 => to_unsigned(588, 10), 868 => to_unsigned(463, 10), 869 => to_unsigned(477, 10), 870 => to_unsigned(662, 10), 871 => to_unsigned(444, 10), 872 => to_unsigned(409, 10), 873 => to_unsigned(540, 10), 874 => to_unsigned(439, 10), 875 => to_unsigned(454, 10), 876 => to_unsigned(464, 10), 877 => to_unsigned(533, 10), 878 => to_unsigned(505, 10), 879 => to_unsigned(449, 10), 880 => to_unsigned(562, 10), 881 => to_unsigned(460, 10), 882 => to_unsigned(449, 10), 883 => to_unsigned(495, 10), 884 => to_unsigned(411, 10), 885 => to_unsigned(358, 10), 886 => to_unsigned(405, 10), 887 => to_unsigned(325, 10), 888 => to_unsigned(667, 10), 889 => to_unsigned(604, 10), 890 => to_unsigned(539, 10), 891 => to_unsigned(571, 10), 892 => to_unsigned(584, 10), 893 => to_unsigned(507, 10), 894 => to_unsigned(499, 10), 895 => to_unsigned(539, 10), 896 => to_unsigned(484, 10), 897 => to_unsigned(422, 10), 898 => to_unsigned(504, 10), 899 => to_unsigned(517, 10), 900 => to_unsigned(671, 10), 901 => to_unsigned(347, 10), 902 => to_unsigned(286, 10), 903 => to_unsigned(665, 10), 904 => to_unsigned(530, 10), 905 => to_unsigned(477, 10), 906 => to_unsigned(466, 10), 907 => to_unsigned(375, 10), 908 => to_unsigned(402, 10), 909 => to_unsigned(412, 10), 910 => to_unsigned(487, 10), 911 => to_unsigned(568, 10), 912 => to_unsigned(388, 10), 913 => to_unsigned(373, 10), 914 => to_unsigned(449, 10), 915 => to_unsigned(479, 10), 916 => to_unsigned(571, 10), 917 => to_unsigned(425, 10), 918 => to_unsigned(374, 10), 919 => to_unsigned(559, 10), 920 => to_unsigned(516, 10), 921 => to_unsigned(407, 10), 922 => to_unsigned(441, 10), 923 => to_unsigned(560, 10), 924 => to_unsigned(611, 10), 925 => to_unsigned(496, 10), 926 => to_unsigned(459, 10), 927 => to_unsigned(440, 10), 928 => to_unsigned(488, 10), 929 => to_unsigned(390, 10), 930 => to_unsigned(616, 10), 931 => to_unsigned(625, 10), 932 => to_unsigned(629, 10), 933 => to_unsigned(430, 10), 934 => to_unsigned(507, 10), 935 => to_unsigned(490, 10), 936 => to_unsigned(554, 10), 937 => to_unsigned(570, 10), 938 => to_unsigned(534, 10), 939 => to_unsigned(520, 10), 940 => to_unsigned(730, 10), 941 => to_unsigned(572, 10), 942 => to_unsigned(321, 10), 943 => to_unsigned(514, 10), 944 => to_unsigned(513, 10), 945 => to_unsigned(612, 10), 946 => to_unsigned(594, 10), 947 => to_unsigned(519, 10), 948 => to_unsigned(559, 10), 949 => to_unsigned(575, 10), 950 => to_unsigned(559, 10), 951 => to_unsigned(577, 10), 952 => to_unsigned(556, 10), 953 => to_unsigned(648, 10), 954 => to_unsigned(328, 10), 955 => to_unsigned(438, 10), 956 => to_unsigned(476, 10), 957 => to_unsigned(637, 10), 958 => to_unsigned(458, 10), 959 => to_unsigned(273, 10), 960 => to_unsigned(689, 10), 961 => to_unsigned(532, 10), 962 => to_unsigned(751, 10), 963 => to_unsigned(392, 10), 964 => to_unsigned(534, 10), 965 => to_unsigned(475, 10), 966 => to_unsigned(484, 10), 967 => to_unsigned(543, 10), 968 => to_unsigned(528, 10), 969 => to_unsigned(381, 10), 970 => to_unsigned(557, 10), 971 => to_unsigned(574, 10), 972 => to_unsigned(493, 10), 973 => to_unsigned(466, 10), 974 => to_unsigned(515, 10), 975 => to_unsigned(412, 10), 976 => to_unsigned(530, 10), 977 => to_unsigned(547, 10), 978 => to_unsigned(412, 10), 979 => to_unsigned(392, 10), 980 => to_unsigned(355, 10), 981 => to_unsigned(439, 10), 982 => to_unsigned(589, 10), 983 => to_unsigned(558, 10), 984 => to_unsigned(493, 10), 985 => to_unsigned(681, 10), 986 => to_unsigned(414, 10), 987 => to_unsigned(489, 10), 988 => to_unsigned(410, 10), 989 => to_unsigned(644, 10), 990 => to_unsigned(430, 10), 991 => to_unsigned(576, 10), 992 => to_unsigned(557, 10), 993 => to_unsigned(425, 10), 994 => to_unsigned(573, 10), 995 => to_unsigned(455, 10), 996 => to_unsigned(575, 10), 997 => to_unsigned(435, 10), 998 => to_unsigned(565, 10), 999 => to_unsigned(604, 10), 1000 => to_unsigned(620, 10), 1001 => to_unsigned(426, 10), 1002 => to_unsigned(438, 10), 1003 => to_unsigned(483, 10), 1004 => to_unsigned(515, 10), 1005 => to_unsigned(326, 10), 1006 => to_unsigned(593, 10), 1007 => to_unsigned(550, 10), 1008 => to_unsigned(554, 10), 1009 => to_unsigned(573, 10), 1010 => to_unsigned(603, 10), 1011 => to_unsigned(433, 10), 1012 => to_unsigned(504, 10), 1013 => to_unsigned(619, 10), 1014 => to_unsigned(264, 10), 1015 => to_unsigned(561, 10), 1016 => to_unsigned(467, 10), 1017 => to_unsigned(582, 10), 1018 => to_unsigned(326, 10), 1019 => to_unsigned(519, 10), 1020 => to_unsigned(436, 10), 1021 => to_unsigned(486, 10), 1022 => to_unsigned(465, 10), 1023 => to_unsigned(545, 10), 1024 => to_unsigned(519, 10), 1025 => to_unsigned(508, 10), 1026 => to_unsigned(444, 10), 1027 => to_unsigned(540, 10), 1028 => to_unsigned(334, 10), 1029 => to_unsigned(538, 10), 1030 => to_unsigned(605, 10), 1031 => to_unsigned(585, 10), 1032 => to_unsigned(672, 10), 1033 => to_unsigned(455, 10), 1034 => to_unsigned(538, 10), 1035 => to_unsigned(521, 10), 1036 => to_unsigned(408, 10), 1037 => to_unsigned(468, 10), 1038 => to_unsigned(575, 10), 1039 => to_unsigned(547, 10), 1040 => to_unsigned(633, 10), 1041 => to_unsigned(441, 10), 1042 => to_unsigned(350, 10), 1043 => to_unsigned(540, 10), 1044 => to_unsigned(532, 10), 1045 => to_unsigned(646, 10), 1046 => to_unsigned(694, 10), 1047 => to_unsigned(491, 10), 1048 => to_unsigned(524, 10), 1049 => to_unsigned(551, 10), 1050 => to_unsigned(403, 10), 1051 => to_unsigned(482, 10), 1052 => to_unsigned(278, 10), 1053 => to_unsigned(515, 10), 1054 => to_unsigned(512, 10), 1055 => to_unsigned(552, 10), 1056 => to_unsigned(529, 10), 1057 => to_unsigned(462, 10), 1058 => to_unsigned(514, 10), 1059 => to_unsigned(602, 10), 1060 => to_unsigned(618, 10), 1061 => to_unsigned(408, 10), 1062 => to_unsigned(480, 10), 1063 => to_unsigned(621, 10), 1064 => to_unsigned(461, 10), 1065 => to_unsigned(590, 10), 1066 => to_unsigned(416, 10), 1067 => to_unsigned(505, 10), 1068 => to_unsigned(381, 10), 1069 => to_unsigned(499, 10), 1070 => to_unsigned(558, 10), 1071 => to_unsigned(601, 10), 1072 => to_unsigned(402, 10), 1073 => to_unsigned(566, 10), 1074 => to_unsigned(562, 10), 1075 => to_unsigned(581, 10), 1076 => to_unsigned(521, 10), 1077 => to_unsigned(406, 10), 1078 => to_unsigned(521, 10), 1079 => to_unsigned(463, 10), 1080 => to_unsigned(574, 10), 1081 => to_unsigned(447, 10), 1082 => to_unsigned(603, 10), 1083 => to_unsigned(494, 10), 1084 => to_unsigned(490, 10), 1085 => to_unsigned(420, 10), 1086 => to_unsigned(587, 10), 1087 => to_unsigned(431, 10), 1088 => to_unsigned(549, 10), 1089 => to_unsigned(546, 10), 1090 => to_unsigned(579, 10), 1091 => to_unsigned(491, 10), 1092 => to_unsigned(574, 10), 1093 => to_unsigned(384, 10), 1094 => to_unsigned(550, 10), 1095 => to_unsigned(363, 10), 1096 => to_unsigned(519, 10), 1097 => to_unsigned(557, 10), 1098 => to_unsigned(427, 10), 1099 => to_unsigned(536, 10), 1100 => to_unsigned(344, 10), 1101 => to_unsigned(479, 10), 1102 => to_unsigned(399, 10), 1103 => to_unsigned(374, 10), 1104 => to_unsigned(400, 10), 1105 => to_unsigned(308, 10), 1106 => to_unsigned(456, 10), 1107 => to_unsigned(392, 10), 1108 => to_unsigned(675, 10), 1109 => to_unsigned(518, 10), 1110 => to_unsigned(465, 10), 1111 => to_unsigned(637, 10), 1112 => to_unsigned(729, 10), 1113 => to_unsigned(664, 10), 1114 => to_unsigned(511, 10), 1115 => to_unsigned(502, 10), 1116 => to_unsigned(546, 10), 1117 => to_unsigned(499, 10), 1118 => to_unsigned(598, 10), 1119 => to_unsigned(444, 10), 1120 => to_unsigned(524, 10), 1121 => to_unsigned(461, 10), 1122 => to_unsigned(581, 10), 1123 => to_unsigned(606, 10), 1124 => to_unsigned(509, 10), 1125 => to_unsigned(535, 10), 1126 => to_unsigned(651, 10), 1127 => to_unsigned(511, 10), 1128 => to_unsigned(524, 10), 1129 => to_unsigned(252, 10), 1130 => to_unsigned(586, 10), 1131 => to_unsigned(620, 10), 1132 => to_unsigned(590, 10), 1133 => to_unsigned(469, 10), 1134 => to_unsigned(501, 10), 1135 => to_unsigned(638, 10), 1136 => to_unsigned(469, 10), 1137 => to_unsigned(528, 10), 1138 => to_unsigned(513, 10), 1139 => to_unsigned(620, 10), 1140 => to_unsigned(503, 10), 1141 => to_unsigned(502, 10), 1142 => to_unsigned(591, 10), 1143 => to_unsigned(381, 10), 1144 => to_unsigned(507, 10), 1145 => to_unsigned(358, 10), 1146 => to_unsigned(504, 10), 1147 => to_unsigned(473, 10), 1148 => to_unsigned(581, 10), 1149 => to_unsigned(545, 10), 1150 => to_unsigned(513, 10), 1151 => to_unsigned(593, 10), 1152 => to_unsigned(621, 10), 1153 => to_unsigned(625, 10), 1154 => to_unsigned(444, 10), 1155 => to_unsigned(457, 10), 1156 => to_unsigned(515, 10), 1157 => to_unsigned(640, 10), 1158 => to_unsigned(488, 10), 1159 => to_unsigned(434, 10), 1160 => to_unsigned(435, 10), 1161 => to_unsigned(472, 10), 1162 => to_unsigned(598, 10), 1163 => to_unsigned(565, 10), 1164 => to_unsigned(487, 10), 1165 => to_unsigned(372, 10), 1166 => to_unsigned(643, 10), 1167 => to_unsigned(354, 10), 1168 => to_unsigned(484, 10), 1169 => to_unsigned(573, 10), 1170 => to_unsigned(582, 10), 1171 => to_unsigned(264, 10), 1172 => to_unsigned(640, 10), 1173 => to_unsigned(545, 10), 1174 => to_unsigned(609, 10), 1175 => to_unsigned(555, 10), 1176 => to_unsigned(578, 10), 1177 => to_unsigned(732, 10), 1178 => to_unsigned(679, 10), 1179 => to_unsigned(397, 10), 1180 => to_unsigned(669, 10), 1181 => to_unsigned(389, 10), 1182 => to_unsigned(485, 10), 1183 => to_unsigned(398, 10), 1184 => to_unsigned(512, 10), 1185 => to_unsigned(367, 10), 1186 => to_unsigned(508, 10), 1187 => to_unsigned(573, 10), 1188 => to_unsigned(409, 10), 1189 => to_unsigned(432, 10), 1190 => to_unsigned(495, 10), 1191 => to_unsigned(637, 10), 1192 => to_unsigned(631, 10), 1193 => to_unsigned(648, 10), 1194 => to_unsigned(561, 10), 1195 => to_unsigned(663, 10), 1196 => to_unsigned(392, 10), 1197 => to_unsigned(607, 10), 1198 => to_unsigned(456, 10), 1199 => to_unsigned(551, 10), 1200 => to_unsigned(461, 10), 1201 => to_unsigned(532, 10), 1202 => to_unsigned(486, 10), 1203 => to_unsigned(588, 10), 1204 => to_unsigned(499, 10), 1205 => to_unsigned(506, 10), 1206 => to_unsigned(422, 10), 1207 => to_unsigned(443, 10), 1208 => to_unsigned(572, 10), 1209 => to_unsigned(388, 10), 1210 => to_unsigned(567, 10), 1211 => to_unsigned(397, 10), 1212 => to_unsigned(525, 10), 1213 => to_unsigned(360, 10), 1214 => to_unsigned(555, 10), 1215 => to_unsigned(541, 10), 1216 => to_unsigned(424, 10), 1217 => to_unsigned(568, 10), 1218 => to_unsigned(412, 10), 1219 => to_unsigned(471, 10), 1220 => to_unsigned(550, 10), 1221 => to_unsigned(545, 10), 1222 => to_unsigned(436, 10), 1223 => to_unsigned(389, 10), 1224 => to_unsigned(669, 10), 1225 => to_unsigned(468, 10), 1226 => to_unsigned(426, 10), 1227 => to_unsigned(465, 10), 1228 => to_unsigned(486, 10), 1229 => to_unsigned(556, 10), 1230 => to_unsigned(708, 10), 1231 => to_unsigned(682, 10), 1232 => to_unsigned(622, 10), 1233 => to_unsigned(512, 10), 1234 => to_unsigned(436, 10), 1235 => to_unsigned(460, 10), 1236 => to_unsigned(553, 10), 1237 => to_unsigned(333, 10), 1238 => to_unsigned(593, 10), 1239 => to_unsigned(590, 10), 1240 => to_unsigned(546, 10), 1241 => to_unsigned(487, 10), 1242 => to_unsigned(451, 10), 1243 => to_unsigned(579, 10), 1244 => to_unsigned(612, 10), 1245 => to_unsigned(594, 10), 1246 => to_unsigned(397, 10), 1247 => to_unsigned(413, 10), 1248 => to_unsigned(480, 10), 1249 => to_unsigned(432, 10), 1250 => to_unsigned(614, 10), 1251 => to_unsigned(417, 10), 1252 => to_unsigned(347, 10), 1253 => to_unsigned(484, 10), 1254 => to_unsigned(474, 10), 1255 => to_unsigned(694, 10), 1256 => to_unsigned(452, 10), 1257 => to_unsigned(571, 10), 1258 => to_unsigned(497, 10), 1259 => to_unsigned(420, 10), 1260 => to_unsigned(631, 10), 1261 => to_unsigned(575, 10), 1262 => to_unsigned(537, 10), 1263 => to_unsigned(383, 10), 1264 => to_unsigned(447, 10), 1265 => to_unsigned(663, 10), 1266 => to_unsigned(651, 10), 1267 => to_unsigned(519, 10), 1268 => to_unsigned(348, 10), 1269 => to_unsigned(523, 10), 1270 => to_unsigned(340, 10), 1271 => to_unsigned(498, 10), 1272 => to_unsigned(452, 10), 1273 => to_unsigned(576, 10), 1274 => to_unsigned(532, 10), 1275 => to_unsigned(399, 10), 1276 => to_unsigned(660, 10), 1277 => to_unsigned(566, 10), 1278 => to_unsigned(405, 10), 1279 => to_unsigned(388, 10), 1280 => to_unsigned(348, 10), 1281 => to_unsigned(536, 10), 1282 => to_unsigned(664, 10), 1283 => to_unsigned(419, 10), 1284 => to_unsigned(426, 10), 1285 => to_unsigned(619, 10), 1286 => to_unsigned(577, 10), 1287 => to_unsigned(605, 10), 1288 => to_unsigned(546, 10), 1289 => to_unsigned(497, 10), 1290 => to_unsigned(481, 10), 1291 => to_unsigned(566, 10), 1292 => to_unsigned(449, 10), 1293 => to_unsigned(424, 10), 1294 => to_unsigned(561, 10), 1295 => to_unsigned(656, 10), 1296 => to_unsigned(668, 10), 1297 => to_unsigned(541, 10), 1298 => to_unsigned(461, 10), 1299 => to_unsigned(477, 10), 1300 => to_unsigned(502, 10), 1301 => to_unsigned(564, 10), 1302 => to_unsigned(651, 10), 1303 => to_unsigned(440, 10), 1304 => to_unsigned(484, 10), 1305 => to_unsigned(513, 10), 1306 => to_unsigned(377, 10), 1307 => to_unsigned(575, 10), 1308 => to_unsigned(541, 10), 1309 => to_unsigned(577, 10), 1310 => to_unsigned(324, 10), 1311 => to_unsigned(578, 10), 1312 => to_unsigned(510, 10), 1313 => to_unsigned(509, 10), 1314 => to_unsigned(406, 10), 1315 => to_unsigned(561, 10), 1316 => to_unsigned(475, 10), 1317 => to_unsigned(485, 10), 1318 => to_unsigned(326, 10), 1319 => to_unsigned(519, 10), 1320 => to_unsigned(353, 10), 1321 => to_unsigned(483, 10), 1322 => to_unsigned(543, 10), 1323 => to_unsigned(574, 10), 1324 => to_unsigned(512, 10), 1325 => to_unsigned(490, 10), 1326 => to_unsigned(530, 10), 1327 => to_unsigned(563, 10), 1328 => to_unsigned(474, 10), 1329 => to_unsigned(556, 10), 1330 => to_unsigned(563, 10), 1331 => to_unsigned(583, 10), 1332 => to_unsigned(577, 10), 1333 => to_unsigned(488, 10), 1334 => to_unsigned(620, 10), 1335 => to_unsigned(685, 10), 1336 => to_unsigned(526, 10), 1337 => to_unsigned(570, 10), 1338 => to_unsigned(396, 10), 1339 => to_unsigned(605, 10), 1340 => to_unsigned(293, 10), 1341 => to_unsigned(448, 10), 1342 => to_unsigned(398, 10), 1343 => to_unsigned(600, 10), 1344 => to_unsigned(422, 10), 1345 => to_unsigned(504, 10), 1346 => to_unsigned(504, 10), 1347 => to_unsigned(636, 10), 1348 => to_unsigned(449, 10), 1349 => to_unsigned(402, 10), 1350 => to_unsigned(593, 10), 1351 => to_unsigned(476, 10), 1352 => to_unsigned(325, 10), 1353 => to_unsigned(606, 10), 1354 => to_unsigned(650, 10), 1355 => to_unsigned(558, 10), 1356 => to_unsigned(417, 10), 1357 => to_unsigned(618, 10), 1358 => to_unsigned(505, 10), 1359 => to_unsigned(647, 10), 1360 => to_unsigned(545, 10), 1361 => to_unsigned(520, 10), 1362 => to_unsigned(477, 10), 1363 => to_unsigned(384, 10), 1364 => to_unsigned(510, 10), 1365 => to_unsigned(336, 10), 1366 => to_unsigned(506, 10), 1367 => to_unsigned(584, 10), 1368 => to_unsigned(521, 10), 1369 => to_unsigned(493, 10), 1370 => to_unsigned(557, 10), 1371 => to_unsigned(443, 10), 1372 => to_unsigned(592, 10), 1373 => to_unsigned(358, 10), 1374 => to_unsigned(591, 10), 1375 => to_unsigned(318, 10), 1376 => to_unsigned(418, 10), 1377 => to_unsigned(433, 10), 1378 => to_unsigned(541, 10), 1379 => to_unsigned(426, 10), 1380 => to_unsigned(580, 10), 1381 => to_unsigned(505, 10), 1382 => to_unsigned(564, 10), 1383 => to_unsigned(569, 10), 1384 => to_unsigned(562, 10), 1385 => to_unsigned(390, 10), 1386 => to_unsigned(573, 10), 1387 => to_unsigned(444, 10), 1388 => to_unsigned(533, 10), 1389 => to_unsigned(462, 10), 1390 => to_unsigned(513, 10), 1391 => to_unsigned(356, 10), 1392 => to_unsigned(519, 10), 1393 => to_unsigned(615, 10), 1394 => to_unsigned(513, 10), 1395 => to_unsigned(472, 10), 1396 => to_unsigned(506, 10), 1397 => to_unsigned(599, 10), 1398 => to_unsigned(405, 10), 1399 => to_unsigned(525, 10), 1400 => to_unsigned(597, 10), 1401 => to_unsigned(420, 10), 1402 => to_unsigned(493, 10), 1403 => to_unsigned(423, 10), 1404 => to_unsigned(348, 10), 1405 => to_unsigned(432, 10), 1406 => to_unsigned(561, 10), 1407 => to_unsigned(588, 10), 1408 => to_unsigned(432, 10), 1409 => to_unsigned(634, 10), 1410 => to_unsigned(287, 10), 1411 => to_unsigned(423, 10), 1412 => to_unsigned(614, 10), 1413 => to_unsigned(427, 10), 1414 => to_unsigned(375, 10), 1415 => to_unsigned(397, 10), 1416 => to_unsigned(439, 10), 1417 => to_unsigned(466, 10), 1418 => to_unsigned(419, 10), 1419 => to_unsigned(469, 10), 1420 => to_unsigned(705, 10), 1421 => to_unsigned(649, 10), 1422 => to_unsigned(514, 10), 1423 => to_unsigned(594, 10), 1424 => to_unsigned(390, 10), 1425 => to_unsigned(564, 10), 1426 => to_unsigned(542, 10), 1427 => to_unsigned(712, 10), 1428 => to_unsigned(384, 10), 1429 => to_unsigned(462, 10), 1430 => to_unsigned(627, 10), 1431 => to_unsigned(539, 10), 1432 => to_unsigned(506, 10), 1433 => to_unsigned(486, 10), 1434 => to_unsigned(537, 10), 1435 => to_unsigned(441, 10), 1436 => to_unsigned(581, 10), 1437 => to_unsigned(555, 10), 1438 => to_unsigned(404, 10), 1439 => to_unsigned(440, 10), 1440 => to_unsigned(531, 10), 1441 => to_unsigned(344, 10), 1442 => to_unsigned(421, 10), 1443 => to_unsigned(588, 10), 1444 => to_unsigned(418, 10), 1445 => to_unsigned(527, 10), 1446 => to_unsigned(292, 10), 1447 => to_unsigned(630, 10), 1448 => to_unsigned(573, 10), 1449 => to_unsigned(589, 10), 1450 => to_unsigned(434, 10), 1451 => to_unsigned(486, 10), 1452 => to_unsigned(547, 10), 1453 => to_unsigned(505, 10), 1454 => to_unsigned(384, 10), 1455 => to_unsigned(559, 10), 1456 => to_unsigned(475, 10), 1457 => to_unsigned(460, 10), 1458 => to_unsigned(565, 10), 1459 => to_unsigned(670, 10), 1460 => to_unsigned(378, 10), 1461 => to_unsigned(515, 10), 1462 => to_unsigned(494, 10), 1463 => to_unsigned(367, 10), 1464 => to_unsigned(625, 10), 1465 => to_unsigned(479, 10), 1466 => to_unsigned(666, 10), 1467 => to_unsigned(553, 10), 1468 => to_unsigned(527, 10), 1469 => to_unsigned(465, 10), 1470 => to_unsigned(493, 10), 1471 => to_unsigned(593, 10), 1472 => to_unsigned(587, 10), 1473 => to_unsigned(619, 10), 1474 => to_unsigned(528, 10), 1475 => to_unsigned(493, 10), 1476 => to_unsigned(475, 10), 1477 => to_unsigned(545, 10), 1478 => to_unsigned(453, 10), 1479 => to_unsigned(383, 10), 1480 => to_unsigned(488, 10), 1481 => to_unsigned(531, 10), 1482 => to_unsigned(485, 10), 1483 => to_unsigned(353, 10), 1484 => to_unsigned(423, 10), 1485 => to_unsigned(456, 10), 1486 => to_unsigned(331, 10), 1487 => to_unsigned(584, 10), 1488 => to_unsigned(581, 10), 1489 => to_unsigned(529, 10), 1490 => to_unsigned(471, 10), 1491 => to_unsigned(498, 10), 1492 => to_unsigned(556, 10), 1493 => to_unsigned(405, 10), 1494 => to_unsigned(382, 10), 1495 => to_unsigned(608, 10), 1496 => to_unsigned(493, 10), 1497 => to_unsigned(467, 10), 1498 => to_unsigned(448, 10), 1499 => to_unsigned(495, 10), 1500 => to_unsigned(459, 10), 1501 => to_unsigned(576, 10), 1502 => to_unsigned(361, 10), 1503 => to_unsigned(635, 10), 1504 => to_unsigned(619, 10), 1505 => to_unsigned(537, 10), 1506 => to_unsigned(463, 10), 1507 => to_unsigned(369, 10), 1508 => to_unsigned(495, 10), 1509 => to_unsigned(407, 10), 1510 => to_unsigned(383, 10), 1511 => to_unsigned(478, 10), 1512 => to_unsigned(500, 10), 1513 => to_unsigned(510, 10), 1514 => to_unsigned(617, 10), 1515 => to_unsigned(539, 10), 1516 => to_unsigned(383, 10), 1517 => to_unsigned(629, 10), 1518 => to_unsigned(479, 10), 1519 => to_unsigned(532, 10), 1520 => to_unsigned(451, 10), 1521 => to_unsigned(405, 10), 1522 => to_unsigned(470, 10), 1523 => to_unsigned(392, 10), 1524 => to_unsigned(608, 10), 1525 => to_unsigned(559, 10), 1526 => to_unsigned(548, 10), 1527 => to_unsigned(564, 10), 1528 => to_unsigned(513, 10), 1529 => to_unsigned(570, 10), 1530 => to_unsigned(580, 10), 1531 => to_unsigned(554, 10), 1532 => to_unsigned(477, 10), 1533 => to_unsigned(409, 10), 1534 => to_unsigned(478, 10), 1535 => to_unsigned(458, 10), 1536 => to_unsigned(622, 10), 1537 => to_unsigned(430, 10), 1538 => to_unsigned(458, 10), 1539 => to_unsigned(622, 10), 1540 => to_unsigned(399, 10), 1541 => to_unsigned(447, 10), 1542 => to_unsigned(672, 10), 1543 => to_unsigned(509, 10), 1544 => to_unsigned(514, 10), 1545 => to_unsigned(456, 10), 1546 => to_unsigned(471, 10), 1547 => to_unsigned(425, 10), 1548 => to_unsigned(264, 10), 1549 => to_unsigned(371, 10), 1550 => to_unsigned(716, 10), 1551 => to_unsigned(430, 10), 1552 => to_unsigned(510, 10), 1553 => to_unsigned(669, 10), 1554 => to_unsigned(536, 10), 1555 => to_unsigned(737, 10), 1556 => to_unsigned(531, 10), 1557 => to_unsigned(321, 10), 1558 => to_unsigned(450, 10), 1559 => to_unsigned(500, 10), 1560 => to_unsigned(398, 10), 1561 => to_unsigned(509, 10), 1562 => to_unsigned(419, 10), 1563 => to_unsigned(350, 10), 1564 => to_unsigned(281, 10), 1565 => to_unsigned(543, 10), 1566 => to_unsigned(576, 10), 1567 => to_unsigned(554, 10), 1568 => to_unsigned(559, 10), 1569 => to_unsigned(551, 10), 1570 => to_unsigned(387, 10), 1571 => to_unsigned(469, 10), 1572 => to_unsigned(540, 10), 1573 => to_unsigned(412, 10), 1574 => to_unsigned(369, 10), 1575 => to_unsigned(669, 10), 1576 => to_unsigned(563, 10), 1577 => to_unsigned(625, 10), 1578 => to_unsigned(594, 10), 1579 => to_unsigned(533, 10), 1580 => to_unsigned(692, 10), 1581 => to_unsigned(470, 10), 1582 => to_unsigned(423, 10), 1583 => to_unsigned(533, 10), 1584 => to_unsigned(443, 10), 1585 => to_unsigned(378, 10), 1586 => to_unsigned(436, 10), 1587 => to_unsigned(565, 10), 1588 => to_unsigned(499, 10), 1589 => to_unsigned(506, 10), 1590 => to_unsigned(513, 10), 1591 => to_unsigned(472, 10), 1592 => to_unsigned(499, 10), 1593 => to_unsigned(464, 10), 1594 => to_unsigned(458, 10), 1595 => to_unsigned(603, 10), 1596 => to_unsigned(468, 10), 1597 => to_unsigned(332, 10), 1598 => to_unsigned(475, 10), 1599 => to_unsigned(323, 10), 1600 => to_unsigned(474, 10), 1601 => to_unsigned(621, 10), 1602 => to_unsigned(449, 10), 1603 => to_unsigned(601, 10), 1604 => to_unsigned(578, 10), 1605 => to_unsigned(523, 10), 1606 => to_unsigned(614, 10), 1607 => to_unsigned(517, 10), 1608 => to_unsigned(487, 10), 1609 => to_unsigned(435, 10), 1610 => to_unsigned(578, 10), 1611 => to_unsigned(551, 10), 1612 => to_unsigned(678, 10), 1613 => to_unsigned(495, 10), 1614 => to_unsigned(402, 10), 1615 => to_unsigned(534, 10), 1616 => to_unsigned(467, 10), 1617 => to_unsigned(510, 10), 1618 => to_unsigned(580, 10), 1619 => to_unsigned(272, 10), 1620 => to_unsigned(323, 10), 1621 => to_unsigned(566, 10), 1622 => to_unsigned(387, 10), 1623 => to_unsigned(489, 10), 1624 => to_unsigned(433, 10), 1625 => to_unsigned(459, 10), 1626 => to_unsigned(536, 10), 1627 => to_unsigned(606, 10), 1628 => to_unsigned(597, 10), 1629 => to_unsigned(454, 10), 1630 => to_unsigned(605, 10), 1631 => to_unsigned(369, 10), 1632 => to_unsigned(529, 10), 1633 => to_unsigned(493, 10), 1634 => to_unsigned(460, 10), 1635 => to_unsigned(594, 10), 1636 => to_unsigned(457, 10), 1637 => to_unsigned(506, 10), 1638 => to_unsigned(364, 10), 1639 => to_unsigned(365, 10), 1640 => to_unsigned(526, 10), 1641 => to_unsigned(585, 10), 1642 => to_unsigned(519, 10), 1643 => to_unsigned(541, 10), 1644 => to_unsigned(554, 10), 1645 => to_unsigned(474, 10), 1646 => to_unsigned(516, 10), 1647 => to_unsigned(614, 10), 1648 => to_unsigned(633, 10), 1649 => to_unsigned(466, 10), 1650 => to_unsigned(555, 10), 1651 => to_unsigned(717, 10), 1652 => to_unsigned(491, 10), 1653 => to_unsigned(591, 10), 1654 => to_unsigned(499, 10), 1655 => to_unsigned(576, 10), 1656 => to_unsigned(624, 10), 1657 => to_unsigned(410, 10), 1658 => to_unsigned(517, 10), 1659 => to_unsigned(536, 10), 1660 => to_unsigned(437, 10), 1661 => to_unsigned(642, 10), 1662 => to_unsigned(527, 10), 1663 => to_unsigned(570, 10), 1664 => to_unsigned(727, 10), 1665 => to_unsigned(571, 10), 1666 => to_unsigned(625, 10), 1667 => to_unsigned(580, 10), 1668 => to_unsigned(742, 10), 1669 => to_unsigned(452, 10), 1670 => to_unsigned(506, 10), 1671 => to_unsigned(475, 10), 1672 => to_unsigned(495, 10), 1673 => to_unsigned(476, 10), 1674 => to_unsigned(419, 10), 1675 => to_unsigned(566, 10), 1676 => to_unsigned(677, 10), 1677 => to_unsigned(443, 10), 1678 => to_unsigned(566, 10), 1679 => to_unsigned(611, 10), 1680 => to_unsigned(522, 10), 1681 => to_unsigned(445, 10), 1682 => to_unsigned(452, 10), 1683 => to_unsigned(494, 10), 1684 => to_unsigned(531, 10), 1685 => to_unsigned(560, 10), 1686 => to_unsigned(659, 10), 1687 => to_unsigned(637, 10), 1688 => to_unsigned(352, 10), 1689 => to_unsigned(566, 10), 1690 => to_unsigned(502, 10), 1691 => to_unsigned(474, 10), 1692 => to_unsigned(500, 10), 1693 => to_unsigned(610, 10), 1694 => to_unsigned(518, 10), 1695 => to_unsigned(588, 10), 1696 => to_unsigned(617, 10), 1697 => to_unsigned(436, 10), 1698 => to_unsigned(527, 10), 1699 => to_unsigned(499, 10), 1700 => to_unsigned(546, 10), 1701 => to_unsigned(285, 10), 1702 => to_unsigned(520, 10), 1703 => to_unsigned(490, 10), 1704 => to_unsigned(442, 10), 1705 => to_unsigned(508, 10), 1706 => to_unsigned(431, 10), 1707 => to_unsigned(503, 10), 1708 => to_unsigned(501, 10), 1709 => to_unsigned(673, 10), 1710 => to_unsigned(433, 10), 1711 => to_unsigned(545, 10), 1712 => to_unsigned(539, 10), 1713 => to_unsigned(497, 10), 1714 => to_unsigned(561, 10), 1715 => to_unsigned(602, 10), 1716 => to_unsigned(720, 10), 1717 => to_unsigned(586, 10), 1718 => to_unsigned(622, 10), 1719 => to_unsigned(631, 10), 1720 => to_unsigned(552, 10), 1721 => to_unsigned(537, 10), 1722 => to_unsigned(554, 10), 1723 => to_unsigned(435, 10), 1724 => to_unsigned(581, 10), 1725 => to_unsigned(517, 10), 1726 => to_unsigned(341, 10), 1727 => to_unsigned(518, 10), 1728 => to_unsigned(553, 10), 1729 => to_unsigned(521, 10), 1730 => to_unsigned(425, 10), 1731 => to_unsigned(554, 10), 1732 => to_unsigned(399, 10), 1733 => to_unsigned(341, 10), 1734 => to_unsigned(487, 10), 1735 => to_unsigned(579, 10), 1736 => to_unsigned(489, 10), 1737 => to_unsigned(505, 10), 1738 => to_unsigned(513, 10), 1739 => to_unsigned(486, 10), 1740 => to_unsigned(336, 10), 1741 => to_unsigned(302, 10), 1742 => to_unsigned(352, 10), 1743 => to_unsigned(637, 10), 1744 => to_unsigned(538, 10), 1745 => to_unsigned(399, 10), 1746 => to_unsigned(460, 10), 1747 => to_unsigned(492, 10), 1748 => to_unsigned(605, 10), 1749 => to_unsigned(348, 10), 1750 => to_unsigned(419, 10), 1751 => to_unsigned(438, 10), 1752 => to_unsigned(432, 10), 1753 => to_unsigned(476, 10), 1754 => to_unsigned(519, 10), 1755 => to_unsigned(471, 10), 1756 => to_unsigned(488, 10), 1757 => to_unsigned(508, 10), 1758 => to_unsigned(561, 10), 1759 => to_unsigned(587, 10), 1760 => to_unsigned(446, 10), 1761 => to_unsigned(638, 10), 1762 => to_unsigned(461, 10), 1763 => to_unsigned(461, 10), 1764 => to_unsigned(528, 10), 1765 => to_unsigned(497, 10), 1766 => to_unsigned(652, 10), 1767 => to_unsigned(505, 10), 1768 => to_unsigned(562, 10), 1769 => to_unsigned(647, 10), 1770 => to_unsigned(510, 10), 1771 => to_unsigned(486, 10), 1772 => to_unsigned(214, 10), 1773 => to_unsigned(482, 10), 1774 => to_unsigned(403, 10), 1775 => to_unsigned(531, 10), 1776 => to_unsigned(611, 10), 1777 => to_unsigned(469, 10), 1778 => to_unsigned(614, 10), 1779 => to_unsigned(469, 10), 1780 => to_unsigned(534, 10), 1781 => to_unsigned(463, 10), 1782 => to_unsigned(528, 10), 1783 => to_unsigned(600, 10), 1784 => to_unsigned(591, 10), 1785 => to_unsigned(553, 10), 1786 => to_unsigned(400, 10), 1787 => to_unsigned(492, 10), 1788 => to_unsigned(453, 10), 1789 => to_unsigned(456, 10), 1790 => to_unsigned(439, 10), 1791 => to_unsigned(469, 10), 1792 => to_unsigned(456, 10), 1793 => to_unsigned(429, 10), 1794 => to_unsigned(435, 10), 1795 => to_unsigned(511, 10), 1796 => to_unsigned(488, 10), 1797 => to_unsigned(344, 10), 1798 => to_unsigned(352, 10), 1799 => to_unsigned(343, 10), 1800 => to_unsigned(471, 10), 1801 => to_unsigned(659, 10), 1802 => to_unsigned(502, 10), 1803 => to_unsigned(539, 10), 1804 => to_unsigned(495, 10), 1805 => to_unsigned(607, 10), 1806 => to_unsigned(536, 10), 1807 => to_unsigned(360, 10), 1808 => to_unsigned(298, 10), 1809 => to_unsigned(486, 10), 1810 => to_unsigned(471, 10), 1811 => to_unsigned(405, 10), 1812 => to_unsigned(455, 10), 1813 => to_unsigned(521, 10), 1814 => to_unsigned(511, 10), 1815 => to_unsigned(484, 10), 1816 => to_unsigned(473, 10), 1817 => to_unsigned(571, 10), 1818 => to_unsigned(400, 10), 1819 => to_unsigned(622, 10), 1820 => to_unsigned(487, 10), 1821 => to_unsigned(488, 10), 1822 => to_unsigned(685, 10), 1823 => to_unsigned(395, 10), 1824 => to_unsigned(454, 10), 1825 => to_unsigned(534, 10), 1826 => to_unsigned(265, 10), 1827 => to_unsigned(510, 10), 1828 => to_unsigned(437, 10), 1829 => to_unsigned(548, 10), 1830 => to_unsigned(613, 10), 1831 => to_unsigned(640, 10), 1832 => to_unsigned(631, 10), 1833 => to_unsigned(599, 10), 1834 => to_unsigned(437, 10), 1835 => to_unsigned(447, 10), 1836 => to_unsigned(366, 10), 1837 => to_unsigned(549, 10), 1838 => to_unsigned(590, 10), 1839 => to_unsigned(388, 10), 1840 => to_unsigned(572, 10), 1841 => to_unsigned(589, 10), 1842 => to_unsigned(528, 10), 1843 => to_unsigned(396, 10), 1844 => to_unsigned(508, 10), 1845 => to_unsigned(586, 10), 1846 => to_unsigned(489, 10), 1847 => to_unsigned(655, 10), 1848 => to_unsigned(712, 10), 1849 => to_unsigned(404, 10), 1850 => to_unsigned(647, 10), 1851 => to_unsigned(550, 10), 1852 => to_unsigned(581, 10), 1853 => to_unsigned(360, 10), 1854 => to_unsigned(497, 10), 1855 => to_unsigned(689, 10), 1856 => to_unsigned(507, 10), 1857 => to_unsigned(544, 10), 1858 => to_unsigned(538, 10), 1859 => to_unsigned(527, 10), 1860 => to_unsigned(548, 10), 1861 => to_unsigned(423, 10), 1862 => to_unsigned(361, 10), 1863 => to_unsigned(590, 10), 1864 => to_unsigned(684, 10), 1865 => to_unsigned(482, 10), 1866 => to_unsigned(470, 10), 1867 => to_unsigned(704, 10), 1868 => to_unsigned(621, 10), 1869 => to_unsigned(565, 10), 1870 => to_unsigned(656, 10), 1871 => to_unsigned(577, 10), 1872 => to_unsigned(525, 10), 1873 => to_unsigned(606, 10), 1874 => to_unsigned(438, 10), 1875 => to_unsigned(552, 10), 1876 => to_unsigned(624, 10), 1877 => to_unsigned(516, 10), 1878 => to_unsigned(498, 10), 1879 => to_unsigned(512, 10), 1880 => to_unsigned(600, 10), 1881 => to_unsigned(582, 10), 1882 => to_unsigned(498, 10), 1883 => to_unsigned(573, 10), 1884 => to_unsigned(417, 10), 1885 => to_unsigned(461, 10), 1886 => to_unsigned(584, 10), 1887 => to_unsigned(433, 10), 1888 => to_unsigned(586, 10), 1889 => to_unsigned(584, 10), 1890 => to_unsigned(547, 10), 1891 => to_unsigned(621, 10), 1892 => to_unsigned(659, 10), 1893 => to_unsigned(527, 10), 1894 => to_unsigned(569, 10), 1895 => to_unsigned(419, 10), 1896 => to_unsigned(558, 10), 1897 => to_unsigned(517, 10), 1898 => to_unsigned(655, 10), 1899 => to_unsigned(523, 10), 1900 => to_unsigned(786, 10), 1901 => to_unsigned(542, 10), 1902 => to_unsigned(386, 10), 1903 => to_unsigned(597, 10), 1904 => to_unsigned(607, 10), 1905 => to_unsigned(519, 10), 1906 => to_unsigned(610, 10), 1907 => to_unsigned(534, 10), 1908 => to_unsigned(433, 10), 1909 => to_unsigned(240, 10), 1910 => to_unsigned(473, 10), 1911 => to_unsigned(694, 10), 1912 => to_unsigned(453, 10), 1913 => to_unsigned(440, 10), 1914 => to_unsigned(581, 10), 1915 => to_unsigned(676, 10), 1916 => to_unsigned(454, 10), 1917 => to_unsigned(467, 10), 1918 => to_unsigned(434, 10), 1919 => to_unsigned(494, 10), 1920 => to_unsigned(378, 10), 1921 => to_unsigned(552, 10), 1922 => to_unsigned(673, 10), 1923 => to_unsigned(368, 10), 1924 => to_unsigned(547, 10), 1925 => to_unsigned(552, 10), 1926 => to_unsigned(465, 10), 1927 => to_unsigned(529, 10), 1928 => to_unsigned(457, 10), 1929 => to_unsigned(691, 10), 1930 => to_unsigned(486, 10), 1931 => to_unsigned(426, 10), 1932 => to_unsigned(523, 10), 1933 => to_unsigned(412, 10), 1934 => to_unsigned(472, 10), 1935 => to_unsigned(327, 10), 1936 => to_unsigned(530, 10), 1937 => to_unsigned(449, 10), 1938 => to_unsigned(467, 10), 1939 => to_unsigned(600, 10), 1940 => to_unsigned(341, 10), 1941 => to_unsigned(459, 10), 1942 => to_unsigned(486, 10), 1943 => to_unsigned(417, 10), 1944 => to_unsigned(546, 10), 1945 => to_unsigned(549, 10), 1946 => to_unsigned(730, 10), 1947 => to_unsigned(529, 10), 1948 => to_unsigned(685, 10), 1949 => to_unsigned(419, 10), 1950 => to_unsigned(379, 10), 1951 => to_unsigned(625, 10), 1952 => to_unsigned(551, 10), 1953 => to_unsigned(546, 10), 1954 => to_unsigned(445, 10), 1955 => to_unsigned(586, 10), 1956 => to_unsigned(516, 10), 1957 => to_unsigned(608, 10), 1958 => to_unsigned(478, 10), 1959 => to_unsigned(479, 10), 1960 => to_unsigned(477, 10), 1961 => to_unsigned(412, 10), 1962 => to_unsigned(496, 10), 1963 => to_unsigned(534, 10), 1964 => to_unsigned(393, 10), 1965 => to_unsigned(556, 10), 1966 => to_unsigned(563, 10), 1967 => to_unsigned(643, 10), 1968 => to_unsigned(577, 10), 1969 => to_unsigned(647, 10), 1970 => to_unsigned(409, 10), 1971 => to_unsigned(545, 10), 1972 => to_unsigned(338, 10), 1973 => to_unsigned(604, 10), 1974 => to_unsigned(491, 10), 1975 => to_unsigned(597, 10), 1976 => to_unsigned(449, 10), 1977 => to_unsigned(512, 10), 1978 => to_unsigned(668, 10), 1979 => to_unsigned(635, 10), 1980 => to_unsigned(572, 10), 1981 => to_unsigned(339, 10), 1982 => to_unsigned(540, 10), 1983 => to_unsigned(608, 10), 1984 => to_unsigned(525, 10), 1985 => to_unsigned(612, 10), 1986 => to_unsigned(483, 10), 1987 => to_unsigned(509, 10), 1988 => to_unsigned(578, 10), 1989 => to_unsigned(555, 10), 1990 => to_unsigned(538, 10), 1991 => to_unsigned(444, 10), 1992 => to_unsigned(622, 10), 1993 => to_unsigned(479, 10), 1994 => to_unsigned(513, 10), 1995 => to_unsigned(542, 10), 1996 => to_unsigned(548, 10), 1997 => to_unsigned(653, 10), 1998 => to_unsigned(427, 10), 1999 => to_unsigned(557, 10), 2000 => to_unsigned(663, 10), 2001 => to_unsigned(572, 10), 2002 => to_unsigned(530, 10), 2003 => to_unsigned(497, 10), 2004 => to_unsigned(289, 10), 2005 => to_unsigned(440, 10), 2006 => to_unsigned(596, 10), 2007 => to_unsigned(283, 10), 2008 => to_unsigned(659, 10), 2009 => to_unsigned(509, 10), 2010 => to_unsigned(509, 10), 2011 => to_unsigned(466, 10), 2012 => to_unsigned(641, 10), 2013 => to_unsigned(555, 10), 2014 => to_unsigned(553, 10), 2015 => to_unsigned(497, 10), 2016 => to_unsigned(628, 10), 2017 => to_unsigned(389, 10), 2018 => to_unsigned(465, 10), 2019 => to_unsigned(727, 10), 2020 => to_unsigned(578, 10), 2021 => to_unsigned(340, 10), 2022 => to_unsigned(361, 10), 2023 => to_unsigned(434, 10), 2024 => to_unsigned(572, 10), 2025 => to_unsigned(446, 10), 2026 => to_unsigned(511, 10), 2027 => to_unsigned(361, 10), 2028 => to_unsigned(450, 10), 2029 => to_unsigned(616, 10), 2030 => to_unsigned(560, 10), 2031 => to_unsigned(402, 10), 2032 => to_unsigned(639, 10), 2033 => to_unsigned(544, 10), 2034 => to_unsigned(458, 10), 2035 => to_unsigned(553, 10), 2036 => to_unsigned(516, 10), 2037 => to_unsigned(319, 10), 2038 => to_unsigned(489, 10), 2039 => to_unsigned(342, 10), 2040 => to_unsigned(614, 10), 2041 => to_unsigned(552, 10), 2042 => to_unsigned(597, 10), 2043 => to_unsigned(676, 10), 2044 => to_unsigned(538, 10), 2045 => to_unsigned(636, 10), 2046 => to_unsigned(513, 10), 2047 => to_unsigned(666, 10)),
        2 => (0 => to_unsigned(390, 10), 1 => to_unsigned(470, 10), 2 => to_unsigned(513, 10), 3 => to_unsigned(447, 10), 4 => to_unsigned(461, 10), 5 => to_unsigned(568, 10), 6 => to_unsigned(593, 10), 7 => to_unsigned(492, 10), 8 => to_unsigned(502, 10), 9 => to_unsigned(404, 10), 10 => to_unsigned(528, 10), 11 => to_unsigned(694, 10), 12 => to_unsigned(625, 10), 13 => to_unsigned(634, 10), 14 => to_unsigned(485, 10), 15 => to_unsigned(557, 10), 16 => to_unsigned(479, 10), 17 => to_unsigned(421, 10), 18 => to_unsigned(511, 10), 19 => to_unsigned(564, 10), 20 => to_unsigned(441, 10), 21 => to_unsigned(415, 10), 22 => to_unsigned(461, 10), 23 => to_unsigned(465, 10), 24 => to_unsigned(437, 10), 25 => to_unsigned(538, 10), 26 => to_unsigned(527, 10), 27 => to_unsigned(580, 10), 28 => to_unsigned(709, 10), 29 => to_unsigned(595, 10), 30 => to_unsigned(553, 10), 31 => to_unsigned(583, 10), 32 => to_unsigned(528, 10), 33 => to_unsigned(370, 10), 34 => to_unsigned(651, 10), 35 => to_unsigned(362, 10), 36 => to_unsigned(544, 10), 37 => to_unsigned(452, 10), 38 => to_unsigned(542, 10), 39 => to_unsigned(453, 10), 40 => to_unsigned(663, 10), 41 => to_unsigned(466, 10), 42 => to_unsigned(427, 10), 43 => to_unsigned(308, 10), 44 => to_unsigned(476, 10), 45 => to_unsigned(516, 10), 46 => to_unsigned(572, 10), 47 => to_unsigned(509, 10), 48 => to_unsigned(528, 10), 49 => to_unsigned(519, 10), 50 => to_unsigned(498, 10), 51 => to_unsigned(471, 10), 52 => to_unsigned(586, 10), 53 => to_unsigned(417, 10), 54 => to_unsigned(556, 10), 55 => to_unsigned(534, 10), 56 => to_unsigned(485, 10), 57 => to_unsigned(552, 10), 58 => to_unsigned(517, 10), 59 => to_unsigned(643, 10), 60 => to_unsigned(502, 10), 61 => to_unsigned(500, 10), 62 => to_unsigned(492, 10), 63 => to_unsigned(456, 10), 64 => to_unsigned(482, 10), 65 => to_unsigned(550, 10), 66 => to_unsigned(540, 10), 67 => to_unsigned(546, 10), 68 => to_unsigned(586, 10), 69 => to_unsigned(483, 10), 70 => to_unsigned(502, 10), 71 => to_unsigned(569, 10), 72 => to_unsigned(479, 10), 73 => to_unsigned(425, 10), 74 => to_unsigned(474, 10), 75 => to_unsigned(336, 10), 76 => to_unsigned(560, 10), 77 => to_unsigned(562, 10), 78 => to_unsigned(480, 10), 79 => to_unsigned(437, 10), 80 => to_unsigned(316, 10), 81 => to_unsigned(565, 10), 82 => to_unsigned(372, 10), 83 => to_unsigned(588, 10), 84 => to_unsigned(575, 10), 85 => to_unsigned(494, 10), 86 => to_unsigned(596, 10), 87 => to_unsigned(627, 10), 88 => to_unsigned(443, 10), 89 => to_unsigned(464, 10), 90 => to_unsigned(511, 10), 91 => to_unsigned(545, 10), 92 => to_unsigned(637, 10), 93 => to_unsigned(544, 10), 94 => to_unsigned(339, 10), 95 => to_unsigned(274, 10), 96 => to_unsigned(639, 10), 97 => to_unsigned(663, 10), 98 => to_unsigned(670, 10), 99 => to_unsigned(600, 10), 100 => to_unsigned(348, 10), 101 => to_unsigned(506, 10), 102 => to_unsigned(320, 10), 103 => to_unsigned(386, 10), 104 => to_unsigned(579, 10), 105 => to_unsigned(521, 10), 106 => to_unsigned(455, 10), 107 => to_unsigned(501, 10), 108 => to_unsigned(372, 10), 109 => to_unsigned(594, 10), 110 => to_unsigned(540, 10), 111 => to_unsigned(495, 10), 112 => to_unsigned(548, 10), 113 => to_unsigned(565, 10), 114 => to_unsigned(438, 10), 115 => to_unsigned(417, 10), 116 => to_unsigned(538, 10), 117 => to_unsigned(638, 10), 118 => to_unsigned(484, 10), 119 => to_unsigned(611, 10), 120 => to_unsigned(302, 10), 121 => to_unsigned(606, 10), 122 => to_unsigned(667, 10), 123 => to_unsigned(539, 10), 124 => to_unsigned(635, 10), 125 => to_unsigned(521, 10), 126 => to_unsigned(505, 10), 127 => to_unsigned(407, 10), 128 => to_unsigned(538, 10), 129 => to_unsigned(599, 10), 130 => to_unsigned(581, 10), 131 => to_unsigned(617, 10), 132 => to_unsigned(598, 10), 133 => to_unsigned(565, 10), 134 => to_unsigned(351, 10), 135 => to_unsigned(532, 10), 136 => to_unsigned(446, 10), 137 => to_unsigned(425, 10), 138 => to_unsigned(446, 10), 139 => to_unsigned(540, 10), 140 => to_unsigned(457, 10), 141 => to_unsigned(530, 10), 142 => to_unsigned(483, 10), 143 => to_unsigned(483, 10), 144 => to_unsigned(610, 10), 145 => to_unsigned(478, 10), 146 => to_unsigned(645, 10), 147 => to_unsigned(645, 10), 148 => to_unsigned(431, 10), 149 => to_unsigned(567, 10), 150 => to_unsigned(335, 10), 151 => to_unsigned(459, 10), 152 => to_unsigned(540, 10), 153 => to_unsigned(533, 10), 154 => to_unsigned(429, 10), 155 => to_unsigned(276, 10), 156 => to_unsigned(651, 10), 157 => to_unsigned(523, 10), 158 => to_unsigned(603, 10), 159 => to_unsigned(556, 10), 160 => to_unsigned(536, 10), 161 => to_unsigned(506, 10), 162 => to_unsigned(226, 10), 163 => to_unsigned(458, 10), 164 => to_unsigned(466, 10), 165 => to_unsigned(471, 10), 166 => to_unsigned(456, 10), 167 => to_unsigned(366, 10), 168 => to_unsigned(534, 10), 169 => to_unsigned(335, 10), 170 => to_unsigned(348, 10), 171 => to_unsigned(373, 10), 172 => to_unsigned(543, 10), 173 => to_unsigned(453, 10), 174 => to_unsigned(417, 10), 175 => to_unsigned(661, 10), 176 => to_unsigned(575, 10), 177 => to_unsigned(510, 10), 178 => to_unsigned(516, 10), 179 => to_unsigned(635, 10), 180 => to_unsigned(507, 10), 181 => to_unsigned(636, 10), 182 => to_unsigned(639, 10), 183 => to_unsigned(482, 10), 184 => to_unsigned(567, 10), 185 => to_unsigned(602, 10), 186 => to_unsigned(448, 10), 187 => to_unsigned(550, 10), 188 => to_unsigned(382, 10), 189 => to_unsigned(583, 10), 190 => to_unsigned(436, 10), 191 => to_unsigned(697, 10), 192 => to_unsigned(567, 10), 193 => to_unsigned(617, 10), 194 => to_unsigned(381, 10), 195 => to_unsigned(426, 10), 196 => to_unsigned(512, 10), 197 => to_unsigned(514, 10), 198 => to_unsigned(302, 10), 199 => to_unsigned(604, 10), 200 => to_unsigned(372, 10), 201 => to_unsigned(413, 10), 202 => to_unsigned(408, 10), 203 => to_unsigned(580, 10), 204 => to_unsigned(601, 10), 205 => to_unsigned(513, 10), 206 => to_unsigned(442, 10), 207 => to_unsigned(358, 10), 208 => to_unsigned(462, 10), 209 => to_unsigned(569, 10), 210 => to_unsigned(432, 10), 211 => to_unsigned(462, 10), 212 => to_unsigned(472, 10), 213 => to_unsigned(417, 10), 214 => to_unsigned(553, 10), 215 => to_unsigned(554, 10), 216 => to_unsigned(497, 10), 217 => to_unsigned(568, 10), 218 => to_unsigned(632, 10), 219 => to_unsigned(507, 10), 220 => to_unsigned(620, 10), 221 => to_unsigned(519, 10), 222 => to_unsigned(548, 10), 223 => to_unsigned(559, 10), 224 => to_unsigned(472, 10), 225 => to_unsigned(566, 10), 226 => to_unsigned(571, 10), 227 => to_unsigned(458, 10), 228 => to_unsigned(438, 10), 229 => to_unsigned(621, 10), 230 => to_unsigned(533, 10), 231 => to_unsigned(601, 10), 232 => to_unsigned(415, 10), 233 => to_unsigned(581, 10), 234 => to_unsigned(471, 10), 235 => to_unsigned(772, 10), 236 => to_unsigned(533, 10), 237 => to_unsigned(398, 10), 238 => to_unsigned(513, 10), 239 => to_unsigned(475, 10), 240 => to_unsigned(469, 10), 241 => to_unsigned(571, 10), 242 => to_unsigned(466, 10), 243 => to_unsigned(447, 10), 244 => to_unsigned(450, 10), 245 => to_unsigned(318, 10), 246 => to_unsigned(514, 10), 247 => to_unsigned(495, 10), 248 => to_unsigned(253, 10), 249 => to_unsigned(625, 10), 250 => to_unsigned(390, 10), 251 => to_unsigned(509, 10), 252 => to_unsigned(493, 10), 253 => to_unsigned(428, 10), 254 => to_unsigned(519, 10), 255 => to_unsigned(706, 10), 256 => to_unsigned(407, 10), 257 => to_unsigned(495, 10), 258 => to_unsigned(618, 10), 259 => to_unsigned(559, 10), 260 => to_unsigned(544, 10), 261 => to_unsigned(509, 10), 262 => to_unsigned(585, 10), 263 => to_unsigned(554, 10), 264 => to_unsigned(521, 10), 265 => to_unsigned(566, 10), 266 => to_unsigned(509, 10), 267 => to_unsigned(617, 10), 268 => to_unsigned(407, 10), 269 => to_unsigned(423, 10), 270 => to_unsigned(592, 10), 271 => to_unsigned(444, 10), 272 => to_unsigned(435, 10), 273 => to_unsigned(443, 10), 274 => to_unsigned(524, 10), 275 => to_unsigned(492, 10), 276 => to_unsigned(490, 10), 277 => to_unsigned(620, 10), 278 => to_unsigned(595, 10), 279 => to_unsigned(494, 10), 280 => to_unsigned(461, 10), 281 => to_unsigned(466, 10), 282 => to_unsigned(408, 10), 283 => to_unsigned(512, 10), 284 => to_unsigned(602, 10), 285 => to_unsigned(519, 10), 286 => to_unsigned(346, 10), 287 => to_unsigned(624, 10), 288 => to_unsigned(530, 10), 289 => to_unsigned(465, 10), 290 => to_unsigned(546, 10), 291 => to_unsigned(633, 10), 292 => to_unsigned(516, 10), 293 => to_unsigned(435, 10), 294 => to_unsigned(246, 10), 295 => to_unsigned(414, 10), 296 => to_unsigned(433, 10), 297 => to_unsigned(453, 10), 298 => to_unsigned(550, 10), 299 => to_unsigned(318, 10), 300 => to_unsigned(496, 10), 301 => to_unsigned(592, 10), 302 => to_unsigned(455, 10), 303 => to_unsigned(563, 10), 304 => to_unsigned(478, 10), 305 => to_unsigned(568, 10), 306 => to_unsigned(614, 10), 307 => to_unsigned(597, 10), 308 => to_unsigned(490, 10), 309 => to_unsigned(530, 10), 310 => to_unsigned(439, 10), 311 => to_unsigned(479, 10), 312 => to_unsigned(353, 10), 313 => to_unsigned(554, 10), 314 => to_unsigned(544, 10), 315 => to_unsigned(533, 10), 316 => to_unsigned(620, 10), 317 => to_unsigned(536, 10), 318 => to_unsigned(541, 10), 319 => to_unsigned(536, 10), 320 => to_unsigned(714, 10), 321 => to_unsigned(472, 10), 322 => to_unsigned(483, 10), 323 => to_unsigned(647, 10), 324 => to_unsigned(444, 10), 325 => to_unsigned(542, 10), 326 => to_unsigned(692, 10), 327 => to_unsigned(409, 10), 328 => to_unsigned(578, 10), 329 => to_unsigned(390, 10), 330 => to_unsigned(506, 10), 331 => to_unsigned(376, 10), 332 => to_unsigned(415, 10), 333 => to_unsigned(572, 10), 334 => to_unsigned(370, 10), 335 => to_unsigned(292, 10), 336 => to_unsigned(492, 10), 337 => to_unsigned(491, 10), 338 => to_unsigned(729, 10), 339 => to_unsigned(668, 10), 340 => to_unsigned(503, 10), 341 => to_unsigned(563, 10), 342 => to_unsigned(603, 10), 343 => to_unsigned(587, 10), 344 => to_unsigned(615, 10), 345 => to_unsigned(513, 10), 346 => to_unsigned(583, 10), 347 => to_unsigned(507, 10), 348 => to_unsigned(563, 10), 349 => to_unsigned(399, 10), 350 => to_unsigned(513, 10), 351 => to_unsigned(567, 10), 352 => to_unsigned(342, 10), 353 => to_unsigned(510, 10), 354 => to_unsigned(303, 10), 355 => to_unsigned(421, 10), 356 => to_unsigned(620, 10), 357 => to_unsigned(480, 10), 358 => to_unsigned(549, 10), 359 => to_unsigned(679, 10), 360 => to_unsigned(435, 10), 361 => to_unsigned(415, 10), 362 => to_unsigned(552, 10), 363 => to_unsigned(519, 10), 364 => to_unsigned(466, 10), 365 => to_unsigned(557, 10), 366 => to_unsigned(444, 10), 367 => to_unsigned(515, 10), 368 => to_unsigned(730, 10), 369 => to_unsigned(495, 10), 370 => to_unsigned(379, 10), 371 => to_unsigned(414, 10), 372 => to_unsigned(522, 10), 373 => to_unsigned(551, 10), 374 => to_unsigned(633, 10), 375 => to_unsigned(484, 10), 376 => to_unsigned(628, 10), 377 => to_unsigned(543, 10), 378 => to_unsigned(413, 10), 379 => to_unsigned(395, 10), 380 => to_unsigned(523, 10), 381 => to_unsigned(255, 10), 382 => to_unsigned(575, 10), 383 => to_unsigned(458, 10), 384 => to_unsigned(509, 10), 385 => to_unsigned(411, 10), 386 => to_unsigned(505, 10), 387 => to_unsigned(574, 10), 388 => to_unsigned(536, 10), 389 => to_unsigned(311, 10), 390 => to_unsigned(632, 10), 391 => to_unsigned(550, 10), 392 => to_unsigned(619, 10), 393 => to_unsigned(376, 10), 394 => to_unsigned(574, 10), 395 => to_unsigned(519, 10), 396 => to_unsigned(317, 10), 397 => to_unsigned(416, 10), 398 => to_unsigned(586, 10), 399 => to_unsigned(543, 10), 400 => to_unsigned(516, 10), 401 => to_unsigned(640, 10), 402 => to_unsigned(557, 10), 403 => to_unsigned(665, 10), 404 => to_unsigned(540, 10), 405 => to_unsigned(498, 10), 406 => to_unsigned(594, 10), 407 => to_unsigned(507, 10), 408 => to_unsigned(580, 10), 409 => to_unsigned(476, 10), 410 => to_unsigned(614, 10), 411 => to_unsigned(534, 10), 412 => to_unsigned(530, 10), 413 => to_unsigned(391, 10), 414 => to_unsigned(555, 10), 415 => to_unsigned(603, 10), 416 => to_unsigned(633, 10), 417 => to_unsigned(555, 10), 418 => to_unsigned(425, 10), 419 => to_unsigned(513, 10), 420 => to_unsigned(441, 10), 421 => to_unsigned(330, 10), 422 => to_unsigned(381, 10), 423 => to_unsigned(468, 10), 424 => to_unsigned(539, 10), 425 => to_unsigned(518, 10), 426 => to_unsigned(526, 10), 427 => to_unsigned(382, 10), 428 => to_unsigned(509, 10), 429 => to_unsigned(436, 10), 430 => to_unsigned(411, 10), 431 => to_unsigned(470, 10), 432 => to_unsigned(509, 10), 433 => to_unsigned(485, 10), 434 => to_unsigned(404, 10), 435 => to_unsigned(509, 10), 436 => to_unsigned(449, 10), 437 => to_unsigned(469, 10), 438 => to_unsigned(335, 10), 439 => to_unsigned(464, 10), 440 => to_unsigned(409, 10), 441 => to_unsigned(505, 10), 442 => to_unsigned(587, 10), 443 => to_unsigned(481, 10), 444 => to_unsigned(573, 10), 445 => to_unsigned(599, 10), 446 => to_unsigned(563, 10), 447 => to_unsigned(536, 10), 448 => to_unsigned(487, 10), 449 => to_unsigned(567, 10), 450 => to_unsigned(454, 10), 451 => to_unsigned(492, 10), 452 => to_unsigned(472, 10), 453 => to_unsigned(574, 10), 454 => to_unsigned(531, 10), 455 => to_unsigned(469, 10), 456 => to_unsigned(453, 10), 457 => to_unsigned(410, 10), 458 => to_unsigned(408, 10), 459 => to_unsigned(543, 10), 460 => to_unsigned(467, 10), 461 => to_unsigned(448, 10), 462 => to_unsigned(403, 10), 463 => to_unsigned(613, 10), 464 => to_unsigned(623, 10), 465 => to_unsigned(430, 10), 466 => to_unsigned(324, 10), 467 => to_unsigned(519, 10), 468 => to_unsigned(451, 10), 469 => to_unsigned(423, 10), 470 => to_unsigned(588, 10), 471 => to_unsigned(576, 10), 472 => to_unsigned(699, 10), 473 => to_unsigned(435, 10), 474 => to_unsigned(492, 10), 475 => to_unsigned(545, 10), 476 => to_unsigned(473, 10), 477 => to_unsigned(573, 10), 478 => to_unsigned(624, 10), 479 => to_unsigned(452, 10), 480 => to_unsigned(549, 10), 481 => to_unsigned(548, 10), 482 => to_unsigned(536, 10), 483 => to_unsigned(514, 10), 484 => to_unsigned(548, 10), 485 => to_unsigned(588, 10), 486 => to_unsigned(627, 10), 487 => to_unsigned(548, 10), 488 => to_unsigned(475, 10), 489 => to_unsigned(453, 10), 490 => to_unsigned(259, 10), 491 => to_unsigned(631, 10), 492 => to_unsigned(482, 10), 493 => to_unsigned(425, 10), 494 => to_unsigned(711, 10), 495 => to_unsigned(445, 10), 496 => to_unsigned(490, 10), 497 => to_unsigned(548, 10), 498 => to_unsigned(542, 10), 499 => to_unsigned(506, 10), 500 => to_unsigned(374, 10), 501 => to_unsigned(646, 10), 502 => to_unsigned(544, 10), 503 => to_unsigned(622, 10), 504 => to_unsigned(577, 10), 505 => to_unsigned(513, 10), 506 => to_unsigned(497, 10), 507 => to_unsigned(573, 10), 508 => to_unsigned(643, 10), 509 => to_unsigned(521, 10), 510 => to_unsigned(596, 10), 511 => to_unsigned(591, 10), 512 => to_unsigned(421, 10), 513 => to_unsigned(500, 10), 514 => to_unsigned(564, 10), 515 => to_unsigned(474, 10), 516 => to_unsigned(449, 10), 517 => to_unsigned(501, 10), 518 => to_unsigned(585, 10), 519 => to_unsigned(529, 10), 520 => to_unsigned(441, 10), 521 => to_unsigned(653, 10), 522 => to_unsigned(430, 10), 523 => to_unsigned(390, 10), 524 => to_unsigned(555, 10), 525 => to_unsigned(325, 10), 526 => to_unsigned(400, 10), 527 => to_unsigned(414, 10), 528 => to_unsigned(453, 10), 529 => to_unsigned(495, 10), 530 => to_unsigned(562, 10), 531 => to_unsigned(616, 10), 532 => to_unsigned(545, 10), 533 => to_unsigned(279, 10), 534 => to_unsigned(703, 10), 535 => to_unsigned(290, 10), 536 => to_unsigned(501, 10), 537 => to_unsigned(446, 10), 538 => to_unsigned(434, 10), 539 => to_unsigned(480, 10), 540 => to_unsigned(569, 10), 541 => to_unsigned(587, 10), 542 => to_unsigned(374, 10), 543 => to_unsigned(314, 10), 544 => to_unsigned(463, 10), 545 => to_unsigned(550, 10), 546 => to_unsigned(536, 10), 547 => to_unsigned(455, 10), 548 => to_unsigned(544, 10), 549 => to_unsigned(399, 10), 550 => to_unsigned(692, 10), 551 => to_unsigned(538, 10), 552 => to_unsigned(497, 10), 553 => to_unsigned(620, 10), 554 => to_unsigned(489, 10), 555 => to_unsigned(501, 10), 556 => to_unsigned(608, 10), 557 => to_unsigned(442, 10), 558 => to_unsigned(520, 10), 559 => to_unsigned(479, 10), 560 => to_unsigned(461, 10), 561 => to_unsigned(633, 10), 562 => to_unsigned(633, 10), 563 => to_unsigned(637, 10), 564 => to_unsigned(376, 10), 565 => to_unsigned(451, 10), 566 => to_unsigned(493, 10), 567 => to_unsigned(477, 10), 568 => to_unsigned(405, 10), 569 => to_unsigned(457, 10), 570 => to_unsigned(321, 10), 571 => to_unsigned(456, 10), 572 => to_unsigned(365, 10), 573 => to_unsigned(480, 10), 574 => to_unsigned(728, 10), 575 => to_unsigned(436, 10), 576 => to_unsigned(423, 10), 577 => to_unsigned(417, 10), 578 => to_unsigned(518, 10), 579 => to_unsigned(467, 10), 580 => to_unsigned(508, 10), 581 => to_unsigned(395, 10), 582 => to_unsigned(359, 10), 583 => to_unsigned(535, 10), 584 => to_unsigned(441, 10), 585 => to_unsigned(340, 10), 586 => to_unsigned(468, 10), 587 => to_unsigned(414, 10), 588 => to_unsigned(405, 10), 589 => to_unsigned(486, 10), 590 => to_unsigned(465, 10), 591 => to_unsigned(512, 10), 592 => to_unsigned(469, 10), 593 => to_unsigned(546, 10), 594 => to_unsigned(511, 10), 595 => to_unsigned(378, 10), 596 => to_unsigned(473, 10), 597 => to_unsigned(502, 10), 598 => to_unsigned(405, 10), 599 => to_unsigned(596, 10), 600 => to_unsigned(458, 10), 601 => to_unsigned(574, 10), 602 => to_unsigned(442, 10), 603 => to_unsigned(516, 10), 604 => to_unsigned(570, 10), 605 => to_unsigned(603, 10), 606 => to_unsigned(449, 10), 607 => to_unsigned(544, 10), 608 => to_unsigned(624, 10), 609 => to_unsigned(723, 10), 610 => to_unsigned(396, 10), 611 => to_unsigned(420, 10), 612 => to_unsigned(544, 10), 613 => to_unsigned(451, 10), 614 => to_unsigned(543, 10), 615 => to_unsigned(472, 10), 616 => to_unsigned(418, 10), 617 => to_unsigned(475, 10), 618 => to_unsigned(522, 10), 619 => to_unsigned(446, 10), 620 => to_unsigned(477, 10), 621 => to_unsigned(547, 10), 622 => to_unsigned(509, 10), 623 => to_unsigned(712, 10), 624 => to_unsigned(435, 10), 625 => to_unsigned(627, 10), 626 => to_unsigned(544, 10), 627 => to_unsigned(684, 10), 628 => to_unsigned(459, 10), 629 => to_unsigned(607, 10), 630 => to_unsigned(398, 10), 631 => to_unsigned(463, 10), 632 => to_unsigned(411, 10), 633 => to_unsigned(641, 10), 634 => to_unsigned(385, 10), 635 => to_unsigned(362, 10), 636 => to_unsigned(520, 10), 637 => to_unsigned(539, 10), 638 => to_unsigned(576, 10), 639 => to_unsigned(632, 10), 640 => to_unsigned(573, 10), 641 => to_unsigned(641, 10), 642 => to_unsigned(460, 10), 643 => to_unsigned(487, 10), 644 => to_unsigned(587, 10), 645 => to_unsigned(449, 10), 646 => to_unsigned(550, 10), 647 => to_unsigned(482, 10), 648 => to_unsigned(446, 10), 649 => to_unsigned(387, 10), 650 => to_unsigned(695, 10), 651 => to_unsigned(649, 10), 652 => to_unsigned(463, 10), 653 => to_unsigned(369, 10), 654 => to_unsigned(468, 10), 655 => to_unsigned(411, 10), 656 => to_unsigned(419, 10), 657 => to_unsigned(588, 10), 658 => to_unsigned(316, 10), 659 => to_unsigned(596, 10), 660 => to_unsigned(493, 10), 661 => to_unsigned(600, 10), 662 => to_unsigned(537, 10), 663 => to_unsigned(497, 10), 664 => to_unsigned(409, 10), 665 => to_unsigned(468, 10), 666 => to_unsigned(323, 10), 667 => to_unsigned(378, 10), 668 => to_unsigned(458, 10), 669 => to_unsigned(684, 10), 670 => to_unsigned(456, 10), 671 => to_unsigned(390, 10), 672 => to_unsigned(542, 10), 673 => to_unsigned(509, 10), 674 => to_unsigned(624, 10), 675 => to_unsigned(638, 10), 676 => to_unsigned(414, 10), 677 => to_unsigned(516, 10), 678 => to_unsigned(479, 10), 679 => to_unsigned(510, 10), 680 => to_unsigned(454, 10), 681 => to_unsigned(605, 10), 682 => to_unsigned(576, 10), 683 => to_unsigned(592, 10), 684 => to_unsigned(557, 10), 685 => to_unsigned(514, 10), 686 => to_unsigned(628, 10), 687 => to_unsigned(528, 10), 688 => to_unsigned(570, 10), 689 => to_unsigned(642, 10), 690 => to_unsigned(495, 10), 691 => to_unsigned(529, 10), 692 => to_unsigned(474, 10), 693 => to_unsigned(555, 10), 694 => to_unsigned(655, 10), 695 => to_unsigned(445, 10), 696 => to_unsigned(613, 10), 697 => to_unsigned(502, 10), 698 => to_unsigned(523, 10), 699 => to_unsigned(350, 10), 700 => to_unsigned(602, 10), 701 => to_unsigned(482, 10), 702 => to_unsigned(570, 10), 703 => to_unsigned(557, 10), 704 => to_unsigned(423, 10), 705 => to_unsigned(498, 10), 706 => to_unsigned(683, 10), 707 => to_unsigned(499, 10), 708 => to_unsigned(589, 10), 709 => to_unsigned(405, 10), 710 => to_unsigned(516, 10), 711 => to_unsigned(426, 10), 712 => to_unsigned(507, 10), 713 => to_unsigned(381, 10), 714 => to_unsigned(546, 10), 715 => to_unsigned(353, 10), 716 => to_unsigned(505, 10), 717 => to_unsigned(460, 10), 718 => to_unsigned(481, 10), 719 => to_unsigned(655, 10), 720 => to_unsigned(647, 10), 721 => to_unsigned(493, 10), 722 => to_unsigned(475, 10), 723 => to_unsigned(498, 10), 724 => to_unsigned(697, 10), 725 => to_unsigned(352, 10), 726 => to_unsigned(404, 10), 727 => to_unsigned(499, 10), 728 => to_unsigned(535, 10), 729 => to_unsigned(508, 10), 730 => to_unsigned(345, 10), 731 => to_unsigned(529, 10), 732 => to_unsigned(479, 10), 733 => to_unsigned(653, 10), 734 => to_unsigned(516, 10), 735 => to_unsigned(658, 10), 736 => to_unsigned(453, 10), 737 => to_unsigned(407, 10), 738 => to_unsigned(328, 10), 739 => to_unsigned(397, 10), 740 => to_unsigned(391, 10), 741 => to_unsigned(394, 10), 742 => to_unsigned(461, 10), 743 => to_unsigned(351, 10), 744 => to_unsigned(602, 10), 745 => to_unsigned(502, 10), 746 => to_unsigned(645, 10), 747 => to_unsigned(442, 10), 748 => to_unsigned(549, 10), 749 => to_unsigned(622, 10), 750 => to_unsigned(469, 10), 751 => to_unsigned(300, 10), 752 => to_unsigned(292, 10), 753 => to_unsigned(542, 10), 754 => to_unsigned(443, 10), 755 => to_unsigned(544, 10), 756 => to_unsigned(469, 10), 757 => to_unsigned(563, 10), 758 => to_unsigned(512, 10), 759 => to_unsigned(361, 10), 760 => to_unsigned(543, 10), 761 => to_unsigned(556, 10), 762 => to_unsigned(640, 10), 763 => to_unsigned(389, 10), 764 => to_unsigned(463, 10), 765 => to_unsigned(601, 10), 766 => to_unsigned(520, 10), 767 => to_unsigned(458, 10), 768 => to_unsigned(329, 10), 769 => to_unsigned(497, 10), 770 => to_unsigned(418, 10), 771 => to_unsigned(481, 10), 772 => to_unsigned(380, 10), 773 => to_unsigned(503, 10), 774 => to_unsigned(502, 10), 775 => to_unsigned(558, 10), 776 => to_unsigned(568, 10), 777 => to_unsigned(469, 10), 778 => to_unsigned(380, 10), 779 => to_unsigned(525, 10), 780 => to_unsigned(432, 10), 781 => to_unsigned(565, 10), 782 => to_unsigned(451, 10), 783 => to_unsigned(531, 10), 784 => to_unsigned(591, 10), 785 => to_unsigned(385, 10), 786 => to_unsigned(573, 10), 787 => to_unsigned(374, 10), 788 => to_unsigned(648, 10), 789 => to_unsigned(425, 10), 790 => to_unsigned(619, 10), 791 => to_unsigned(460, 10), 792 => to_unsigned(621, 10), 793 => to_unsigned(637, 10), 794 => to_unsigned(659, 10), 795 => to_unsigned(529, 10), 796 => to_unsigned(469, 10), 797 => to_unsigned(709, 10), 798 => to_unsigned(443, 10), 799 => to_unsigned(545, 10), 800 => to_unsigned(486, 10), 801 => to_unsigned(616, 10), 802 => to_unsigned(455, 10), 803 => to_unsigned(442, 10), 804 => to_unsigned(451, 10), 805 => to_unsigned(377, 10), 806 => to_unsigned(457, 10), 807 => to_unsigned(427, 10), 808 => to_unsigned(580, 10), 809 => to_unsigned(510, 10), 810 => to_unsigned(547, 10), 811 => to_unsigned(462, 10), 812 => to_unsigned(504, 10), 813 => to_unsigned(399, 10), 814 => to_unsigned(526, 10), 815 => to_unsigned(328, 10), 816 => to_unsigned(423, 10), 817 => to_unsigned(544, 10), 818 => to_unsigned(586, 10), 819 => to_unsigned(511, 10), 820 => to_unsigned(415, 10), 821 => to_unsigned(566, 10), 822 => to_unsigned(350, 10), 823 => to_unsigned(575, 10), 824 => to_unsigned(461, 10), 825 => to_unsigned(386, 10), 826 => to_unsigned(393, 10), 827 => to_unsigned(509, 10), 828 => to_unsigned(580, 10), 829 => to_unsigned(547, 10), 830 => to_unsigned(304, 10), 831 => to_unsigned(482, 10), 832 => to_unsigned(551, 10), 833 => to_unsigned(504, 10), 834 => to_unsigned(565, 10), 835 => to_unsigned(223, 10), 836 => to_unsigned(507, 10), 837 => to_unsigned(414, 10), 838 => to_unsigned(687, 10), 839 => to_unsigned(494, 10), 840 => to_unsigned(514, 10), 841 => to_unsigned(484, 10), 842 => to_unsigned(572, 10), 843 => to_unsigned(580, 10), 844 => to_unsigned(439, 10), 845 => to_unsigned(402, 10), 846 => to_unsigned(478, 10), 847 => to_unsigned(628, 10), 848 => to_unsigned(472, 10), 849 => to_unsigned(518, 10), 850 => to_unsigned(415, 10), 851 => to_unsigned(420, 10), 852 => to_unsigned(500, 10), 853 => to_unsigned(518, 10), 854 => to_unsigned(452, 10), 855 => to_unsigned(548, 10), 856 => to_unsigned(501, 10), 857 => to_unsigned(376, 10), 858 => to_unsigned(475, 10), 859 => to_unsigned(359, 10), 860 => to_unsigned(603, 10), 861 => to_unsigned(443, 10), 862 => to_unsigned(530, 10), 863 => to_unsigned(394, 10), 864 => to_unsigned(546, 10), 865 => to_unsigned(608, 10), 866 => to_unsigned(595, 10), 867 => to_unsigned(542, 10), 868 => to_unsigned(376, 10), 869 => to_unsigned(445, 10), 870 => to_unsigned(479, 10), 871 => to_unsigned(448, 10), 872 => to_unsigned(511, 10), 873 => to_unsigned(453, 10), 874 => to_unsigned(422, 10), 875 => to_unsigned(571, 10), 876 => to_unsigned(460, 10), 877 => to_unsigned(586, 10), 878 => to_unsigned(635, 10), 879 => to_unsigned(503, 10), 880 => to_unsigned(624, 10), 881 => to_unsigned(425, 10), 882 => to_unsigned(550, 10), 883 => to_unsigned(436, 10), 884 => to_unsigned(587, 10), 885 => to_unsigned(546, 10), 886 => to_unsigned(639, 10), 887 => to_unsigned(591, 10), 888 => to_unsigned(419, 10), 889 => to_unsigned(440, 10), 890 => to_unsigned(556, 10), 891 => to_unsigned(586, 10), 892 => to_unsigned(589, 10), 893 => to_unsigned(392, 10), 894 => to_unsigned(566, 10), 895 => to_unsigned(529, 10), 896 => to_unsigned(410, 10), 897 => to_unsigned(626, 10), 898 => to_unsigned(477, 10), 899 => to_unsigned(636, 10), 900 => to_unsigned(461, 10), 901 => to_unsigned(366, 10), 902 => to_unsigned(453, 10), 903 => to_unsigned(371, 10), 904 => to_unsigned(640, 10), 905 => to_unsigned(463, 10), 906 => to_unsigned(554, 10), 907 => to_unsigned(309, 10), 908 => to_unsigned(478, 10), 909 => to_unsigned(604, 10), 910 => to_unsigned(585, 10), 911 => to_unsigned(528, 10), 912 => to_unsigned(466, 10), 913 => to_unsigned(675, 10), 914 => to_unsigned(532, 10), 915 => to_unsigned(526, 10), 916 => to_unsigned(508, 10), 917 => to_unsigned(554, 10), 918 => to_unsigned(555, 10), 919 => to_unsigned(461, 10), 920 => to_unsigned(550, 10), 921 => to_unsigned(320, 10), 922 => to_unsigned(713, 10), 923 => to_unsigned(427, 10), 924 => to_unsigned(372, 10), 925 => to_unsigned(519, 10), 926 => to_unsigned(772, 10), 927 => to_unsigned(484, 10), 928 => to_unsigned(538, 10), 929 => to_unsigned(526, 10), 930 => to_unsigned(580, 10), 931 => to_unsigned(509, 10), 932 => to_unsigned(520, 10), 933 => to_unsigned(475, 10), 934 => to_unsigned(625, 10), 935 => to_unsigned(368, 10), 936 => to_unsigned(712, 10), 937 => to_unsigned(523, 10), 938 => to_unsigned(602, 10), 939 => to_unsigned(600, 10), 940 => to_unsigned(390, 10), 941 => to_unsigned(451, 10), 942 => to_unsigned(418, 10), 943 => to_unsigned(436, 10), 944 => to_unsigned(536, 10), 945 => to_unsigned(437, 10), 946 => to_unsigned(440, 10), 947 => to_unsigned(596, 10), 948 => to_unsigned(441, 10), 949 => to_unsigned(510, 10), 950 => to_unsigned(444, 10), 951 => to_unsigned(504, 10), 952 => to_unsigned(485, 10), 953 => to_unsigned(703, 10), 954 => to_unsigned(330, 10), 955 => to_unsigned(547, 10), 956 => to_unsigned(484, 10), 957 => to_unsigned(409, 10), 958 => to_unsigned(695, 10), 959 => to_unsigned(454, 10), 960 => to_unsigned(360, 10), 961 => to_unsigned(613, 10), 962 => to_unsigned(608, 10), 963 => to_unsigned(597, 10), 964 => to_unsigned(457, 10), 965 => to_unsigned(555, 10), 966 => to_unsigned(527, 10), 967 => to_unsigned(421, 10), 968 => to_unsigned(519, 10), 969 => to_unsigned(446, 10), 970 => to_unsigned(556, 10), 971 => to_unsigned(518, 10), 972 => to_unsigned(436, 10), 973 => to_unsigned(453, 10), 974 => to_unsigned(460, 10), 975 => to_unsigned(432, 10), 976 => to_unsigned(447, 10), 977 => to_unsigned(542, 10), 978 => to_unsigned(525, 10), 979 => to_unsigned(571, 10), 980 => to_unsigned(408, 10), 981 => to_unsigned(564, 10), 982 => to_unsigned(419, 10), 983 => to_unsigned(491, 10), 984 => to_unsigned(449, 10), 985 => to_unsigned(450, 10), 986 => to_unsigned(444, 10), 987 => to_unsigned(596, 10), 988 => to_unsigned(468, 10), 989 => to_unsigned(627, 10), 990 => to_unsigned(639, 10), 991 => to_unsigned(621, 10), 992 => to_unsigned(403, 10), 993 => to_unsigned(412, 10), 994 => to_unsigned(536, 10), 995 => to_unsigned(663, 10), 996 => to_unsigned(581, 10), 997 => to_unsigned(656, 10), 998 => to_unsigned(440, 10), 999 => to_unsigned(610, 10), 1000 => to_unsigned(524, 10), 1001 => to_unsigned(492, 10), 1002 => to_unsigned(560, 10), 1003 => to_unsigned(540, 10), 1004 => to_unsigned(616, 10), 1005 => to_unsigned(445, 10), 1006 => to_unsigned(551, 10), 1007 => to_unsigned(532, 10), 1008 => to_unsigned(462, 10), 1009 => to_unsigned(597, 10), 1010 => to_unsigned(400, 10), 1011 => to_unsigned(567, 10), 1012 => to_unsigned(599, 10), 1013 => to_unsigned(499, 10), 1014 => to_unsigned(583, 10), 1015 => to_unsigned(564, 10), 1016 => to_unsigned(455, 10), 1017 => to_unsigned(352, 10), 1018 => to_unsigned(608, 10), 1019 => to_unsigned(626, 10), 1020 => to_unsigned(607, 10), 1021 => to_unsigned(434, 10), 1022 => to_unsigned(546, 10), 1023 => to_unsigned(679, 10), 1024 => to_unsigned(544, 10), 1025 => to_unsigned(567, 10), 1026 => to_unsigned(537, 10), 1027 => to_unsigned(556, 10), 1028 => to_unsigned(543, 10), 1029 => to_unsigned(630, 10), 1030 => to_unsigned(394, 10), 1031 => to_unsigned(558, 10), 1032 => to_unsigned(399, 10), 1033 => to_unsigned(486, 10), 1034 => to_unsigned(526, 10), 1035 => to_unsigned(533, 10), 1036 => to_unsigned(315, 10), 1037 => to_unsigned(465, 10), 1038 => to_unsigned(512, 10), 1039 => to_unsigned(610, 10), 1040 => to_unsigned(504, 10), 1041 => to_unsigned(524, 10), 1042 => to_unsigned(510, 10), 1043 => to_unsigned(415, 10), 1044 => to_unsigned(401, 10), 1045 => to_unsigned(403, 10), 1046 => to_unsigned(361, 10), 1047 => to_unsigned(552, 10), 1048 => to_unsigned(481, 10), 1049 => to_unsigned(702, 10), 1050 => to_unsigned(396, 10), 1051 => to_unsigned(506, 10), 1052 => to_unsigned(462, 10), 1053 => to_unsigned(505, 10), 1054 => to_unsigned(536, 10), 1055 => to_unsigned(505, 10), 1056 => to_unsigned(578, 10), 1057 => to_unsigned(592, 10), 1058 => to_unsigned(545, 10), 1059 => to_unsigned(570, 10), 1060 => to_unsigned(648, 10), 1061 => to_unsigned(618, 10), 1062 => to_unsigned(607, 10), 1063 => to_unsigned(555, 10), 1064 => to_unsigned(479, 10), 1065 => to_unsigned(709, 10), 1066 => to_unsigned(488, 10), 1067 => to_unsigned(514, 10), 1068 => to_unsigned(321, 10), 1069 => to_unsigned(520, 10), 1070 => to_unsigned(519, 10), 1071 => to_unsigned(517, 10), 1072 => to_unsigned(649, 10), 1073 => to_unsigned(428, 10), 1074 => to_unsigned(498, 10), 1075 => to_unsigned(499, 10), 1076 => to_unsigned(378, 10), 1077 => to_unsigned(562, 10), 1078 => to_unsigned(594, 10), 1079 => to_unsigned(381, 10), 1080 => to_unsigned(570, 10), 1081 => to_unsigned(560, 10), 1082 => to_unsigned(561, 10), 1083 => to_unsigned(573, 10), 1084 => to_unsigned(506, 10), 1085 => to_unsigned(384, 10), 1086 => to_unsigned(537, 10), 1087 => to_unsigned(632, 10), 1088 => to_unsigned(480, 10), 1089 => to_unsigned(421, 10), 1090 => to_unsigned(501, 10), 1091 => to_unsigned(467, 10), 1092 => to_unsigned(425, 10), 1093 => to_unsigned(519, 10), 1094 => to_unsigned(489, 10), 1095 => to_unsigned(528, 10), 1096 => to_unsigned(575, 10), 1097 => to_unsigned(366, 10), 1098 => to_unsigned(504, 10), 1099 => to_unsigned(556, 10), 1100 => to_unsigned(566, 10), 1101 => to_unsigned(352, 10), 1102 => to_unsigned(542, 10), 1103 => to_unsigned(428, 10), 1104 => to_unsigned(463, 10), 1105 => to_unsigned(531, 10), 1106 => to_unsigned(385, 10), 1107 => to_unsigned(603, 10), 1108 => to_unsigned(521, 10), 1109 => to_unsigned(651, 10), 1110 => to_unsigned(538, 10), 1111 => to_unsigned(510, 10), 1112 => to_unsigned(588, 10), 1113 => to_unsigned(384, 10), 1114 => to_unsigned(384, 10), 1115 => to_unsigned(496, 10), 1116 => to_unsigned(573, 10), 1117 => to_unsigned(623, 10), 1118 => to_unsigned(642, 10), 1119 => to_unsigned(496, 10), 1120 => to_unsigned(631, 10), 1121 => to_unsigned(600, 10), 1122 => to_unsigned(503, 10), 1123 => to_unsigned(536, 10), 1124 => to_unsigned(486, 10), 1125 => to_unsigned(476, 10), 1126 => to_unsigned(570, 10), 1127 => to_unsigned(613, 10), 1128 => to_unsigned(505, 10), 1129 => to_unsigned(558, 10), 1130 => to_unsigned(502, 10), 1131 => to_unsigned(461, 10), 1132 => to_unsigned(594, 10), 1133 => to_unsigned(455, 10), 1134 => to_unsigned(433, 10), 1135 => to_unsigned(634, 10), 1136 => to_unsigned(527, 10), 1137 => to_unsigned(453, 10), 1138 => to_unsigned(523, 10), 1139 => to_unsigned(578, 10), 1140 => to_unsigned(602, 10), 1141 => to_unsigned(620, 10), 1142 => to_unsigned(700, 10), 1143 => to_unsigned(546, 10), 1144 => to_unsigned(610, 10), 1145 => to_unsigned(622, 10), 1146 => to_unsigned(506, 10), 1147 => to_unsigned(497, 10), 1148 => to_unsigned(609, 10), 1149 => to_unsigned(590, 10), 1150 => to_unsigned(590, 10), 1151 => to_unsigned(443, 10), 1152 => to_unsigned(437, 10), 1153 => to_unsigned(506, 10), 1154 => to_unsigned(560, 10), 1155 => to_unsigned(501, 10), 1156 => to_unsigned(606, 10), 1157 => to_unsigned(536, 10), 1158 => to_unsigned(407, 10), 1159 => to_unsigned(456, 10), 1160 => to_unsigned(626, 10), 1161 => to_unsigned(582, 10), 1162 => to_unsigned(566, 10), 1163 => to_unsigned(538, 10), 1164 => to_unsigned(515, 10), 1165 => to_unsigned(703, 10), 1166 => to_unsigned(537, 10), 1167 => to_unsigned(534, 10), 1168 => to_unsigned(600, 10), 1169 => to_unsigned(439, 10), 1170 => to_unsigned(394, 10), 1171 => to_unsigned(378, 10), 1172 => to_unsigned(346, 10), 1173 => to_unsigned(687, 10), 1174 => to_unsigned(634, 10), 1175 => to_unsigned(477, 10), 1176 => to_unsigned(273, 10), 1177 => to_unsigned(594, 10), 1178 => to_unsigned(398, 10), 1179 => to_unsigned(333, 10), 1180 => to_unsigned(411, 10), 1181 => to_unsigned(637, 10), 1182 => to_unsigned(412, 10), 1183 => to_unsigned(593, 10), 1184 => to_unsigned(388, 10), 1185 => to_unsigned(475, 10), 1186 => to_unsigned(558, 10), 1187 => to_unsigned(461, 10), 1188 => to_unsigned(496, 10), 1189 => to_unsigned(519, 10), 1190 => to_unsigned(458, 10), 1191 => to_unsigned(445, 10), 1192 => to_unsigned(425, 10), 1193 => to_unsigned(418, 10), 1194 => to_unsigned(813, 10), 1195 => to_unsigned(507, 10), 1196 => to_unsigned(524, 10), 1197 => to_unsigned(652, 10), 1198 => to_unsigned(694, 10), 1199 => to_unsigned(539, 10), 1200 => to_unsigned(440, 10), 1201 => to_unsigned(561, 10), 1202 => to_unsigned(633, 10), 1203 => to_unsigned(625, 10), 1204 => to_unsigned(762, 10), 1205 => to_unsigned(601, 10), 1206 => to_unsigned(598, 10), 1207 => to_unsigned(477, 10), 1208 => to_unsigned(492, 10), 1209 => to_unsigned(551, 10), 1210 => to_unsigned(491, 10), 1211 => to_unsigned(476, 10), 1212 => to_unsigned(524, 10), 1213 => to_unsigned(467, 10), 1214 => to_unsigned(632, 10), 1215 => to_unsigned(503, 10), 1216 => to_unsigned(455, 10), 1217 => to_unsigned(531, 10), 1218 => to_unsigned(599, 10), 1219 => to_unsigned(559, 10), 1220 => to_unsigned(548, 10), 1221 => to_unsigned(438, 10), 1222 => to_unsigned(364, 10), 1223 => to_unsigned(476, 10), 1224 => to_unsigned(407, 10), 1225 => to_unsigned(551, 10), 1226 => to_unsigned(399, 10), 1227 => to_unsigned(388, 10), 1228 => to_unsigned(624, 10), 1229 => to_unsigned(529, 10), 1230 => to_unsigned(451, 10), 1231 => to_unsigned(537, 10), 1232 => to_unsigned(608, 10), 1233 => to_unsigned(556, 10), 1234 => to_unsigned(521, 10), 1235 => to_unsigned(470, 10), 1236 => to_unsigned(624, 10), 1237 => to_unsigned(602, 10), 1238 => to_unsigned(458, 10), 1239 => to_unsigned(501, 10), 1240 => to_unsigned(463, 10), 1241 => to_unsigned(504, 10), 1242 => to_unsigned(501, 10), 1243 => to_unsigned(609, 10), 1244 => to_unsigned(564, 10), 1245 => to_unsigned(491, 10), 1246 => to_unsigned(523, 10), 1247 => to_unsigned(646, 10), 1248 => to_unsigned(556, 10), 1249 => to_unsigned(616, 10), 1250 => to_unsigned(633, 10), 1251 => to_unsigned(456, 10), 1252 => to_unsigned(552, 10), 1253 => to_unsigned(550, 10), 1254 => to_unsigned(532, 10), 1255 => to_unsigned(409, 10), 1256 => to_unsigned(432, 10), 1257 => to_unsigned(524, 10), 1258 => to_unsigned(542, 10), 1259 => to_unsigned(473, 10), 1260 => to_unsigned(468, 10), 1261 => to_unsigned(391, 10), 1262 => to_unsigned(439, 10), 1263 => to_unsigned(462, 10), 1264 => to_unsigned(514, 10), 1265 => to_unsigned(402, 10), 1266 => to_unsigned(563, 10), 1267 => to_unsigned(494, 10), 1268 => to_unsigned(421, 10), 1269 => to_unsigned(589, 10), 1270 => to_unsigned(459, 10), 1271 => to_unsigned(527, 10), 1272 => to_unsigned(438, 10), 1273 => to_unsigned(503, 10), 1274 => to_unsigned(519, 10), 1275 => to_unsigned(583, 10), 1276 => to_unsigned(521, 10), 1277 => to_unsigned(743, 10), 1278 => to_unsigned(508, 10), 1279 => to_unsigned(454, 10), 1280 => to_unsigned(638, 10), 1281 => to_unsigned(681, 10), 1282 => to_unsigned(492, 10), 1283 => to_unsigned(557, 10), 1284 => to_unsigned(446, 10), 1285 => to_unsigned(542, 10), 1286 => to_unsigned(471, 10), 1287 => to_unsigned(457, 10), 1288 => to_unsigned(366, 10), 1289 => to_unsigned(601, 10), 1290 => to_unsigned(589, 10), 1291 => to_unsigned(455, 10), 1292 => to_unsigned(532, 10), 1293 => to_unsigned(520, 10), 1294 => to_unsigned(346, 10), 1295 => to_unsigned(629, 10), 1296 => to_unsigned(468, 10), 1297 => to_unsigned(498, 10), 1298 => to_unsigned(471, 10), 1299 => to_unsigned(596, 10), 1300 => to_unsigned(527, 10), 1301 => to_unsigned(567, 10), 1302 => to_unsigned(578, 10), 1303 => to_unsigned(487, 10), 1304 => to_unsigned(496, 10), 1305 => to_unsigned(509, 10), 1306 => to_unsigned(494, 10), 1307 => to_unsigned(453, 10), 1308 => to_unsigned(514, 10), 1309 => to_unsigned(533, 10), 1310 => to_unsigned(466, 10), 1311 => to_unsigned(441, 10), 1312 => to_unsigned(428, 10), 1313 => to_unsigned(647, 10), 1314 => to_unsigned(565, 10), 1315 => to_unsigned(440, 10), 1316 => to_unsigned(514, 10), 1317 => to_unsigned(403, 10), 1318 => to_unsigned(510, 10), 1319 => to_unsigned(324, 10), 1320 => to_unsigned(509, 10), 1321 => to_unsigned(414, 10), 1322 => to_unsigned(439, 10), 1323 => to_unsigned(463, 10), 1324 => to_unsigned(635, 10), 1325 => to_unsigned(655, 10), 1326 => to_unsigned(530, 10), 1327 => to_unsigned(342, 10), 1328 => to_unsigned(382, 10), 1329 => to_unsigned(550, 10), 1330 => to_unsigned(673, 10), 1331 => to_unsigned(554, 10), 1332 => to_unsigned(420, 10), 1333 => to_unsigned(341, 10), 1334 => to_unsigned(413, 10), 1335 => to_unsigned(538, 10), 1336 => to_unsigned(573, 10), 1337 => to_unsigned(440, 10), 1338 => to_unsigned(629, 10), 1339 => to_unsigned(600, 10), 1340 => to_unsigned(425, 10), 1341 => to_unsigned(641, 10), 1342 => to_unsigned(561, 10), 1343 => to_unsigned(542, 10), 1344 => to_unsigned(429, 10), 1345 => to_unsigned(629, 10), 1346 => to_unsigned(471, 10), 1347 => to_unsigned(630, 10), 1348 => to_unsigned(570, 10), 1349 => to_unsigned(441, 10), 1350 => to_unsigned(589, 10), 1351 => to_unsigned(500, 10), 1352 => to_unsigned(402, 10), 1353 => to_unsigned(542, 10), 1354 => to_unsigned(473, 10), 1355 => to_unsigned(609, 10), 1356 => to_unsigned(502, 10), 1357 => to_unsigned(470, 10), 1358 => to_unsigned(478, 10), 1359 => to_unsigned(338, 10), 1360 => to_unsigned(647, 10), 1361 => to_unsigned(491, 10), 1362 => to_unsigned(438, 10), 1363 => to_unsigned(635, 10), 1364 => to_unsigned(532, 10), 1365 => to_unsigned(462, 10), 1366 => to_unsigned(588, 10), 1367 => to_unsigned(526, 10), 1368 => to_unsigned(319, 10), 1369 => to_unsigned(461, 10), 1370 => to_unsigned(572, 10), 1371 => to_unsigned(569, 10), 1372 => to_unsigned(623, 10), 1373 => to_unsigned(585, 10), 1374 => to_unsigned(472, 10), 1375 => to_unsigned(477, 10), 1376 => to_unsigned(661, 10), 1377 => to_unsigned(674, 10), 1378 => to_unsigned(529, 10), 1379 => to_unsigned(371, 10), 1380 => to_unsigned(548, 10), 1381 => to_unsigned(429, 10), 1382 => to_unsigned(290, 10), 1383 => to_unsigned(374, 10), 1384 => to_unsigned(524, 10), 1385 => to_unsigned(536, 10), 1386 => to_unsigned(614, 10), 1387 => to_unsigned(484, 10), 1388 => to_unsigned(384, 10), 1389 => to_unsigned(492, 10), 1390 => to_unsigned(596, 10), 1391 => to_unsigned(547, 10), 1392 => to_unsigned(675, 10), 1393 => to_unsigned(307, 10), 1394 => to_unsigned(386, 10), 1395 => to_unsigned(543, 10), 1396 => to_unsigned(531, 10), 1397 => to_unsigned(532, 10), 1398 => to_unsigned(338, 10), 1399 => to_unsigned(513, 10), 1400 => to_unsigned(453, 10), 1401 => to_unsigned(594, 10), 1402 => to_unsigned(376, 10), 1403 => to_unsigned(529, 10), 1404 => to_unsigned(494, 10), 1405 => to_unsigned(693, 10), 1406 => to_unsigned(705, 10), 1407 => to_unsigned(333, 10), 1408 => to_unsigned(595, 10), 1409 => to_unsigned(652, 10), 1410 => to_unsigned(476, 10), 1411 => to_unsigned(571, 10), 1412 => to_unsigned(563, 10), 1413 => to_unsigned(553, 10), 1414 => to_unsigned(470, 10), 1415 => to_unsigned(529, 10), 1416 => to_unsigned(519, 10), 1417 => to_unsigned(555, 10), 1418 => to_unsigned(482, 10), 1419 => to_unsigned(523, 10), 1420 => to_unsigned(663, 10), 1421 => to_unsigned(485, 10), 1422 => to_unsigned(347, 10), 1423 => to_unsigned(572, 10), 1424 => to_unsigned(530, 10), 1425 => to_unsigned(404, 10), 1426 => to_unsigned(321, 10), 1427 => to_unsigned(455, 10), 1428 => to_unsigned(486, 10), 1429 => to_unsigned(548, 10), 1430 => to_unsigned(344, 10), 1431 => to_unsigned(559, 10), 1432 => to_unsigned(620, 10), 1433 => to_unsigned(576, 10), 1434 => to_unsigned(653, 10), 1435 => to_unsigned(315, 10), 1436 => to_unsigned(522, 10), 1437 => to_unsigned(527, 10), 1438 => to_unsigned(577, 10), 1439 => to_unsigned(348, 10), 1440 => to_unsigned(455, 10), 1441 => to_unsigned(516, 10), 1442 => to_unsigned(405, 10), 1443 => to_unsigned(534, 10), 1444 => to_unsigned(466, 10), 1445 => to_unsigned(633, 10), 1446 => to_unsigned(432, 10), 1447 => to_unsigned(458, 10), 1448 => to_unsigned(652, 10), 1449 => to_unsigned(599, 10), 1450 => to_unsigned(691, 10), 1451 => to_unsigned(585, 10), 1452 => to_unsigned(487, 10), 1453 => to_unsigned(628, 10), 1454 => to_unsigned(502, 10), 1455 => to_unsigned(586, 10), 1456 => to_unsigned(516, 10), 1457 => to_unsigned(565, 10), 1458 => to_unsigned(593, 10), 1459 => to_unsigned(488, 10), 1460 => to_unsigned(585, 10), 1461 => to_unsigned(476, 10), 1462 => to_unsigned(480, 10), 1463 => to_unsigned(485, 10), 1464 => to_unsigned(594, 10), 1465 => to_unsigned(522, 10), 1466 => to_unsigned(585, 10), 1467 => to_unsigned(599, 10), 1468 => to_unsigned(250, 10), 1469 => to_unsigned(400, 10), 1470 => to_unsigned(594, 10), 1471 => to_unsigned(694, 10), 1472 => to_unsigned(597, 10), 1473 => to_unsigned(577, 10), 1474 => to_unsigned(558, 10), 1475 => to_unsigned(530, 10), 1476 => to_unsigned(582, 10), 1477 => to_unsigned(419, 10), 1478 => to_unsigned(693, 10), 1479 => to_unsigned(446, 10), 1480 => to_unsigned(638, 10), 1481 => to_unsigned(452, 10), 1482 => to_unsigned(583, 10), 1483 => to_unsigned(611, 10), 1484 => to_unsigned(292, 10), 1485 => to_unsigned(451, 10), 1486 => to_unsigned(384, 10), 1487 => to_unsigned(593, 10), 1488 => to_unsigned(424, 10), 1489 => to_unsigned(599, 10), 1490 => to_unsigned(477, 10), 1491 => to_unsigned(522, 10), 1492 => to_unsigned(508, 10), 1493 => to_unsigned(449, 10), 1494 => to_unsigned(460, 10), 1495 => to_unsigned(526, 10), 1496 => to_unsigned(628, 10), 1497 => to_unsigned(517, 10), 1498 => to_unsigned(410, 10), 1499 => to_unsigned(485, 10), 1500 => to_unsigned(510, 10), 1501 => to_unsigned(501, 10), 1502 => to_unsigned(348, 10), 1503 => to_unsigned(448, 10), 1504 => to_unsigned(588, 10), 1505 => to_unsigned(607, 10), 1506 => to_unsigned(601, 10), 1507 => to_unsigned(373, 10), 1508 => to_unsigned(600, 10), 1509 => to_unsigned(615, 10), 1510 => to_unsigned(463, 10), 1511 => to_unsigned(620, 10), 1512 => to_unsigned(510, 10), 1513 => to_unsigned(570, 10), 1514 => to_unsigned(417, 10), 1515 => to_unsigned(485, 10), 1516 => to_unsigned(523, 10), 1517 => to_unsigned(538, 10), 1518 => to_unsigned(490, 10), 1519 => to_unsigned(444, 10), 1520 => to_unsigned(389, 10), 1521 => to_unsigned(362, 10), 1522 => to_unsigned(661, 10), 1523 => to_unsigned(443, 10), 1524 => to_unsigned(414, 10), 1525 => to_unsigned(680, 10), 1526 => to_unsigned(542, 10), 1527 => to_unsigned(528, 10), 1528 => to_unsigned(461, 10), 1529 => to_unsigned(373, 10), 1530 => to_unsigned(502, 10), 1531 => to_unsigned(542, 10), 1532 => to_unsigned(451, 10), 1533 => to_unsigned(460, 10), 1534 => to_unsigned(533, 10), 1535 => to_unsigned(462, 10), 1536 => to_unsigned(611, 10), 1537 => to_unsigned(602, 10), 1538 => to_unsigned(505, 10), 1539 => to_unsigned(656, 10), 1540 => to_unsigned(464, 10), 1541 => to_unsigned(395, 10), 1542 => to_unsigned(479, 10), 1543 => to_unsigned(548, 10), 1544 => to_unsigned(454, 10), 1545 => to_unsigned(520, 10), 1546 => to_unsigned(592, 10), 1547 => to_unsigned(540, 10), 1548 => to_unsigned(434, 10), 1549 => to_unsigned(520, 10), 1550 => to_unsigned(653, 10), 1551 => to_unsigned(466, 10), 1552 => to_unsigned(646, 10), 1553 => to_unsigned(619, 10), 1554 => to_unsigned(460, 10), 1555 => to_unsigned(533, 10), 1556 => to_unsigned(577, 10), 1557 => to_unsigned(559, 10), 1558 => to_unsigned(441, 10), 1559 => to_unsigned(525, 10), 1560 => to_unsigned(481, 10), 1561 => to_unsigned(646, 10), 1562 => to_unsigned(302, 10), 1563 => to_unsigned(456, 10), 1564 => to_unsigned(461, 10), 1565 => to_unsigned(482, 10), 1566 => to_unsigned(499, 10), 1567 => to_unsigned(539, 10), 1568 => to_unsigned(419, 10), 1569 => to_unsigned(459, 10), 1570 => to_unsigned(412, 10), 1571 => to_unsigned(314, 10), 1572 => to_unsigned(459, 10), 1573 => to_unsigned(654, 10), 1574 => to_unsigned(553, 10), 1575 => to_unsigned(444, 10), 1576 => to_unsigned(698, 10), 1577 => to_unsigned(629, 10), 1578 => to_unsigned(543, 10), 1579 => to_unsigned(512, 10), 1580 => to_unsigned(494, 10), 1581 => to_unsigned(383, 10), 1582 => to_unsigned(461, 10), 1583 => to_unsigned(588, 10), 1584 => to_unsigned(408, 10), 1585 => to_unsigned(664, 10), 1586 => to_unsigned(519, 10), 1587 => to_unsigned(493, 10), 1588 => to_unsigned(492, 10), 1589 => to_unsigned(574, 10), 1590 => to_unsigned(544, 10), 1591 => to_unsigned(525, 10), 1592 => to_unsigned(603, 10), 1593 => to_unsigned(669, 10), 1594 => to_unsigned(527, 10), 1595 => to_unsigned(664, 10), 1596 => to_unsigned(466, 10), 1597 => to_unsigned(590, 10), 1598 => to_unsigned(581, 10), 1599 => to_unsigned(400, 10), 1600 => to_unsigned(506, 10), 1601 => to_unsigned(501, 10), 1602 => to_unsigned(452, 10), 1603 => to_unsigned(722, 10), 1604 => to_unsigned(511, 10), 1605 => to_unsigned(379, 10), 1606 => to_unsigned(617, 10), 1607 => to_unsigned(575, 10), 1608 => to_unsigned(469, 10), 1609 => to_unsigned(388, 10), 1610 => to_unsigned(720, 10), 1611 => to_unsigned(381, 10), 1612 => to_unsigned(368, 10), 1613 => to_unsigned(562, 10), 1614 => to_unsigned(478, 10), 1615 => to_unsigned(385, 10), 1616 => to_unsigned(669, 10), 1617 => to_unsigned(495, 10), 1618 => to_unsigned(561, 10), 1619 => to_unsigned(506, 10), 1620 => to_unsigned(481, 10), 1621 => to_unsigned(503, 10), 1622 => to_unsigned(626, 10), 1623 => to_unsigned(395, 10), 1624 => to_unsigned(496, 10), 1625 => to_unsigned(498, 10), 1626 => to_unsigned(515, 10), 1627 => to_unsigned(471, 10), 1628 => to_unsigned(416, 10), 1629 => to_unsigned(515, 10), 1630 => to_unsigned(617, 10), 1631 => to_unsigned(386, 10), 1632 => to_unsigned(548, 10), 1633 => to_unsigned(700, 10), 1634 => to_unsigned(445, 10), 1635 => to_unsigned(617, 10), 1636 => to_unsigned(487, 10), 1637 => to_unsigned(671, 10), 1638 => to_unsigned(496, 10), 1639 => to_unsigned(683, 10), 1640 => to_unsigned(395, 10), 1641 => to_unsigned(418, 10), 1642 => to_unsigned(545, 10), 1643 => to_unsigned(555, 10), 1644 => to_unsigned(489, 10), 1645 => to_unsigned(531, 10), 1646 => to_unsigned(735, 10), 1647 => to_unsigned(510, 10), 1648 => to_unsigned(668, 10), 1649 => to_unsigned(580, 10), 1650 => to_unsigned(578, 10), 1651 => to_unsigned(495, 10), 1652 => to_unsigned(525, 10), 1653 => to_unsigned(533, 10), 1654 => to_unsigned(401, 10), 1655 => to_unsigned(629, 10), 1656 => to_unsigned(473, 10), 1657 => to_unsigned(355, 10), 1658 => to_unsigned(529, 10), 1659 => to_unsigned(600, 10), 1660 => to_unsigned(441, 10), 1661 => to_unsigned(574, 10), 1662 => to_unsigned(490, 10), 1663 => to_unsigned(489, 10), 1664 => to_unsigned(523, 10), 1665 => to_unsigned(596, 10), 1666 => to_unsigned(531, 10), 1667 => to_unsigned(558, 10), 1668 => to_unsigned(670, 10), 1669 => to_unsigned(509, 10), 1670 => to_unsigned(626, 10), 1671 => to_unsigned(485, 10), 1672 => to_unsigned(573, 10), 1673 => to_unsigned(343, 10), 1674 => to_unsigned(627, 10), 1675 => to_unsigned(585, 10), 1676 => to_unsigned(527, 10), 1677 => to_unsigned(688, 10), 1678 => to_unsigned(509, 10), 1679 => to_unsigned(550, 10), 1680 => to_unsigned(496, 10), 1681 => to_unsigned(481, 10), 1682 => to_unsigned(461, 10), 1683 => to_unsigned(548, 10), 1684 => to_unsigned(460, 10), 1685 => to_unsigned(451, 10), 1686 => to_unsigned(528, 10), 1687 => to_unsigned(468, 10), 1688 => to_unsigned(494, 10), 1689 => to_unsigned(520, 10), 1690 => to_unsigned(552, 10), 1691 => to_unsigned(442, 10), 1692 => to_unsigned(483, 10), 1693 => to_unsigned(508, 10), 1694 => to_unsigned(414, 10), 1695 => to_unsigned(617, 10), 1696 => to_unsigned(618, 10), 1697 => to_unsigned(385, 10), 1698 => to_unsigned(306, 10), 1699 => to_unsigned(494, 10), 1700 => to_unsigned(553, 10), 1701 => to_unsigned(490, 10), 1702 => to_unsigned(432, 10), 1703 => to_unsigned(530, 10), 1704 => to_unsigned(731, 10), 1705 => to_unsigned(572, 10), 1706 => to_unsigned(514, 10), 1707 => to_unsigned(415, 10), 1708 => to_unsigned(424, 10), 1709 => to_unsigned(531, 10), 1710 => to_unsigned(545, 10), 1711 => to_unsigned(428, 10), 1712 => to_unsigned(370, 10), 1713 => to_unsigned(447, 10), 1714 => to_unsigned(660, 10), 1715 => to_unsigned(408, 10), 1716 => to_unsigned(440, 10), 1717 => to_unsigned(369, 10), 1718 => to_unsigned(394, 10), 1719 => to_unsigned(414, 10), 1720 => to_unsigned(386, 10), 1721 => to_unsigned(463, 10), 1722 => to_unsigned(418, 10), 1723 => to_unsigned(585, 10), 1724 => to_unsigned(472, 10), 1725 => to_unsigned(358, 10), 1726 => to_unsigned(553, 10), 1727 => to_unsigned(378, 10), 1728 => to_unsigned(547, 10), 1729 => to_unsigned(555, 10), 1730 => to_unsigned(402, 10), 1731 => to_unsigned(475, 10), 1732 => to_unsigned(382, 10), 1733 => to_unsigned(367, 10), 1734 => to_unsigned(464, 10), 1735 => to_unsigned(606, 10), 1736 => to_unsigned(453, 10), 1737 => to_unsigned(446, 10), 1738 => to_unsigned(530, 10), 1739 => to_unsigned(508, 10), 1740 => to_unsigned(488, 10), 1741 => to_unsigned(471, 10), 1742 => to_unsigned(671, 10), 1743 => to_unsigned(632, 10), 1744 => to_unsigned(493, 10), 1745 => to_unsigned(469, 10), 1746 => to_unsigned(541, 10), 1747 => to_unsigned(534, 10), 1748 => to_unsigned(422, 10), 1749 => to_unsigned(592, 10), 1750 => to_unsigned(491, 10), 1751 => to_unsigned(489, 10), 1752 => to_unsigned(482, 10), 1753 => to_unsigned(370, 10), 1754 => to_unsigned(487, 10), 1755 => to_unsigned(553, 10), 1756 => to_unsigned(445, 10), 1757 => to_unsigned(642, 10), 1758 => to_unsigned(411, 10), 1759 => to_unsigned(598, 10), 1760 => to_unsigned(348, 10), 1761 => to_unsigned(448, 10), 1762 => to_unsigned(434, 10), 1763 => to_unsigned(455, 10), 1764 => to_unsigned(499, 10), 1765 => to_unsigned(594, 10), 1766 => to_unsigned(333, 10), 1767 => to_unsigned(616, 10), 1768 => to_unsigned(383, 10), 1769 => to_unsigned(674, 10), 1770 => to_unsigned(577, 10), 1771 => to_unsigned(569, 10), 1772 => to_unsigned(663, 10), 1773 => to_unsigned(636, 10), 1774 => to_unsigned(483, 10), 1775 => to_unsigned(511, 10), 1776 => to_unsigned(489, 10), 1777 => to_unsigned(573, 10), 1778 => to_unsigned(588, 10), 1779 => to_unsigned(473, 10), 1780 => to_unsigned(511, 10), 1781 => to_unsigned(404, 10), 1782 => to_unsigned(502, 10), 1783 => to_unsigned(657, 10), 1784 => to_unsigned(569, 10), 1785 => to_unsigned(719, 10), 1786 => to_unsigned(604, 10), 1787 => to_unsigned(628, 10), 1788 => to_unsigned(662, 10), 1789 => to_unsigned(352, 10), 1790 => to_unsigned(649, 10), 1791 => to_unsigned(615, 10), 1792 => to_unsigned(525, 10), 1793 => to_unsigned(429, 10), 1794 => to_unsigned(555, 10), 1795 => to_unsigned(565, 10), 1796 => to_unsigned(516, 10), 1797 => to_unsigned(524, 10), 1798 => to_unsigned(596, 10), 1799 => to_unsigned(533, 10), 1800 => to_unsigned(530, 10), 1801 => to_unsigned(460, 10), 1802 => to_unsigned(619, 10), 1803 => to_unsigned(539, 10), 1804 => to_unsigned(597, 10), 1805 => to_unsigned(555, 10), 1806 => to_unsigned(497, 10), 1807 => to_unsigned(601, 10), 1808 => to_unsigned(290, 10), 1809 => to_unsigned(443, 10), 1810 => to_unsigned(485, 10), 1811 => to_unsigned(520, 10), 1812 => to_unsigned(420, 10), 1813 => to_unsigned(445, 10), 1814 => to_unsigned(666, 10), 1815 => to_unsigned(401, 10), 1816 => to_unsigned(411, 10), 1817 => to_unsigned(489, 10), 1818 => to_unsigned(604, 10), 1819 => to_unsigned(624, 10), 1820 => to_unsigned(545, 10), 1821 => to_unsigned(424, 10), 1822 => to_unsigned(605, 10), 1823 => to_unsigned(481, 10), 1824 => to_unsigned(345, 10), 1825 => to_unsigned(541, 10), 1826 => to_unsigned(385, 10), 1827 => to_unsigned(416, 10), 1828 => to_unsigned(360, 10), 1829 => to_unsigned(654, 10), 1830 => to_unsigned(561, 10), 1831 => to_unsigned(603, 10), 1832 => to_unsigned(548, 10), 1833 => to_unsigned(625, 10), 1834 => to_unsigned(428, 10), 1835 => to_unsigned(479, 10), 1836 => to_unsigned(501, 10), 1837 => to_unsigned(430, 10), 1838 => to_unsigned(456, 10), 1839 => to_unsigned(596, 10), 1840 => to_unsigned(510, 10), 1841 => to_unsigned(469, 10), 1842 => to_unsigned(404, 10), 1843 => to_unsigned(406, 10), 1844 => to_unsigned(569, 10), 1845 => to_unsigned(460, 10), 1846 => to_unsigned(401, 10), 1847 => to_unsigned(475, 10), 1848 => to_unsigned(503, 10), 1849 => to_unsigned(482, 10), 1850 => to_unsigned(623, 10), 1851 => to_unsigned(575, 10), 1852 => to_unsigned(568, 10), 1853 => to_unsigned(551, 10), 1854 => to_unsigned(498, 10), 1855 => to_unsigned(534, 10), 1856 => to_unsigned(423, 10), 1857 => to_unsigned(546, 10), 1858 => to_unsigned(508, 10), 1859 => to_unsigned(330, 10), 1860 => to_unsigned(666, 10), 1861 => to_unsigned(489, 10), 1862 => to_unsigned(476, 10), 1863 => to_unsigned(548, 10), 1864 => to_unsigned(662, 10), 1865 => to_unsigned(397, 10), 1866 => to_unsigned(650, 10), 1867 => to_unsigned(588, 10), 1868 => to_unsigned(619, 10), 1869 => to_unsigned(490, 10), 1870 => to_unsigned(389, 10), 1871 => to_unsigned(631, 10), 1872 => to_unsigned(533, 10), 1873 => to_unsigned(527, 10), 1874 => to_unsigned(638, 10), 1875 => to_unsigned(431, 10), 1876 => to_unsigned(642, 10), 1877 => to_unsigned(502, 10), 1878 => to_unsigned(518, 10), 1879 => to_unsigned(447, 10), 1880 => to_unsigned(385, 10), 1881 => to_unsigned(456, 10), 1882 => to_unsigned(574, 10), 1883 => to_unsigned(656, 10), 1884 => to_unsigned(549, 10), 1885 => to_unsigned(635, 10), 1886 => to_unsigned(427, 10), 1887 => to_unsigned(437, 10), 1888 => to_unsigned(451, 10), 1889 => to_unsigned(438, 10), 1890 => to_unsigned(464, 10), 1891 => to_unsigned(576, 10), 1892 => to_unsigned(642, 10), 1893 => to_unsigned(457, 10), 1894 => to_unsigned(419, 10), 1895 => to_unsigned(683, 10), 1896 => to_unsigned(471, 10), 1897 => to_unsigned(612, 10), 1898 => to_unsigned(590, 10), 1899 => to_unsigned(554, 10), 1900 => to_unsigned(563, 10), 1901 => to_unsigned(476, 10), 1902 => to_unsigned(540, 10), 1903 => to_unsigned(508, 10), 1904 => to_unsigned(590, 10), 1905 => to_unsigned(498, 10), 1906 => to_unsigned(570, 10), 1907 => to_unsigned(504, 10), 1908 => to_unsigned(479, 10), 1909 => to_unsigned(556, 10), 1910 => to_unsigned(512, 10), 1911 => to_unsigned(620, 10), 1912 => to_unsigned(506, 10), 1913 => to_unsigned(440, 10), 1914 => to_unsigned(553, 10), 1915 => to_unsigned(735, 10), 1916 => to_unsigned(495, 10), 1917 => to_unsigned(588, 10), 1918 => to_unsigned(593, 10), 1919 => to_unsigned(650, 10), 1920 => to_unsigned(521, 10), 1921 => to_unsigned(392, 10), 1922 => to_unsigned(537, 10), 1923 => to_unsigned(631, 10), 1924 => to_unsigned(520, 10), 1925 => to_unsigned(405, 10), 1926 => to_unsigned(444, 10), 1927 => to_unsigned(660, 10), 1928 => to_unsigned(680, 10), 1929 => to_unsigned(650, 10), 1930 => to_unsigned(519, 10), 1931 => to_unsigned(674, 10), 1932 => to_unsigned(505, 10), 1933 => to_unsigned(609, 10), 1934 => to_unsigned(463, 10), 1935 => to_unsigned(549, 10), 1936 => to_unsigned(451, 10), 1937 => to_unsigned(769, 10), 1938 => to_unsigned(363, 10), 1939 => to_unsigned(558, 10), 1940 => to_unsigned(524, 10), 1941 => to_unsigned(485, 10), 1942 => to_unsigned(521, 10), 1943 => to_unsigned(720, 10), 1944 => to_unsigned(364, 10), 1945 => to_unsigned(654, 10), 1946 => to_unsigned(468, 10), 1947 => to_unsigned(590, 10), 1948 => to_unsigned(528, 10), 1949 => to_unsigned(526, 10), 1950 => to_unsigned(543, 10), 1951 => to_unsigned(513, 10), 1952 => to_unsigned(598, 10), 1953 => to_unsigned(332, 10), 1954 => to_unsigned(493, 10), 1955 => to_unsigned(567, 10), 1956 => to_unsigned(597, 10), 1957 => to_unsigned(542, 10), 1958 => to_unsigned(336, 10), 1959 => to_unsigned(694, 10), 1960 => to_unsigned(588, 10), 1961 => to_unsigned(406, 10), 1962 => to_unsigned(415, 10), 1963 => to_unsigned(536, 10), 1964 => to_unsigned(437, 10), 1965 => to_unsigned(484, 10), 1966 => to_unsigned(364, 10), 1967 => to_unsigned(367, 10), 1968 => to_unsigned(431, 10), 1969 => to_unsigned(778, 10), 1970 => to_unsigned(575, 10), 1971 => to_unsigned(548, 10), 1972 => to_unsigned(613, 10), 1973 => to_unsigned(534, 10), 1974 => to_unsigned(323, 10), 1975 => to_unsigned(290, 10), 1976 => to_unsigned(345, 10), 1977 => to_unsigned(564, 10), 1978 => to_unsigned(516, 10), 1979 => to_unsigned(489, 10), 1980 => to_unsigned(484, 10), 1981 => to_unsigned(433, 10), 1982 => to_unsigned(560, 10), 1983 => to_unsigned(472, 10), 1984 => to_unsigned(474, 10), 1985 => to_unsigned(557, 10), 1986 => to_unsigned(657, 10), 1987 => to_unsigned(439, 10), 1988 => to_unsigned(553, 10), 1989 => to_unsigned(444, 10), 1990 => to_unsigned(640, 10), 1991 => to_unsigned(598, 10), 1992 => to_unsigned(628, 10), 1993 => to_unsigned(595, 10), 1994 => to_unsigned(635, 10), 1995 => to_unsigned(557, 10), 1996 => to_unsigned(565, 10), 1997 => to_unsigned(577, 10), 1998 => to_unsigned(573, 10), 1999 => to_unsigned(571, 10), 2000 => to_unsigned(510, 10), 2001 => to_unsigned(529, 10), 2002 => to_unsigned(302, 10), 2003 => to_unsigned(509, 10), 2004 => to_unsigned(508, 10), 2005 => to_unsigned(527, 10), 2006 => to_unsigned(729, 10), 2007 => to_unsigned(508, 10), 2008 => to_unsigned(579, 10), 2009 => to_unsigned(477, 10), 2010 => to_unsigned(594, 10), 2011 => to_unsigned(354, 10), 2012 => to_unsigned(229, 10), 2013 => to_unsigned(790, 10), 2014 => to_unsigned(401, 10), 2015 => to_unsigned(469, 10), 2016 => to_unsigned(521, 10), 2017 => to_unsigned(657, 10), 2018 => to_unsigned(353, 10), 2019 => to_unsigned(397, 10), 2020 => to_unsigned(519, 10), 2021 => to_unsigned(502, 10), 2022 => to_unsigned(538, 10), 2023 => to_unsigned(543, 10), 2024 => to_unsigned(479, 10), 2025 => to_unsigned(487, 10), 2026 => to_unsigned(384, 10), 2027 => to_unsigned(680, 10), 2028 => to_unsigned(473, 10), 2029 => to_unsigned(597, 10), 2030 => to_unsigned(386, 10), 2031 => to_unsigned(386, 10), 2032 => to_unsigned(415, 10), 2033 => to_unsigned(533, 10), 2034 => to_unsigned(539, 10), 2035 => to_unsigned(553, 10), 2036 => to_unsigned(625, 10), 2037 => to_unsigned(489, 10), 2038 => to_unsigned(541, 10), 2039 => to_unsigned(512, 10), 2040 => to_unsigned(521, 10), 2041 => to_unsigned(414, 10), 2042 => to_unsigned(578, 10), 2043 => to_unsigned(422, 10), 2044 => to_unsigned(581, 10), 2045 => to_unsigned(438, 10), 2046 => to_unsigned(402, 10), 2047 => to_unsigned(430, 10))
    );

begin

	-- Generate main clock signal
    clock_gen : process
        constant clock_period : time := 20 ns;
	begin
		wait for clock_period / 2;
		clock <= not clock;
	end process clock_gen;

    test : process
        constant fragment_size : integer := vnir_row_width / vnir_lvds_data_width;
        variable tests_passed : boolean := true;
    begin
        reset_n <= '0';
        wait until rising_edge(clock);
        reset_n <= '1';

        config.window_blue <= (lo => window_size * 0, hi => window_size * 1 - 1);
        config.window_red  <= (lo => window_size * 1, hi => window_size * 2 - 1);
        config.window_nir  <= (lo => window_size * 2, hi => window_size * 3 - 1);
        read_config <= '1';
        wait until rising_edge(clock);
        read_config <= '0';

        report "Uploading started";
        pixels_available <= '1';
        for color in 0 to n_colours-1 loop
            for row in 0 to window_size-1 loop
                for fragment in 0 to fragment_size-1 loop
                    for i in 0 to vnir_lvds_data_width-1 loop
                        pixels(i) <= data(color)(row)(fragment + fragment_size * i);
                    end loop;
                    wait until rising_edge(clock);
                end loop;
            end loop;
        end loop;
        pixels_available <= '0';
        report "Uploading finished";
        
        wait until rising_edge(clock);
        tests_passed := tests_passed and test_report(rows_available = '1', "rows available");
        tests_passed := tests_passed and test_report(rows.red = averages(0), "red row");
        tests_passed := tests_passed and test_report(rows.blue = averages(1), "blue row");
        tests_passed := tests_passed and test_report(rows.nir = averages(2), "NIR row");

        test_end(tests_passed);
        wait;
    end process test;

    row_collator_component : row_collator port map (
        clock => clock,
        reset_n => reset_n,
        config => config,
        read_config => read_config,
        pixels => pixels,
        pixels_available => pixels_available,
        rows => rows,
        rows_available => rows_available
    );

end tests;
