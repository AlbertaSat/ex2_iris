----------------------------------------------------------------
-- Copyright 2020 University of Alberta

-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at

--     http://www.apache.org/licenses/LICENSE-2.0

-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
----------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.spi_types.all;
use work.vnir_types.all;
use work.test_util.all;

use work.row_collector_pkg.all;


entity row_collector_tb is
end entity row_collector_tb;

architecture tests of row_collector_tb is
	signal clock                : std_logic := '0';
	signal config               : vnir_config_t;
    signal read_config          : std_logic := '0';
    signal start                : std_logic := '0';
    signal fragment             : fragment_t;
	signal fragment_available   : std_logic := '0';
	signal rows                 : vnir_rows_t;
	signal rows_available       : std_logic := '0';

    component row_collector is
    port (
        clock               : in std_logic;
        config              : in vnir_config_t;
        read_config         : in std_logic;
        start               : in std_logic;
        fragment            : in fragment_t;
        fragment_available  : in std_logic;
        rows                : out vnir_rows_t;
        rows_available      : out std_logic
    );
    end component row_collector;

    type vnir_row_vector_t is array(integer range <>) of vnir_row_t;
    
    constant data : vnir_row_vector_t(2 downto 0) := (
        0 => (0 => to_unsigned(684, 10), 1 => to_unsigned(559, 10), 2 => to_unsigned(629, 10), 3 => to_unsigned(192, 10), 4 => to_unsigned(835, 10), 5 => to_unsigned(763, 10), 6 => to_unsigned(707, 10), 7 => to_unsigned(359, 10), 8 => to_unsigned(9, 10), 9 => to_unsigned(723, 10), 10 => to_unsigned(277, 10), 11 => to_unsigned(754, 10), 12 => to_unsigned(804, 10), 13 => to_unsigned(599, 10), 14 => to_unsigned(70, 10), 15 => to_unsigned(472, 10), 16 => to_unsigned(600, 10), 17 => to_unsigned(396, 10), 18 => to_unsigned(314, 10), 19 => to_unsigned(705, 10), 20 => to_unsigned(486, 10), 21 => to_unsigned(551, 10), 22 => to_unsigned(87, 10), 23 => to_unsigned(174, 10), 24 => to_unsigned(600, 10), 25 => to_unsigned(849, 10), 26 => to_unsigned(677, 10), 27 => to_unsigned(537, 10), 28 => to_unsigned(845, 10), 29 => to_unsigned(72, 10), 30 => to_unsigned(777, 10), 31 => to_unsigned(916, 10), 32 => to_unsigned(115, 10), 33 => to_unsigned(976, 10), 34 => to_unsigned(755, 10), 35 => to_unsigned(709, 10), 36 => to_unsigned(1022, 10), 37 => to_unsigned(847, 10), 38 => to_unsigned(431, 10), 39 => to_unsigned(448, 10), 40 => to_unsigned(850, 10), 41 => to_unsigned(99, 10), 42 => to_unsigned(984, 10), 43 => to_unsigned(177, 10), 44 => to_unsigned(755, 10), 45 => to_unsigned(797, 10), 46 => to_unsigned(659, 10), 47 => to_unsigned(147, 10), 48 => to_unsigned(910, 10), 49 => to_unsigned(423, 10), 50 => to_unsigned(288, 10), 51 => to_unsigned(961, 10), 52 => to_unsigned(265, 10), 53 => to_unsigned(697, 10), 54 => to_unsigned(639, 10), 55 => to_unsigned(544, 10), 56 => to_unsigned(543, 10), 57 => to_unsigned(714, 10), 58 => to_unsigned(244, 10), 59 => to_unsigned(151, 10), 60 => to_unsigned(675, 10), 61 => to_unsigned(510, 10), 62 => to_unsigned(459, 10), 63 => to_unsigned(882, 10), 64 => to_unsigned(183, 10), 65 => to_unsigned(28, 10), 66 => to_unsigned(802, 10), 67 => to_unsigned(128, 10), 68 => to_unsigned(128, 10), 69 => to_unsigned(932, 10), 70 => to_unsigned(53, 10), 71 => to_unsigned(901, 10), 72 => to_unsigned(550, 10), 73 => to_unsigned(488, 10), 74 => to_unsigned(756, 10), 75 => to_unsigned(273, 10), 76 => to_unsigned(335, 10), 77 => to_unsigned(388, 10), 78 => to_unsigned(617, 10), 79 => to_unsigned(42, 10), 80 => to_unsigned(442, 10), 81 => to_unsigned(543, 10), 82 => to_unsigned(888, 10), 83 => to_unsigned(257, 10), 84 => to_unsigned(321, 10), 85 => to_unsigned(999, 10), 86 => to_unsigned(937, 10), 87 => to_unsigned(57, 10), 88 => to_unsigned(291, 10), 89 => to_unsigned(870, 10), 90 => to_unsigned(119, 10), 91 => to_unsigned(779, 10), 92 => to_unsigned(430, 10), 93 => to_unsigned(82, 10), 94 => to_unsigned(91, 10), 95 => to_unsigned(896, 10), 96 => to_unsigned(398, 10), 97 => to_unsigned(611, 10), 98 => to_unsigned(565, 10), 99 => to_unsigned(908, 10), 100 => to_unsigned(633, 10), 101 => to_unsigned(938, 10), 102 => to_unsigned(84, 10), 103 => to_unsigned(203, 10), 104 => to_unsigned(324, 10), 105 => to_unsigned(774, 10), 106 => to_unsigned(964, 10), 107 => to_unsigned(47, 10), 108 => to_unsigned(639, 10), 109 => to_unsigned(1012, 10), 110 => to_unsigned(131, 10), 111 => to_unsigned(972, 10), 112 => to_unsigned(868, 10), 113 => to_unsigned(180, 10), 114 => to_unsigned(1000, 10), 115 => to_unsigned(846, 10), 116 => to_unsigned(143, 10), 117 => to_unsigned(660, 10), 118 => to_unsigned(227, 10), 119 => to_unsigned(954, 10), 120 => to_unsigned(791, 10), 121 => to_unsigned(719, 10), 122 => to_unsigned(909, 10), 123 => to_unsigned(373, 10), 124 => to_unsigned(853, 10), 125 => to_unsigned(560, 10), 126 => to_unsigned(305, 10), 127 => to_unsigned(581, 10), 128 => to_unsigned(169, 10), 129 => to_unsigned(675, 10), 130 => to_unsigned(448, 10), 131 => to_unsigned(95, 10), 132 => to_unsigned(197, 10), 133 => to_unsigned(606, 10), 134 => to_unsigned(256, 10), 135 => to_unsigned(881, 10), 136 => to_unsigned(690, 10), 137 => to_unsigned(292, 10), 138 => to_unsigned(930, 10), 139 => to_unsigned(816, 10), 140 => to_unsigned(861, 10), 141 => to_unsigned(387, 10), 142 => to_unsigned(610, 10), 143 => to_unsigned(554, 10), 144 => to_unsigned(973, 10), 145 => to_unsigned(368, 10), 146 => to_unsigned(999, 10), 147 => to_unsigned(917, 10), 148 => to_unsigned(201, 10), 149 => to_unsigned(383, 10), 150 => to_unsigned(512, 10), 151 => to_unsigned(906, 10), 152 => to_unsigned(370, 10), 153 => to_unsigned(555, 10), 154 => to_unsigned(954, 10), 155 => to_unsigned(383, 10), 156 => to_unsigned(23, 10), 157 => to_unsigned(699, 10), 158 => to_unsigned(130, 10), 159 => to_unsigned(377, 10), 160 => to_unsigned(98, 10), 161 => to_unsigned(574, 10), 162 => to_unsigned(931, 10), 163 => to_unsigned(734, 10), 164 => to_unsigned(123, 10), 165 => to_unsigned(963, 10), 166 => to_unsigned(594, 10), 167 => to_unsigned(942, 10), 168 => to_unsigned(739, 10), 169 => to_unsigned(148, 10), 170 => to_unsigned(209, 10), 171 => to_unsigned(562, 10), 172 => to_unsigned(411, 10), 173 => to_unsigned(782, 10), 174 => to_unsigned(41, 10), 175 => to_unsigned(58, 10), 176 => to_unsigned(705, 10), 177 => to_unsigned(36, 10), 178 => to_unsigned(778, 10), 179 => to_unsigned(86, 10), 180 => to_unsigned(43, 10), 181 => to_unsigned(872, 10), 182 => to_unsigned(11, 10), 183 => to_unsigned(770, 10), 184 => to_unsigned(307, 10), 185 => to_unsigned(80, 10), 186 => to_unsigned(32, 10), 187 => to_unsigned(182, 10), 188 => to_unsigned(128, 10), 189 => to_unsigned(806, 10), 190 => to_unsigned(275, 10), 191 => to_unsigned(174, 10), 192 => to_unsigned(554, 10), 193 => to_unsigned(371, 10), 194 => to_unsigned(184, 10), 195 => to_unsigned(444, 10), 196 => to_unsigned(488, 10), 197 => to_unsigned(589, 10), 198 => to_unsigned(286, 10), 199 => to_unsigned(280, 10), 200 => to_unsigned(637, 10), 201 => to_unsigned(770, 10), 202 => to_unsigned(515, 10), 203 => to_unsigned(94, 10), 204 => to_unsigned(226, 10), 205 => to_unsigned(875, 10), 206 => to_unsigned(269, 10), 207 => to_unsigned(880, 10), 208 => to_unsigned(296, 10), 209 => to_unsigned(328, 10), 210 => to_unsigned(19, 10), 211 => to_unsigned(607, 10), 212 => to_unsigned(840, 10), 213 => to_unsigned(410, 10), 214 => to_unsigned(450, 10), 215 => to_unsigned(248, 10), 216 => to_unsigned(180, 10), 217 => to_unsigned(323, 10), 218 => to_unsigned(1004, 10), 219 => to_unsigned(829, 10), 220 => to_unsigned(782, 10), 221 => to_unsigned(864, 10), 222 => to_unsigned(260, 10), 223 => to_unsigned(963, 10), 224 => to_unsigned(749, 10), 225 => to_unsigned(139, 10), 226 => to_unsigned(1020, 10), 227 => to_unsigned(598, 10), 228 => to_unsigned(461, 10), 229 => to_unsigned(889, 10), 230 => to_unsigned(621, 10), 231 => to_unsigned(843, 10), 232 => to_unsigned(696, 10), 233 => to_unsigned(528, 10), 234 => to_unsigned(152, 10), 235 => to_unsigned(925, 10), 236 => to_unsigned(149, 10), 237 => to_unsigned(110, 10), 238 => to_unsigned(25, 10), 239 => to_unsigned(464, 10), 240 => to_unsigned(956, 10), 241 => to_unsigned(889, 10), 242 => to_unsigned(886, 10), 243 => to_unsigned(117, 10), 244 => to_unsigned(445, 10), 245 => to_unsigned(595, 10), 246 => to_unsigned(673, 10), 247 => to_unsigned(872, 10), 248 => to_unsigned(928, 10), 249 => to_unsigned(228, 10), 250 => to_unsigned(507, 10), 251 => to_unsigned(763, 10), 252 => to_unsigned(121, 10), 253 => to_unsigned(326, 10), 254 => to_unsigned(469, 10), 255 => to_unsigned(287, 10), 256 => to_unsigned(525, 10), 257 => to_unsigned(839, 10), 258 => to_unsigned(696, 10), 259 => to_unsigned(152, 10), 260 => to_unsigned(591, 10), 261 => to_unsigned(41, 10), 262 => to_unsigned(274, 10), 263 => to_unsigned(552, 10), 264 => to_unsigned(438, 10), 265 => to_unsigned(207, 10), 266 => to_unsigned(779, 10), 267 => to_unsigned(166, 10), 268 => to_unsigned(111, 10), 269 => to_unsigned(349, 10), 270 => to_unsigned(1017, 10), 271 => to_unsigned(129, 10), 272 => to_unsigned(735, 10), 273 => to_unsigned(886, 10), 274 => to_unsigned(812, 10), 275 => to_unsigned(216, 10), 276 => to_unsigned(381, 10), 277 => to_unsigned(24, 10), 278 => to_unsigned(67, 10), 279 => to_unsigned(978, 10), 280 => to_unsigned(1007, 10), 281 => to_unsigned(771, 10), 282 => to_unsigned(234, 10), 283 => to_unsigned(716, 10), 284 => to_unsigned(998, 10), 285 => to_unsigned(291, 10), 286 => to_unsigned(726, 10), 287 => to_unsigned(1022, 10), 288 => to_unsigned(701, 10), 289 => to_unsigned(709, 10), 290 => to_unsigned(727, 10), 291 => to_unsigned(555, 10), 292 => to_unsigned(32, 10), 293 => to_unsigned(11, 10), 294 => to_unsigned(616, 10), 295 => to_unsigned(212, 10), 296 => to_unsigned(138, 10), 297 => to_unsigned(694, 10), 298 => to_unsigned(1003, 10), 299 => to_unsigned(421, 10), 300 => to_unsigned(637, 10), 301 => to_unsigned(668, 10), 302 => to_unsigned(623, 10), 303 => to_unsigned(488, 10), 304 => to_unsigned(770, 10), 305 => to_unsigned(539, 10), 306 => to_unsigned(979, 10), 307 => to_unsigned(217, 10), 308 => to_unsigned(663, 10), 309 => to_unsigned(821, 10), 310 => to_unsigned(307, 10), 311 => to_unsigned(174, 10), 312 => to_unsigned(148, 10), 313 => to_unsigned(949, 10), 314 => to_unsigned(541, 10), 315 => to_unsigned(579, 10), 316 => to_unsigned(547, 10), 317 => to_unsigned(807, 10), 318 => to_unsigned(393, 10), 319 => to_unsigned(73, 10), 320 => to_unsigned(297, 10), 321 => to_unsigned(919, 10), 322 => to_unsigned(899, 10), 323 => to_unsigned(814, 10), 324 => to_unsigned(730, 10), 325 => to_unsigned(946, 10), 326 => to_unsigned(876, 10), 327 => to_unsigned(771, 10), 328 => to_unsigned(799, 10), 329 => to_unsigned(777, 10), 330 => to_unsigned(394, 10), 331 => to_unsigned(539, 10), 332 => to_unsigned(429, 10), 333 => to_unsigned(199, 10), 334 => to_unsigned(423, 10), 335 => to_unsigned(61, 10), 336 => to_unsigned(341, 10), 337 => to_unsigned(865, 10), 338 => to_unsigned(44, 10), 339 => to_unsigned(802, 10), 340 => to_unsigned(930, 10), 341 => to_unsigned(88, 10), 342 => to_unsigned(33, 10), 343 => to_unsigned(645, 10), 344 => to_unsigned(232, 10), 345 => to_unsigned(767, 10), 346 => to_unsigned(36, 10), 347 => to_unsigned(768, 10), 348 => to_unsigned(459, 10), 349 => to_unsigned(290, 10), 350 => to_unsigned(197, 10), 351 => to_unsigned(894, 10), 352 => to_unsigned(949, 10), 353 => to_unsigned(254, 10), 354 => to_unsigned(80, 10), 355 => to_unsigned(446, 10), 356 => to_unsigned(136, 10), 357 => to_unsigned(189, 10), 358 => to_unsigned(129, 10), 359 => to_unsigned(209, 10), 360 => to_unsigned(368, 10), 361 => to_unsigned(291, 10), 362 => to_unsigned(376, 10), 363 => to_unsigned(347, 10), 364 => to_unsigned(168, 10), 365 => to_unsigned(884, 10), 366 => to_unsigned(804, 10), 367 => to_unsigned(176, 10), 368 => to_unsigned(537, 10), 369 => to_unsigned(323, 10), 370 => to_unsigned(871, 10), 371 => to_unsigned(508, 10), 372 => to_unsigned(803, 10), 373 => to_unsigned(114, 10), 374 => to_unsigned(798, 10), 375 => to_unsigned(29, 10), 376 => to_unsigned(753, 10), 377 => to_unsigned(289, 10), 378 => to_unsigned(146, 10), 379 => to_unsigned(273, 10), 380 => to_unsigned(221, 10), 381 => to_unsigned(340, 10), 382 => to_unsigned(509, 10), 383 => to_unsigned(514, 10), 384 => to_unsigned(69, 10), 385 => to_unsigned(357, 10), 386 => to_unsigned(908, 10), 387 => to_unsigned(556, 10), 388 => to_unsigned(885, 10), 389 => to_unsigned(765, 10), 390 => to_unsigned(322, 10), 391 => to_unsigned(623, 10), 392 => to_unsigned(91, 10), 393 => to_unsigned(341, 10), 394 => to_unsigned(423, 10), 395 => to_unsigned(551, 10), 396 => to_unsigned(971, 10), 397 => to_unsigned(662, 10), 398 => to_unsigned(414, 10), 399 => to_unsigned(657, 10), 400 => to_unsigned(710, 10), 401 => to_unsigned(967, 10), 402 => to_unsigned(274, 10), 403 => to_unsigned(860, 10), 404 => to_unsigned(43, 10), 405 => to_unsigned(83, 10), 406 => to_unsigned(433, 10), 407 => to_unsigned(809, 10), 408 => to_unsigned(93, 10), 409 => to_unsigned(174, 10), 410 => to_unsigned(405, 10), 411 => to_unsigned(201, 10), 412 => to_unsigned(857, 10), 413 => to_unsigned(498, 10), 414 => to_unsigned(480, 10), 415 => to_unsigned(987, 10), 416 => to_unsigned(329, 10), 417 => to_unsigned(540, 10), 418 => to_unsigned(1003, 10), 419 => to_unsigned(209, 10), 420 => to_unsigned(617, 10), 421 => to_unsigned(954, 10), 422 => to_unsigned(896, 10), 423 => to_unsigned(982, 10), 424 => to_unsigned(575, 10), 425 => to_unsigned(16, 10), 426 => to_unsigned(106, 10), 427 => to_unsigned(164, 10), 428 => to_unsigned(606, 10), 429 => to_unsigned(536, 10), 430 => to_unsigned(628, 10), 431 => to_unsigned(191, 10), 432 => to_unsigned(195, 10), 433 => to_unsigned(307, 10), 434 => to_unsigned(136, 10), 435 => to_unsigned(952, 10), 436 => to_unsigned(859, 10), 437 => to_unsigned(93, 10), 438 => to_unsigned(891, 10), 439 => to_unsigned(750, 10), 440 => to_unsigned(87, 10), 441 => to_unsigned(160, 10), 442 => to_unsigned(147, 10), 443 => to_unsigned(584, 10), 444 => to_unsigned(455, 10), 445 => to_unsigned(87, 10), 446 => to_unsigned(13, 10), 447 => to_unsigned(314, 10), 448 => to_unsigned(593, 10), 449 => to_unsigned(120, 10), 450 => to_unsigned(884, 10), 451 => to_unsigned(951, 10), 452 => to_unsigned(832, 10), 453 => to_unsigned(715, 10), 454 => to_unsigned(732, 10), 455 => to_unsigned(932, 10), 456 => to_unsigned(281, 10), 457 => to_unsigned(800, 10), 458 => to_unsigned(426, 10), 459 => to_unsigned(782, 10), 460 => to_unsigned(470, 10), 461 => to_unsigned(284, 10), 462 => to_unsigned(276, 10), 463 => to_unsigned(978, 10), 464 => to_unsigned(324, 10), 465 => to_unsigned(534, 10), 466 => to_unsigned(227, 10), 467 => to_unsigned(890, 10), 468 => to_unsigned(595, 10), 469 => to_unsigned(647, 10), 470 => to_unsigned(968, 10), 471 => to_unsigned(573, 10), 472 => to_unsigned(653, 10), 473 => to_unsigned(517, 10), 474 => to_unsigned(256, 10), 475 => to_unsigned(136, 10), 476 => to_unsigned(207, 10), 477 => to_unsigned(463, 10), 478 => to_unsigned(949, 10), 479 => to_unsigned(139, 10), 480 => to_unsigned(4, 10), 481 => to_unsigned(423, 10), 482 => to_unsigned(348, 10), 483 => to_unsigned(941, 10), 484 => to_unsigned(282, 10), 485 => to_unsigned(586, 10), 486 => to_unsigned(820, 10), 487 => to_unsigned(1006, 10), 488 => to_unsigned(433, 10), 489 => to_unsigned(219, 10), 490 => to_unsigned(819, 10), 491 => to_unsigned(739, 10), 492 => to_unsigned(873, 10), 493 => to_unsigned(786, 10), 494 => to_unsigned(373, 10), 495 => to_unsigned(290, 10), 496 => to_unsigned(563, 10), 497 => to_unsigned(670, 10), 498 => to_unsigned(437, 10), 499 => to_unsigned(826, 10), 500 => to_unsigned(939, 10), 501 => to_unsigned(823, 10), 502 => to_unsigned(508, 10), 503 => to_unsigned(1020, 10), 504 => to_unsigned(786, 10), 505 => to_unsigned(941, 10), 506 => to_unsigned(855, 10), 507 => to_unsigned(449, 10), 508 => to_unsigned(326, 10), 509 => to_unsigned(490, 10), 510 => to_unsigned(53, 10), 511 => to_unsigned(816, 10), 512 => to_unsigned(94, 10), 513 => to_unsigned(59, 10), 514 => to_unsigned(336, 10), 515 => to_unsigned(666, 10), 516 => to_unsigned(636, 10), 517 => to_unsigned(163, 10), 518 => to_unsigned(570, 10), 519 => to_unsigned(945, 10), 520 => to_unsigned(106, 10), 521 => to_unsigned(201, 10), 522 => to_unsigned(300, 10), 523 => to_unsigned(781, 10), 524 => to_unsigned(889, 10), 525 => to_unsigned(838, 10), 526 => to_unsigned(550, 10), 527 => to_unsigned(679, 10), 528 => to_unsigned(648, 10), 529 => to_unsigned(13, 10), 530 => to_unsigned(1016, 10), 531 => to_unsigned(903, 10), 532 => to_unsigned(720, 10), 533 => to_unsigned(1016, 10), 534 => to_unsigned(534, 10), 535 => to_unsigned(504, 10), 536 => to_unsigned(847, 10), 537 => to_unsigned(985, 10), 538 => to_unsigned(776, 10), 539 => to_unsigned(739, 10), 540 => to_unsigned(774, 10), 541 => to_unsigned(209, 10), 542 => to_unsigned(455, 10), 543 => to_unsigned(468, 10), 544 => to_unsigned(473, 10), 545 => to_unsigned(962, 10), 546 => to_unsigned(572, 10), 547 => to_unsigned(400, 10), 548 => to_unsigned(56, 10), 549 => to_unsigned(882, 10), 550 => to_unsigned(749, 10), 551 => to_unsigned(663, 10), 552 => to_unsigned(280, 10), 553 => to_unsigned(4, 10), 554 => to_unsigned(612, 10), 555 => to_unsigned(1004, 10), 556 => to_unsigned(305, 10), 557 => to_unsigned(343, 10), 558 => to_unsigned(542, 10), 559 => to_unsigned(566, 10), 560 => to_unsigned(153, 10), 561 => to_unsigned(788, 10), 562 => to_unsigned(353, 10), 563 => to_unsigned(357, 10), 564 => to_unsigned(697, 10), 565 => to_unsigned(407, 10), 566 => to_unsigned(411, 10), 567 => to_unsigned(29, 10), 568 => to_unsigned(929, 10), 569 => to_unsigned(371, 10), 570 => to_unsigned(821, 10), 571 => to_unsigned(631, 10), 572 => to_unsigned(947, 10), 573 => to_unsigned(854, 10), 574 => to_unsigned(502, 10), 575 => to_unsigned(7, 10), 576 => to_unsigned(617, 10), 577 => to_unsigned(1009, 10), 578 => to_unsigned(137, 10), 579 => to_unsigned(694, 10), 580 => to_unsigned(896, 10), 581 => to_unsigned(851, 10), 582 => to_unsigned(376, 10), 583 => to_unsigned(932, 10), 584 => to_unsigned(721, 10), 585 => to_unsigned(148, 10), 586 => to_unsigned(885, 10), 587 => to_unsigned(1008, 10), 588 => to_unsigned(259, 10), 589 => to_unsigned(126, 10), 590 => to_unsigned(810, 10), 591 => to_unsigned(577, 10), 592 => to_unsigned(532, 10), 593 => to_unsigned(804, 10), 594 => to_unsigned(324, 10), 595 => to_unsigned(976, 10), 596 => to_unsigned(112, 10), 597 => to_unsigned(943, 10), 598 => to_unsigned(650, 10), 599 => to_unsigned(237, 10), 600 => to_unsigned(360, 10), 601 => to_unsigned(990, 10), 602 => to_unsigned(859, 10), 603 => to_unsigned(555, 10), 604 => to_unsigned(63, 10), 605 => to_unsigned(927, 10), 606 => to_unsigned(916, 10), 607 => to_unsigned(454, 10), 608 => to_unsigned(265, 10), 609 => to_unsigned(444, 10), 610 => to_unsigned(603, 10), 611 => to_unsigned(623, 10), 612 => to_unsigned(419, 10), 613 => to_unsigned(339, 10), 614 => to_unsigned(844, 10), 615 => to_unsigned(274, 10), 616 => to_unsigned(369, 10), 617 => to_unsigned(842, 10), 618 => to_unsigned(226, 10), 619 => to_unsigned(225, 10), 620 => to_unsigned(939, 10), 621 => to_unsigned(643, 10), 622 => to_unsigned(908, 10), 623 => to_unsigned(228, 10), 624 => to_unsigned(826, 10), 625 => to_unsigned(897, 10), 626 => to_unsigned(369, 10), 627 => to_unsigned(128, 10), 628 => to_unsigned(807, 10), 629 => to_unsigned(24, 10), 630 => to_unsigned(698, 10), 631 => to_unsigned(292, 10), 632 => to_unsigned(355, 10), 633 => to_unsigned(837, 10), 634 => to_unsigned(134, 10), 635 => to_unsigned(3, 10), 636 => to_unsigned(226, 10), 637 => to_unsigned(889, 10), 638 => to_unsigned(680, 10), 639 => to_unsigned(444, 10), 640 => to_unsigned(417, 10), 641 => to_unsigned(284, 10), 642 => to_unsigned(836, 10), 643 => to_unsigned(26, 10), 644 => to_unsigned(736, 10), 645 => to_unsigned(248, 10), 646 => to_unsigned(365, 10), 647 => to_unsigned(947, 10), 648 => to_unsigned(201, 10), 649 => to_unsigned(437, 10), 650 => to_unsigned(197, 10), 651 => to_unsigned(929, 10), 652 => to_unsigned(647, 10), 653 => to_unsigned(637, 10), 654 => to_unsigned(606, 10), 655 => to_unsigned(72, 10), 656 => to_unsigned(246, 10), 657 => to_unsigned(852, 10), 658 => to_unsigned(135, 10), 659 => to_unsigned(707, 10), 660 => to_unsigned(213, 10), 661 => to_unsigned(475, 10), 662 => to_unsigned(620, 10), 663 => to_unsigned(323, 10), 664 => to_unsigned(102, 10), 665 => to_unsigned(852, 10), 666 => to_unsigned(327, 10), 667 => to_unsigned(595, 10), 668 => to_unsigned(223, 10), 669 => to_unsigned(256, 10), 670 => to_unsigned(645, 10), 671 => to_unsigned(347, 10), 672 => to_unsigned(107, 10), 673 => to_unsigned(926, 10), 674 => to_unsigned(969, 10), 675 => to_unsigned(979, 10), 676 => to_unsigned(519, 10), 677 => to_unsigned(149, 10), 678 => to_unsigned(997, 10), 679 => to_unsigned(476, 10), 680 => to_unsigned(392, 10), 681 => to_unsigned(683, 10), 682 => to_unsigned(558, 10), 683 => to_unsigned(0, 10), 684 => to_unsigned(360, 10), 685 => to_unsigned(691, 10), 686 => to_unsigned(550, 10), 687 => to_unsigned(89, 10), 688 => to_unsigned(74, 10), 689 => to_unsigned(499, 10), 690 => to_unsigned(738, 10), 691 => to_unsigned(635, 10), 692 => to_unsigned(343, 10), 693 => to_unsigned(96, 10), 694 => to_unsigned(851, 10), 695 => to_unsigned(282, 10), 696 => to_unsigned(718, 10), 697 => to_unsigned(32, 10), 698 => to_unsigned(115, 10), 699 => to_unsigned(454, 10), 700 => to_unsigned(865, 10), 701 => to_unsigned(428, 10), 702 => to_unsigned(827, 10), 703 => to_unsigned(825, 10), 704 => to_unsigned(690, 10), 705 => to_unsigned(173, 10), 706 => to_unsigned(745, 10), 707 => to_unsigned(132, 10), 708 => to_unsigned(441, 10), 709 => to_unsigned(93, 10), 710 => to_unsigned(347, 10), 711 => to_unsigned(401, 10), 712 => to_unsigned(419, 10), 713 => to_unsigned(706, 10), 714 => to_unsigned(404, 10), 715 => to_unsigned(941, 10), 716 => to_unsigned(185, 10), 717 => to_unsigned(975, 10), 718 => to_unsigned(375, 10), 719 => to_unsigned(676, 10), 720 => to_unsigned(873, 10), 721 => to_unsigned(702, 10), 722 => to_unsigned(516, 10), 723 => to_unsigned(497, 10), 724 => to_unsigned(498, 10), 725 => to_unsigned(205, 10), 726 => to_unsigned(414, 10), 727 => to_unsigned(365, 10), 728 => to_unsigned(855, 10), 729 => to_unsigned(738, 10), 730 => to_unsigned(419, 10), 731 => to_unsigned(585, 10), 732 => to_unsigned(218, 10), 733 => to_unsigned(951, 10), 734 => to_unsigned(538, 10), 735 => to_unsigned(374, 10), 736 => to_unsigned(22, 10), 737 => to_unsigned(460, 10), 738 => to_unsigned(719, 10), 739 => to_unsigned(354, 10), 740 => to_unsigned(602, 10), 741 => to_unsigned(51, 10), 742 => to_unsigned(998, 10), 743 => to_unsigned(814, 10), 744 => to_unsigned(720, 10), 745 => to_unsigned(573, 10), 746 => to_unsigned(444, 10), 747 => to_unsigned(815, 10), 748 => to_unsigned(1018, 10), 749 => to_unsigned(104, 10), 750 => to_unsigned(640, 10), 751 => to_unsigned(394, 10), 752 => to_unsigned(971, 10), 753 => to_unsigned(909, 10), 754 => to_unsigned(327, 10), 755 => to_unsigned(606, 10), 756 => to_unsigned(518, 10), 757 => to_unsigned(685, 10), 758 => to_unsigned(245, 10), 759 => to_unsigned(414, 10), 760 => to_unsigned(527, 10), 761 => to_unsigned(169, 10), 762 => to_unsigned(166, 10), 763 => to_unsigned(309, 10), 764 => to_unsigned(939, 10), 765 => to_unsigned(594, 10), 766 => to_unsigned(391, 10), 767 => to_unsigned(220, 10), 768 => to_unsigned(833, 10), 769 => to_unsigned(681, 10), 770 => to_unsigned(834, 10), 771 => to_unsigned(114, 10), 772 => to_unsigned(860, 10), 773 => to_unsigned(334, 10), 774 => to_unsigned(741, 10), 775 => to_unsigned(219, 10), 776 => to_unsigned(246, 10), 777 => to_unsigned(100, 10), 778 => to_unsigned(415, 10), 779 => to_unsigned(221, 10), 780 => to_unsigned(178, 10), 781 => to_unsigned(508, 10), 782 => to_unsigned(174, 10), 783 => to_unsigned(605, 10), 784 => to_unsigned(626, 10), 785 => to_unsigned(673, 10), 786 => to_unsigned(780, 10), 787 => to_unsigned(736, 10), 788 => to_unsigned(745, 10), 789 => to_unsigned(848, 10), 790 => to_unsigned(66, 10), 791 => to_unsigned(456, 10), 792 => to_unsigned(1011, 10), 793 => to_unsigned(125, 10), 794 => to_unsigned(138, 10), 795 => to_unsigned(624, 10), 796 => to_unsigned(730, 10), 797 => to_unsigned(155, 10), 798 => to_unsigned(696, 10), 799 => to_unsigned(120, 10), 800 => to_unsigned(321, 10), 801 => to_unsigned(448, 10), 802 => to_unsigned(709, 10), 803 => to_unsigned(856, 10), 804 => to_unsigned(290, 10), 805 => to_unsigned(975, 10), 806 => to_unsigned(3, 10), 807 => to_unsigned(700, 10), 808 => to_unsigned(238, 10), 809 => to_unsigned(677, 10), 810 => to_unsigned(171, 10), 811 => to_unsigned(723, 10), 812 => to_unsigned(856, 10), 813 => to_unsigned(582, 10), 814 => to_unsigned(660, 10), 815 => to_unsigned(902, 10), 816 => to_unsigned(796, 10), 817 => to_unsigned(627, 10), 818 => to_unsigned(902, 10), 819 => to_unsigned(834, 10), 820 => to_unsigned(604, 10), 821 => to_unsigned(988, 10), 822 => to_unsigned(614, 10), 823 => to_unsigned(869, 10), 824 => to_unsigned(379, 10), 825 => to_unsigned(709, 10), 826 => to_unsigned(109, 10), 827 => to_unsigned(329, 10), 828 => to_unsigned(100, 10), 829 => to_unsigned(694, 10), 830 => to_unsigned(845, 10), 831 => to_unsigned(917, 10), 832 => to_unsigned(507, 10), 833 => to_unsigned(671, 10), 834 => to_unsigned(593, 10), 835 => to_unsigned(35, 10), 836 => to_unsigned(237, 10), 837 => to_unsigned(243, 10), 838 => to_unsigned(250, 10), 839 => to_unsigned(392, 10), 840 => to_unsigned(766, 10), 841 => to_unsigned(281, 10), 842 => to_unsigned(21, 10), 843 => to_unsigned(429, 10), 844 => to_unsigned(229, 10), 845 => to_unsigned(982, 10), 846 => to_unsigned(400, 10), 847 => to_unsigned(153, 10), 848 => to_unsigned(1006, 10), 849 => to_unsigned(119, 10), 850 => to_unsigned(677, 10), 851 => to_unsigned(895, 10), 852 => to_unsigned(385, 10), 853 => to_unsigned(389, 10), 854 => to_unsigned(710, 10), 855 => to_unsigned(396, 10), 856 => to_unsigned(346, 10), 857 => to_unsigned(586, 10), 858 => to_unsigned(1019, 10), 859 => to_unsigned(950, 10), 860 => to_unsigned(78, 10), 861 => to_unsigned(830, 10), 862 => to_unsigned(584, 10), 863 => to_unsigned(199, 10), 864 => to_unsigned(813, 10), 865 => to_unsigned(133, 10), 866 => to_unsigned(559, 10), 867 => to_unsigned(699, 10), 868 => to_unsigned(170, 10), 869 => to_unsigned(451, 10), 870 => to_unsigned(138, 10), 871 => to_unsigned(754, 10), 872 => to_unsigned(313, 10), 873 => to_unsigned(475, 10), 874 => to_unsigned(345, 10), 875 => to_unsigned(387, 10), 876 => to_unsigned(125, 10), 877 => to_unsigned(718, 10), 878 => to_unsigned(850, 10), 879 => to_unsigned(197, 10), 880 => to_unsigned(698, 10), 881 => to_unsigned(900, 10), 882 => to_unsigned(17, 10), 883 => to_unsigned(709, 10), 884 => to_unsigned(447, 10), 885 => to_unsigned(350, 10), 886 => to_unsigned(664, 10), 887 => to_unsigned(643, 10), 888 => to_unsigned(325, 10), 889 => to_unsigned(424, 10), 890 => to_unsigned(164, 10), 891 => to_unsigned(570, 10), 892 => to_unsigned(177, 10), 893 => to_unsigned(439, 10), 894 => to_unsigned(664, 10), 895 => to_unsigned(673, 10), 896 => to_unsigned(914, 10), 897 => to_unsigned(865, 10), 898 => to_unsigned(462, 10), 899 => to_unsigned(753, 10), 900 => to_unsigned(135, 10), 901 => to_unsigned(949, 10), 902 => to_unsigned(747, 10), 903 => to_unsigned(46, 10), 904 => to_unsigned(496, 10), 905 => to_unsigned(1012, 10), 906 => to_unsigned(639, 10), 907 => to_unsigned(929, 10), 908 => to_unsigned(337, 10), 909 => to_unsigned(157, 10), 910 => to_unsigned(524, 10), 911 => to_unsigned(630, 10), 912 => to_unsigned(814, 10), 913 => to_unsigned(886, 10), 914 => to_unsigned(288, 10), 915 => to_unsigned(802, 10), 916 => to_unsigned(115, 10), 917 => to_unsigned(599, 10), 918 => to_unsigned(636, 10), 919 => to_unsigned(409, 10), 920 => to_unsigned(174, 10), 921 => to_unsigned(498, 10), 922 => to_unsigned(875, 10), 923 => to_unsigned(564, 10), 924 => to_unsigned(1001, 10), 925 => to_unsigned(622, 10), 926 => to_unsigned(576, 10), 927 => to_unsigned(332, 10), 928 => to_unsigned(886, 10), 929 => to_unsigned(585, 10), 930 => to_unsigned(146, 10), 931 => to_unsigned(772, 10), 932 => to_unsigned(775, 10), 933 => to_unsigned(643, 10), 934 => to_unsigned(48, 10), 935 => to_unsigned(76, 10), 936 => to_unsigned(293, 10), 937 => to_unsigned(116, 10), 938 => to_unsigned(493, 10), 939 => to_unsigned(560, 10), 940 => to_unsigned(109, 10), 941 => to_unsigned(978, 10), 942 => to_unsigned(179, 10), 943 => to_unsigned(561, 10), 944 => to_unsigned(71, 10), 945 => to_unsigned(858, 10), 946 => to_unsigned(433, 10), 947 => to_unsigned(1006, 10), 948 => to_unsigned(285, 10), 949 => to_unsigned(515, 10), 950 => to_unsigned(74, 10), 951 => to_unsigned(596, 10), 952 => to_unsigned(490, 10), 953 => to_unsigned(321, 10), 954 => to_unsigned(887, 10), 955 => to_unsigned(532, 10), 956 => to_unsigned(208, 10), 957 => to_unsigned(42, 10), 958 => to_unsigned(498, 10), 959 => to_unsigned(28, 10), 960 => to_unsigned(410, 10), 961 => to_unsigned(855, 10), 962 => to_unsigned(180, 10), 963 => to_unsigned(304, 10), 964 => to_unsigned(962, 10), 965 => to_unsigned(614, 10), 966 => to_unsigned(777, 10), 967 => to_unsigned(258, 10), 968 => to_unsigned(372, 10), 969 => to_unsigned(876, 10), 970 => to_unsigned(745, 10), 971 => to_unsigned(857, 10), 972 => to_unsigned(380, 10), 973 => to_unsigned(885, 10), 974 => to_unsigned(612, 10), 975 => to_unsigned(90, 10), 976 => to_unsigned(68, 10), 977 => to_unsigned(617, 10), 978 => to_unsigned(522, 10), 979 => to_unsigned(12, 10), 980 => to_unsigned(616, 10), 981 => to_unsigned(225, 10), 982 => to_unsigned(421, 10), 983 => to_unsigned(167, 10), 984 => to_unsigned(928, 10), 985 => to_unsigned(378, 10), 986 => to_unsigned(289, 10), 987 => to_unsigned(922, 10), 988 => to_unsigned(99, 10), 989 => to_unsigned(217, 10), 990 => to_unsigned(306, 10), 991 => to_unsigned(344, 10), 992 => to_unsigned(210, 10), 993 => to_unsigned(788, 10), 994 => to_unsigned(734, 10), 995 => to_unsigned(668, 10), 996 => to_unsigned(584, 10), 997 => to_unsigned(274, 10), 998 => to_unsigned(409, 10), 999 => to_unsigned(920, 10), 1000 => to_unsigned(551, 10), 1001 => to_unsigned(234, 10), 1002 => to_unsigned(635, 10), 1003 => to_unsigned(284, 10), 1004 => to_unsigned(664, 10), 1005 => to_unsigned(658, 10), 1006 => to_unsigned(707, 10), 1007 => to_unsigned(172, 10), 1008 => to_unsigned(723, 10), 1009 => to_unsigned(301, 10), 1010 => to_unsigned(822, 10), 1011 => to_unsigned(0, 10), 1012 => to_unsigned(138, 10), 1013 => to_unsigned(707, 10), 1014 => to_unsigned(902, 10), 1015 => to_unsigned(731, 10), 1016 => to_unsigned(867, 10), 1017 => to_unsigned(441, 10), 1018 => to_unsigned(966, 10), 1019 => to_unsigned(915, 10), 1020 => to_unsigned(162, 10), 1021 => to_unsigned(50, 10), 1022 => to_unsigned(242, 10), 1023 => to_unsigned(870, 10), 1024 => to_unsigned(20, 10), 1025 => to_unsigned(683, 10), 1026 => to_unsigned(630, 10), 1027 => to_unsigned(128, 10), 1028 => to_unsigned(484, 10), 1029 => to_unsigned(365, 10), 1030 => to_unsigned(105, 10), 1031 => to_unsigned(706, 10), 1032 => to_unsigned(225, 10), 1033 => to_unsigned(652, 10), 1034 => to_unsigned(783, 10), 1035 => to_unsigned(118, 10), 1036 => to_unsigned(545, 10), 1037 => to_unsigned(151, 10), 1038 => to_unsigned(908, 10), 1039 => to_unsigned(901, 10), 1040 => to_unsigned(38, 10), 1041 => to_unsigned(769, 10), 1042 => to_unsigned(266, 10), 1043 => to_unsigned(6, 10), 1044 => to_unsigned(893, 10), 1045 => to_unsigned(262, 10), 1046 => to_unsigned(614, 10), 1047 => to_unsigned(934, 10), 1048 => to_unsigned(331, 10), 1049 => to_unsigned(370, 10), 1050 => to_unsigned(341, 10), 1051 => to_unsigned(382, 10), 1052 => to_unsigned(370, 10), 1053 => to_unsigned(690, 10), 1054 => to_unsigned(819, 10), 1055 => to_unsigned(258, 10), 1056 => to_unsigned(332, 10), 1057 => to_unsigned(669, 10), 1058 => to_unsigned(521, 10), 1059 => to_unsigned(627, 10), 1060 => to_unsigned(968, 10), 1061 => to_unsigned(389, 10), 1062 => to_unsigned(628, 10), 1063 => to_unsigned(181, 10), 1064 => to_unsigned(235, 10), 1065 => to_unsigned(193, 10), 1066 => to_unsigned(811, 10), 1067 => to_unsigned(591, 10), 1068 => to_unsigned(62, 10), 1069 => to_unsigned(332, 10), 1070 => to_unsigned(559, 10), 1071 => to_unsigned(588, 10), 1072 => to_unsigned(661, 10), 1073 => to_unsigned(120, 10), 1074 => to_unsigned(786, 10), 1075 => to_unsigned(345, 10), 1076 => to_unsigned(525, 10), 1077 => to_unsigned(222, 10), 1078 => to_unsigned(604, 10), 1079 => to_unsigned(236, 10), 1080 => to_unsigned(105, 10), 1081 => to_unsigned(213, 10), 1082 => to_unsigned(518, 10), 1083 => to_unsigned(612, 10), 1084 => to_unsigned(560, 10), 1085 => to_unsigned(552, 10), 1086 => to_unsigned(922, 10), 1087 => to_unsigned(158, 10), 1088 => to_unsigned(389, 10), 1089 => to_unsigned(143, 10), 1090 => to_unsigned(959, 10), 1091 => to_unsigned(485, 10), 1092 => to_unsigned(37, 10), 1093 => to_unsigned(571, 10), 1094 => to_unsigned(625, 10), 1095 => to_unsigned(95, 10), 1096 => to_unsigned(352, 10), 1097 => to_unsigned(496, 10), 1098 => to_unsigned(208, 10), 1099 => to_unsigned(288, 10), 1100 => to_unsigned(62, 10), 1101 => to_unsigned(394, 10), 1102 => to_unsigned(396, 10), 1103 => to_unsigned(605, 10), 1104 => to_unsigned(832, 10), 1105 => to_unsigned(413, 10), 1106 => to_unsigned(346, 10), 1107 => to_unsigned(999, 10), 1108 => to_unsigned(150, 10), 1109 => to_unsigned(403, 10), 1110 => to_unsigned(389, 10), 1111 => to_unsigned(804, 10), 1112 => to_unsigned(595, 10), 1113 => to_unsigned(127, 10), 1114 => to_unsigned(484, 10), 1115 => to_unsigned(773, 10), 1116 => to_unsigned(348, 10), 1117 => to_unsigned(460, 10), 1118 => to_unsigned(154, 10), 1119 => to_unsigned(753, 10), 1120 => to_unsigned(83, 10), 1121 => to_unsigned(908, 10), 1122 => to_unsigned(998, 10), 1123 => to_unsigned(135, 10), 1124 => to_unsigned(180, 10), 1125 => to_unsigned(592, 10), 1126 => to_unsigned(413, 10), 1127 => to_unsigned(0, 10), 1128 => to_unsigned(727, 10), 1129 => to_unsigned(719, 10), 1130 => to_unsigned(842, 10), 1131 => to_unsigned(764, 10), 1132 => to_unsigned(643, 10), 1133 => to_unsigned(573, 10), 1134 => to_unsigned(323, 10), 1135 => to_unsigned(144, 10), 1136 => to_unsigned(880, 10), 1137 => to_unsigned(457, 10), 1138 => to_unsigned(596, 10), 1139 => to_unsigned(116, 10), 1140 => to_unsigned(741, 10), 1141 => to_unsigned(767, 10), 1142 => to_unsigned(824, 10), 1143 => to_unsigned(318, 10), 1144 => to_unsigned(952, 10), 1145 => to_unsigned(560, 10), 1146 => to_unsigned(145, 10), 1147 => to_unsigned(885, 10), 1148 => to_unsigned(953, 10), 1149 => to_unsigned(521, 10), 1150 => to_unsigned(492, 10), 1151 => to_unsigned(190, 10), 1152 => to_unsigned(79, 10), 1153 => to_unsigned(742, 10), 1154 => to_unsigned(206, 10), 1155 => to_unsigned(417, 10), 1156 => to_unsigned(900, 10), 1157 => to_unsigned(912, 10), 1158 => to_unsigned(228, 10), 1159 => to_unsigned(839, 10), 1160 => to_unsigned(318, 10), 1161 => to_unsigned(791, 10), 1162 => to_unsigned(859, 10), 1163 => to_unsigned(366, 10), 1164 => to_unsigned(7, 10), 1165 => to_unsigned(509, 10), 1166 => to_unsigned(790, 10), 1167 => to_unsigned(866, 10), 1168 => to_unsigned(158, 10), 1169 => to_unsigned(758, 10), 1170 => to_unsigned(592, 10), 1171 => to_unsigned(155, 10), 1172 => to_unsigned(559, 10), 1173 => to_unsigned(495, 10), 1174 => to_unsigned(626, 10), 1175 => to_unsigned(523, 10), 1176 => to_unsigned(983, 10), 1177 => to_unsigned(846, 10), 1178 => to_unsigned(999, 10), 1179 => to_unsigned(798, 10), 1180 => to_unsigned(90, 10), 1181 => to_unsigned(290, 10), 1182 => to_unsigned(566, 10), 1183 => to_unsigned(849, 10), 1184 => to_unsigned(675, 10), 1185 => to_unsigned(71, 10), 1186 => to_unsigned(877, 10), 1187 => to_unsigned(827, 10), 1188 => to_unsigned(624, 10), 1189 => to_unsigned(421, 10), 1190 => to_unsigned(68, 10), 1191 => to_unsigned(437, 10), 1192 => to_unsigned(13, 10), 1193 => to_unsigned(101, 10), 1194 => to_unsigned(787, 10), 1195 => to_unsigned(875, 10), 1196 => to_unsigned(264, 10), 1197 => to_unsigned(864, 10), 1198 => to_unsigned(721, 10), 1199 => to_unsigned(197, 10), 1200 => to_unsigned(380, 10), 1201 => to_unsigned(100, 10), 1202 => to_unsigned(385, 10), 1203 => to_unsigned(765, 10), 1204 => to_unsigned(157, 10), 1205 => to_unsigned(901, 10), 1206 => to_unsigned(976, 10), 1207 => to_unsigned(230, 10), 1208 => to_unsigned(504, 10), 1209 => to_unsigned(936, 10), 1210 => to_unsigned(662, 10), 1211 => to_unsigned(30, 10), 1212 => to_unsigned(255, 10), 1213 => to_unsigned(531, 10), 1214 => to_unsigned(772, 10), 1215 => to_unsigned(660, 10), 1216 => to_unsigned(874, 10), 1217 => to_unsigned(586, 10), 1218 => to_unsigned(123, 10), 1219 => to_unsigned(451, 10), 1220 => to_unsigned(214, 10), 1221 => to_unsigned(316, 10), 1222 => to_unsigned(741, 10), 1223 => to_unsigned(250, 10), 1224 => to_unsigned(605, 10), 1225 => to_unsigned(681, 10), 1226 => to_unsigned(552, 10), 1227 => to_unsigned(188, 10), 1228 => to_unsigned(209, 10), 1229 => to_unsigned(691, 10), 1230 => to_unsigned(296, 10), 1231 => to_unsigned(59, 10), 1232 => to_unsigned(490, 10), 1233 => to_unsigned(478, 10), 1234 => to_unsigned(541, 10), 1235 => to_unsigned(225, 10), 1236 => to_unsigned(606, 10), 1237 => to_unsigned(238, 10), 1238 => to_unsigned(677, 10), 1239 => to_unsigned(382, 10), 1240 => to_unsigned(216, 10), 1241 => to_unsigned(272, 10), 1242 => to_unsigned(867, 10), 1243 => to_unsigned(167, 10), 1244 => to_unsigned(669, 10), 1245 => to_unsigned(508, 10), 1246 => to_unsigned(65, 10), 1247 => to_unsigned(791, 10), 1248 => to_unsigned(200, 10), 1249 => to_unsigned(384, 10), 1250 => to_unsigned(87, 10), 1251 => to_unsigned(805, 10), 1252 => to_unsigned(367, 10), 1253 => to_unsigned(447, 10), 1254 => to_unsigned(410, 10), 1255 => to_unsigned(729, 10), 1256 => to_unsigned(345, 10), 1257 => to_unsigned(134, 10), 1258 => to_unsigned(216, 10), 1259 => to_unsigned(503, 10), 1260 => to_unsigned(463, 10), 1261 => to_unsigned(101, 10), 1262 => to_unsigned(297, 10), 1263 => to_unsigned(913, 10), 1264 => to_unsigned(976, 10), 1265 => to_unsigned(880, 10), 1266 => to_unsigned(43, 10), 1267 => to_unsigned(110, 10), 1268 => to_unsigned(453, 10), 1269 => to_unsigned(374, 10), 1270 => to_unsigned(915, 10), 1271 => to_unsigned(751, 10), 1272 => to_unsigned(790, 10), 1273 => to_unsigned(365, 10), 1274 => to_unsigned(907, 10), 1275 => to_unsigned(523, 10), 1276 => to_unsigned(929, 10), 1277 => to_unsigned(903, 10), 1278 => to_unsigned(119, 10), 1279 => to_unsigned(282, 10), 1280 => to_unsigned(560, 10), 1281 => to_unsigned(199, 10), 1282 => to_unsigned(239, 10), 1283 => to_unsigned(694, 10), 1284 => to_unsigned(608, 10), 1285 => to_unsigned(356, 10), 1286 => to_unsigned(850, 10), 1287 => to_unsigned(599, 10), 1288 => to_unsigned(405, 10), 1289 => to_unsigned(510, 10), 1290 => to_unsigned(514, 10), 1291 => to_unsigned(264, 10), 1292 => to_unsigned(266, 10), 1293 => to_unsigned(261, 10), 1294 => to_unsigned(294, 10), 1295 => to_unsigned(934, 10), 1296 => to_unsigned(612, 10), 1297 => to_unsigned(449, 10), 1298 => to_unsigned(629, 10), 1299 => to_unsigned(571, 10), 1300 => to_unsigned(676, 10), 1301 => to_unsigned(901, 10), 1302 => to_unsigned(261, 10), 1303 => to_unsigned(38, 10), 1304 => to_unsigned(675, 10), 1305 => to_unsigned(88, 10), 1306 => to_unsigned(945, 10), 1307 => to_unsigned(719, 10), 1308 => to_unsigned(340, 10), 1309 => to_unsigned(370, 10), 1310 => to_unsigned(265, 10), 1311 => to_unsigned(1015, 10), 1312 => to_unsigned(132, 10), 1313 => to_unsigned(945, 10), 1314 => to_unsigned(24, 10), 1315 => to_unsigned(606, 10), 1316 => to_unsigned(386, 10), 1317 => to_unsigned(851, 10), 1318 => to_unsigned(899, 10), 1319 => to_unsigned(589, 10), 1320 => to_unsigned(267, 10), 1321 => to_unsigned(397, 10), 1322 => to_unsigned(484, 10), 1323 => to_unsigned(81, 10), 1324 => to_unsigned(154, 10), 1325 => to_unsigned(966, 10), 1326 => to_unsigned(687, 10), 1327 => to_unsigned(610, 10), 1328 => to_unsigned(533, 10), 1329 => to_unsigned(916, 10), 1330 => to_unsigned(682, 10), 1331 => to_unsigned(890, 10), 1332 => to_unsigned(441, 10), 1333 => to_unsigned(145, 10), 1334 => to_unsigned(613, 10), 1335 => to_unsigned(985, 10), 1336 => to_unsigned(244, 10), 1337 => to_unsigned(469, 10), 1338 => to_unsigned(183, 10), 1339 => to_unsigned(612, 10), 1340 => to_unsigned(196, 10), 1341 => to_unsigned(111, 10), 1342 => to_unsigned(226, 10), 1343 => to_unsigned(779, 10), 1344 => to_unsigned(994, 10), 1345 => to_unsigned(97, 10), 1346 => to_unsigned(238, 10), 1347 => to_unsigned(403, 10), 1348 => to_unsigned(880, 10), 1349 => to_unsigned(11, 10), 1350 => to_unsigned(993, 10), 1351 => to_unsigned(537, 10), 1352 => to_unsigned(97, 10), 1353 => to_unsigned(351, 10), 1354 => to_unsigned(301, 10), 1355 => to_unsigned(774, 10), 1356 => to_unsigned(601, 10), 1357 => to_unsigned(856, 10), 1358 => to_unsigned(493, 10), 1359 => to_unsigned(550, 10), 1360 => to_unsigned(51, 10), 1361 => to_unsigned(16, 10), 1362 => to_unsigned(919, 10), 1363 => to_unsigned(730, 10), 1364 => to_unsigned(771, 10), 1365 => to_unsigned(858, 10), 1366 => to_unsigned(430, 10), 1367 => to_unsigned(634, 10), 1368 => to_unsigned(413, 10), 1369 => to_unsigned(770, 10), 1370 => to_unsigned(645, 10), 1371 => to_unsigned(377, 10), 1372 => to_unsigned(967, 10), 1373 => to_unsigned(783, 10), 1374 => to_unsigned(846, 10), 1375 => to_unsigned(419, 10), 1376 => to_unsigned(180, 10), 1377 => to_unsigned(359, 10), 1378 => to_unsigned(886, 10), 1379 => to_unsigned(263, 10), 1380 => to_unsigned(691, 10), 1381 => to_unsigned(358, 10), 1382 => to_unsigned(761, 10), 1383 => to_unsigned(947, 10), 1384 => to_unsigned(925, 10), 1385 => to_unsigned(695, 10), 1386 => to_unsigned(625, 10), 1387 => to_unsigned(395, 10), 1388 => to_unsigned(451, 10), 1389 => to_unsigned(717, 10), 1390 => to_unsigned(890, 10), 1391 => to_unsigned(311, 10), 1392 => to_unsigned(600, 10), 1393 => to_unsigned(507, 10), 1394 => to_unsigned(252, 10), 1395 => to_unsigned(504, 10), 1396 => to_unsigned(836, 10), 1397 => to_unsigned(117, 10), 1398 => to_unsigned(371, 10), 1399 => to_unsigned(470, 10), 1400 => to_unsigned(185, 10), 1401 => to_unsigned(349, 10), 1402 => to_unsigned(614, 10), 1403 => to_unsigned(907, 10), 1404 => to_unsigned(718, 10), 1405 => to_unsigned(594, 10), 1406 => to_unsigned(985, 10), 1407 => to_unsigned(236, 10), 1408 => to_unsigned(3, 10), 1409 => to_unsigned(165, 10), 1410 => to_unsigned(391, 10), 1411 => to_unsigned(797, 10), 1412 => to_unsigned(78, 10), 1413 => to_unsigned(779, 10), 1414 => to_unsigned(969, 10), 1415 => to_unsigned(523, 10), 1416 => to_unsigned(784, 10), 1417 => to_unsigned(60, 10), 1418 => to_unsigned(635, 10), 1419 => to_unsigned(103, 10), 1420 => to_unsigned(703, 10), 1421 => to_unsigned(699, 10), 1422 => to_unsigned(129, 10), 1423 => to_unsigned(914, 10), 1424 => to_unsigned(693, 10), 1425 => to_unsigned(284, 10), 1426 => to_unsigned(448, 10), 1427 => to_unsigned(853, 10), 1428 => to_unsigned(728, 10), 1429 => to_unsigned(585, 10), 1430 => to_unsigned(904, 10), 1431 => to_unsigned(978, 10), 1432 => to_unsigned(395, 10), 1433 => to_unsigned(476, 10), 1434 => to_unsigned(373, 10), 1435 => to_unsigned(947, 10), 1436 => to_unsigned(849, 10), 1437 => to_unsigned(439, 10), 1438 => to_unsigned(15, 10), 1439 => to_unsigned(131, 10), 1440 => to_unsigned(106, 10), 1441 => to_unsigned(472, 10), 1442 => to_unsigned(213, 10), 1443 => to_unsigned(284, 10), 1444 => to_unsigned(826, 10), 1445 => to_unsigned(725, 10), 1446 => to_unsigned(590, 10), 1447 => to_unsigned(879, 10), 1448 => to_unsigned(833, 10), 1449 => to_unsigned(844, 10), 1450 => to_unsigned(267, 10), 1451 => to_unsigned(281, 10), 1452 => to_unsigned(359, 10), 1453 => to_unsigned(779, 10), 1454 => to_unsigned(858, 10), 1455 => to_unsigned(749, 10), 1456 => to_unsigned(418, 10), 1457 => to_unsigned(897, 10), 1458 => to_unsigned(1022, 10), 1459 => to_unsigned(656, 10), 1460 => to_unsigned(257, 10), 1461 => to_unsigned(528, 10), 1462 => to_unsigned(545, 10), 1463 => to_unsigned(33, 10), 1464 => to_unsigned(172, 10), 1465 => to_unsigned(486, 10), 1466 => to_unsigned(808, 10), 1467 => to_unsigned(328, 10), 1468 => to_unsigned(205, 10), 1469 => to_unsigned(106, 10), 1470 => to_unsigned(595, 10), 1471 => to_unsigned(754, 10), 1472 => to_unsigned(416, 10), 1473 => to_unsigned(919, 10), 1474 => to_unsigned(324, 10), 1475 => to_unsigned(415, 10), 1476 => to_unsigned(662, 10), 1477 => to_unsigned(64, 10), 1478 => to_unsigned(741, 10), 1479 => to_unsigned(287, 10), 1480 => to_unsigned(79, 10), 1481 => to_unsigned(83, 10), 1482 => to_unsigned(783, 10), 1483 => to_unsigned(819, 10), 1484 => to_unsigned(505, 10), 1485 => to_unsigned(396, 10), 1486 => to_unsigned(685, 10), 1487 => to_unsigned(10, 10), 1488 => to_unsigned(500, 10), 1489 => to_unsigned(617, 10), 1490 => to_unsigned(848, 10), 1491 => to_unsigned(70, 10), 1492 => to_unsigned(21, 10), 1493 => to_unsigned(734, 10), 1494 => to_unsigned(707, 10), 1495 => to_unsigned(336, 10), 1496 => to_unsigned(320, 10), 1497 => to_unsigned(129, 10), 1498 => to_unsigned(818, 10), 1499 => to_unsigned(864, 10), 1500 => to_unsigned(363, 10), 1501 => to_unsigned(1019, 10), 1502 => to_unsigned(466, 10), 1503 => to_unsigned(338, 10), 1504 => to_unsigned(697, 10), 1505 => to_unsigned(406, 10), 1506 => to_unsigned(783, 10), 1507 => to_unsigned(911, 10), 1508 => to_unsigned(540, 10), 1509 => to_unsigned(327, 10), 1510 => to_unsigned(283, 10), 1511 => to_unsigned(216, 10), 1512 => to_unsigned(313, 10), 1513 => to_unsigned(826, 10), 1514 => to_unsigned(216, 10), 1515 => to_unsigned(972, 10), 1516 => to_unsigned(269, 10), 1517 => to_unsigned(914, 10), 1518 => to_unsigned(78, 10), 1519 => to_unsigned(974, 10), 1520 => to_unsigned(788, 10), 1521 => to_unsigned(583, 10), 1522 => to_unsigned(695, 10), 1523 => to_unsigned(300, 10), 1524 => to_unsigned(235, 10), 1525 => to_unsigned(245, 10), 1526 => to_unsigned(91, 10), 1527 => to_unsigned(44, 10), 1528 => to_unsigned(783, 10), 1529 => to_unsigned(1021, 10), 1530 => to_unsigned(599, 10), 1531 => to_unsigned(971, 10), 1532 => to_unsigned(589, 10), 1533 => to_unsigned(510, 10), 1534 => to_unsigned(413, 10), 1535 => to_unsigned(607, 10), 1536 => to_unsigned(110, 10), 1537 => to_unsigned(722, 10), 1538 => to_unsigned(644, 10), 1539 => to_unsigned(540, 10), 1540 => to_unsigned(705, 10), 1541 => to_unsigned(49, 10), 1542 => to_unsigned(945, 10), 1543 => to_unsigned(343, 10), 1544 => to_unsigned(569, 10), 1545 => to_unsigned(720, 10), 1546 => to_unsigned(41, 10), 1547 => to_unsigned(474, 10), 1548 => to_unsigned(752, 10), 1549 => to_unsigned(194, 10), 1550 => to_unsigned(943, 10), 1551 => to_unsigned(273, 10), 1552 => to_unsigned(20, 10), 1553 => to_unsigned(678, 10), 1554 => to_unsigned(320, 10), 1555 => to_unsigned(646, 10), 1556 => to_unsigned(236, 10), 1557 => to_unsigned(662, 10), 1558 => to_unsigned(79, 10), 1559 => to_unsigned(74, 10), 1560 => to_unsigned(162, 10), 1561 => to_unsigned(680, 10), 1562 => to_unsigned(678, 10), 1563 => to_unsigned(1014, 10), 1564 => to_unsigned(661, 10), 1565 => to_unsigned(802, 10), 1566 => to_unsigned(373, 10), 1567 => to_unsigned(160, 10), 1568 => to_unsigned(426, 10), 1569 => to_unsigned(383, 10), 1570 => to_unsigned(300, 10), 1571 => to_unsigned(611, 10), 1572 => to_unsigned(809, 10), 1573 => to_unsigned(761, 10), 1574 => to_unsigned(871, 10), 1575 => to_unsigned(923, 10), 1576 => to_unsigned(763, 10), 1577 => to_unsigned(304, 10), 1578 => to_unsigned(383, 10), 1579 => to_unsigned(650, 10), 1580 => to_unsigned(324, 10), 1581 => to_unsigned(273, 10), 1582 => to_unsigned(771, 10), 1583 => to_unsigned(613, 10), 1584 => to_unsigned(606, 10), 1585 => to_unsigned(471, 10), 1586 => to_unsigned(285, 10), 1587 => to_unsigned(614, 10), 1588 => to_unsigned(635, 10), 1589 => to_unsigned(158, 10), 1590 => to_unsigned(203, 10), 1591 => to_unsigned(450, 10), 1592 => to_unsigned(477, 10), 1593 => to_unsigned(316, 10), 1594 => to_unsigned(647, 10), 1595 => to_unsigned(691, 10), 1596 => to_unsigned(244, 10), 1597 => to_unsigned(585, 10), 1598 => to_unsigned(471, 10), 1599 => to_unsigned(960, 10), 1600 => to_unsigned(1008, 10), 1601 => to_unsigned(401, 10), 1602 => to_unsigned(680, 10), 1603 => to_unsigned(243, 10), 1604 => to_unsigned(533, 10), 1605 => to_unsigned(606, 10), 1606 => to_unsigned(922, 10), 1607 => to_unsigned(143, 10), 1608 => to_unsigned(752, 10), 1609 => to_unsigned(785, 10), 1610 => to_unsigned(266, 10), 1611 => to_unsigned(657, 10), 1612 => to_unsigned(131, 10), 1613 => to_unsigned(999, 10), 1614 => to_unsigned(585, 10), 1615 => to_unsigned(797, 10), 1616 => to_unsigned(195, 10), 1617 => to_unsigned(455, 10), 1618 => to_unsigned(464, 10), 1619 => to_unsigned(226, 10), 1620 => to_unsigned(644, 10), 1621 => to_unsigned(445, 10), 1622 => to_unsigned(858, 10), 1623 => to_unsigned(100, 10), 1624 => to_unsigned(134, 10), 1625 => to_unsigned(32, 10), 1626 => to_unsigned(81, 10), 1627 => to_unsigned(631, 10), 1628 => to_unsigned(374, 10), 1629 => to_unsigned(757, 10), 1630 => to_unsigned(293, 10), 1631 => to_unsigned(631, 10), 1632 => to_unsigned(283, 10), 1633 => to_unsigned(51, 10), 1634 => to_unsigned(590, 10), 1635 => to_unsigned(955, 10), 1636 => to_unsigned(598, 10), 1637 => to_unsigned(607, 10), 1638 => to_unsigned(8, 10), 1639 => to_unsigned(312, 10), 1640 => to_unsigned(797, 10), 1641 => to_unsigned(668, 10), 1642 => to_unsigned(991, 10), 1643 => to_unsigned(418, 10), 1644 => to_unsigned(186, 10), 1645 => to_unsigned(895, 10), 1646 => to_unsigned(894, 10), 1647 => to_unsigned(977, 10), 1648 => to_unsigned(476, 10), 1649 => to_unsigned(111, 10), 1650 => to_unsigned(656, 10), 1651 => to_unsigned(968, 10), 1652 => to_unsigned(571, 10), 1653 => to_unsigned(247, 10), 1654 => to_unsigned(1004, 10), 1655 => to_unsigned(7, 10), 1656 => to_unsigned(908, 10), 1657 => to_unsigned(288, 10), 1658 => to_unsigned(724, 10), 1659 => to_unsigned(747, 10), 1660 => to_unsigned(75, 10), 1661 => to_unsigned(221, 10), 1662 => to_unsigned(40, 10), 1663 => to_unsigned(0, 10), 1664 => to_unsigned(212, 10), 1665 => to_unsigned(109, 10), 1666 => to_unsigned(604, 10), 1667 => to_unsigned(205, 10), 1668 => to_unsigned(165, 10), 1669 => to_unsigned(431, 10), 1670 => to_unsigned(573, 10), 1671 => to_unsigned(103, 10), 1672 => to_unsigned(946, 10), 1673 => to_unsigned(580, 10), 1674 => to_unsigned(494, 10), 1675 => to_unsigned(972, 10), 1676 => to_unsigned(697, 10), 1677 => to_unsigned(887, 10), 1678 => to_unsigned(997, 10), 1679 => to_unsigned(1008, 10), 1680 => to_unsigned(132, 10), 1681 => to_unsigned(617, 10), 1682 => to_unsigned(548, 10), 1683 => to_unsigned(336, 10), 1684 => to_unsigned(466, 10), 1685 => to_unsigned(165, 10), 1686 => to_unsigned(734, 10), 1687 => to_unsigned(373, 10), 1688 => to_unsigned(494, 10), 1689 => to_unsigned(291, 10), 1690 => to_unsigned(944, 10), 1691 => to_unsigned(640, 10), 1692 => to_unsigned(561, 10), 1693 => to_unsigned(185, 10), 1694 => to_unsigned(265, 10), 1695 => to_unsigned(50, 10), 1696 => to_unsigned(737, 10), 1697 => to_unsigned(176, 10), 1698 => to_unsigned(1009, 10), 1699 => to_unsigned(524, 10), 1700 => to_unsigned(710, 10), 1701 => to_unsigned(636, 10), 1702 => to_unsigned(499, 10), 1703 => to_unsigned(932, 10), 1704 => to_unsigned(99, 10), 1705 => to_unsigned(358, 10), 1706 => to_unsigned(36, 10), 1707 => to_unsigned(286, 10), 1708 => to_unsigned(626, 10), 1709 => to_unsigned(147, 10), 1710 => to_unsigned(422, 10), 1711 => to_unsigned(428, 10), 1712 => to_unsigned(35, 10), 1713 => to_unsigned(782, 10), 1714 => to_unsigned(29, 10), 1715 => to_unsigned(947, 10), 1716 => to_unsigned(60, 10), 1717 => to_unsigned(1016, 10), 1718 => to_unsigned(337, 10), 1719 => to_unsigned(835, 10), 1720 => to_unsigned(797, 10), 1721 => to_unsigned(155, 10), 1722 => to_unsigned(131, 10), 1723 => to_unsigned(33, 10), 1724 => to_unsigned(757, 10), 1725 => to_unsigned(435, 10), 1726 => to_unsigned(886, 10), 1727 => to_unsigned(411, 10), 1728 => to_unsigned(228, 10), 1729 => to_unsigned(56, 10), 1730 => to_unsigned(277, 10), 1731 => to_unsigned(679, 10), 1732 => to_unsigned(746, 10), 1733 => to_unsigned(330, 10), 1734 => to_unsigned(541, 10), 1735 => to_unsigned(241, 10), 1736 => to_unsigned(925, 10), 1737 => to_unsigned(957, 10), 1738 => to_unsigned(570, 10), 1739 => to_unsigned(792, 10), 1740 => to_unsigned(114, 10), 1741 => to_unsigned(272, 10), 1742 => to_unsigned(448, 10), 1743 => to_unsigned(868, 10), 1744 => to_unsigned(994, 10), 1745 => to_unsigned(635, 10), 1746 => to_unsigned(13, 10), 1747 => to_unsigned(769, 10), 1748 => to_unsigned(763, 10), 1749 => to_unsigned(258, 10), 1750 => to_unsigned(834, 10), 1751 => to_unsigned(147, 10), 1752 => to_unsigned(500, 10), 1753 => to_unsigned(762, 10), 1754 => to_unsigned(460, 10), 1755 => to_unsigned(670, 10), 1756 => to_unsigned(551, 10), 1757 => to_unsigned(469, 10), 1758 => to_unsigned(589, 10), 1759 => to_unsigned(945, 10), 1760 => to_unsigned(282, 10), 1761 => to_unsigned(371, 10), 1762 => to_unsigned(140, 10), 1763 => to_unsigned(241, 10), 1764 => to_unsigned(960, 10), 1765 => to_unsigned(257, 10), 1766 => to_unsigned(420, 10), 1767 => to_unsigned(778, 10), 1768 => to_unsigned(874, 10), 1769 => to_unsigned(288, 10), 1770 => to_unsigned(510, 10), 1771 => to_unsigned(284, 10), 1772 => to_unsigned(698, 10), 1773 => to_unsigned(706, 10), 1774 => to_unsigned(732, 10), 1775 => to_unsigned(65, 10), 1776 => to_unsigned(205, 10), 1777 => to_unsigned(339, 10), 1778 => to_unsigned(559, 10), 1779 => to_unsigned(593, 10), 1780 => to_unsigned(420, 10), 1781 => to_unsigned(199, 10), 1782 => to_unsigned(309, 10), 1783 => to_unsigned(710, 10), 1784 => to_unsigned(649, 10), 1785 => to_unsigned(527, 10), 1786 => to_unsigned(786, 10), 1787 => to_unsigned(157, 10), 1788 => to_unsigned(693, 10), 1789 => to_unsigned(956, 10), 1790 => to_unsigned(554, 10), 1791 => to_unsigned(466, 10), 1792 => to_unsigned(642, 10), 1793 => to_unsigned(797, 10), 1794 => to_unsigned(401, 10), 1795 => to_unsigned(35, 10), 1796 => to_unsigned(888, 10), 1797 => to_unsigned(275, 10), 1798 => to_unsigned(912, 10), 1799 => to_unsigned(535, 10), 1800 => to_unsigned(652, 10), 1801 => to_unsigned(355, 10), 1802 => to_unsigned(877, 10), 1803 => to_unsigned(696, 10), 1804 => to_unsigned(706, 10), 1805 => to_unsigned(788, 10), 1806 => to_unsigned(131, 10), 1807 => to_unsigned(81, 10), 1808 => to_unsigned(940, 10), 1809 => to_unsigned(38, 10), 1810 => to_unsigned(42, 10), 1811 => to_unsigned(970, 10), 1812 => to_unsigned(549, 10), 1813 => to_unsigned(362, 10), 1814 => to_unsigned(552, 10), 1815 => to_unsigned(879, 10), 1816 => to_unsigned(795, 10), 1817 => to_unsigned(644, 10), 1818 => to_unsigned(435, 10), 1819 => to_unsigned(406, 10), 1820 => to_unsigned(677, 10), 1821 => to_unsigned(803, 10), 1822 => to_unsigned(542, 10), 1823 => to_unsigned(775, 10), 1824 => to_unsigned(984, 10), 1825 => to_unsigned(600, 10), 1826 => to_unsigned(239, 10), 1827 => to_unsigned(911, 10), 1828 => to_unsigned(394, 10), 1829 => to_unsigned(147, 10), 1830 => to_unsigned(845, 10), 1831 => to_unsigned(999, 10), 1832 => to_unsigned(824, 10), 1833 => to_unsigned(997, 10), 1834 => to_unsigned(999, 10), 1835 => to_unsigned(914, 10), 1836 => to_unsigned(455, 10), 1837 => to_unsigned(60, 10), 1838 => to_unsigned(24, 10), 1839 => to_unsigned(160, 10), 1840 => to_unsigned(364, 10), 1841 => to_unsigned(295, 10), 1842 => to_unsigned(884, 10), 1843 => to_unsigned(104, 10), 1844 => to_unsigned(382, 10), 1845 => to_unsigned(367, 10), 1846 => to_unsigned(116, 10), 1847 => to_unsigned(996, 10), 1848 => to_unsigned(1002, 10), 1849 => to_unsigned(16, 10), 1850 => to_unsigned(948, 10), 1851 => to_unsigned(218, 10), 1852 => to_unsigned(1000, 10), 1853 => to_unsigned(208, 10), 1854 => to_unsigned(814, 10), 1855 => to_unsigned(224, 10), 1856 => to_unsigned(606, 10), 1857 => to_unsigned(852, 10), 1858 => to_unsigned(791, 10), 1859 => to_unsigned(655, 10), 1860 => to_unsigned(172, 10), 1861 => to_unsigned(595, 10), 1862 => to_unsigned(119, 10), 1863 => to_unsigned(567, 10), 1864 => to_unsigned(354, 10), 1865 => to_unsigned(411, 10), 1866 => to_unsigned(301, 10), 1867 => to_unsigned(994, 10), 1868 => to_unsigned(337, 10), 1869 => to_unsigned(727, 10), 1870 => to_unsigned(411, 10), 1871 => to_unsigned(589, 10), 1872 => to_unsigned(432, 10), 1873 => to_unsigned(983, 10), 1874 => to_unsigned(862, 10), 1875 => to_unsigned(389, 10), 1876 => to_unsigned(377, 10), 1877 => to_unsigned(231, 10), 1878 => to_unsigned(737, 10), 1879 => to_unsigned(881, 10), 1880 => to_unsigned(994, 10), 1881 => to_unsigned(796, 10), 1882 => to_unsigned(244, 10), 1883 => to_unsigned(65, 10), 1884 => to_unsigned(68, 10), 1885 => to_unsigned(725, 10), 1886 => to_unsigned(456, 10), 1887 => to_unsigned(764, 10), 1888 => to_unsigned(370, 10), 1889 => to_unsigned(929, 10), 1890 => to_unsigned(374, 10), 1891 => to_unsigned(483, 10), 1892 => to_unsigned(560, 10), 1893 => to_unsigned(99, 10), 1894 => to_unsigned(985, 10), 1895 => to_unsigned(581, 10), 1896 => to_unsigned(961, 10), 1897 => to_unsigned(611, 10), 1898 => to_unsigned(71, 10), 1899 => to_unsigned(513, 10), 1900 => to_unsigned(129, 10), 1901 => to_unsigned(199, 10), 1902 => to_unsigned(665, 10), 1903 => to_unsigned(100, 10), 1904 => to_unsigned(589, 10), 1905 => to_unsigned(620, 10), 1906 => to_unsigned(178, 10), 1907 => to_unsigned(411, 10), 1908 => to_unsigned(96, 10), 1909 => to_unsigned(555, 10), 1910 => to_unsigned(787, 10), 1911 => to_unsigned(354, 10), 1912 => to_unsigned(301, 10), 1913 => to_unsigned(100, 10), 1914 => to_unsigned(336, 10), 1915 => to_unsigned(112, 10), 1916 => to_unsigned(234, 10), 1917 => to_unsigned(889, 10), 1918 => to_unsigned(939, 10), 1919 => to_unsigned(451, 10), 1920 => to_unsigned(520, 10), 1921 => to_unsigned(211, 10), 1922 => to_unsigned(942, 10), 1923 => to_unsigned(576, 10), 1924 => to_unsigned(372, 10), 1925 => to_unsigned(916, 10), 1926 => to_unsigned(96, 10), 1927 => to_unsigned(482, 10), 1928 => to_unsigned(875, 10), 1929 => to_unsigned(389, 10), 1930 => to_unsigned(341, 10), 1931 => to_unsigned(280, 10), 1932 => to_unsigned(2, 10), 1933 => to_unsigned(509, 10), 1934 => to_unsigned(1021, 10), 1935 => to_unsigned(455, 10), 1936 => to_unsigned(108, 10), 1937 => to_unsigned(203, 10), 1938 => to_unsigned(243, 10), 1939 => to_unsigned(796, 10), 1940 => to_unsigned(374, 10), 1941 => to_unsigned(863, 10), 1942 => to_unsigned(65, 10), 1943 => to_unsigned(464, 10), 1944 => to_unsigned(370, 10), 1945 => to_unsigned(210, 10), 1946 => to_unsigned(398, 10), 1947 => to_unsigned(533, 10), 1948 => to_unsigned(111, 10), 1949 => to_unsigned(879, 10), 1950 => to_unsigned(197, 10), 1951 => to_unsigned(801, 10), 1952 => to_unsigned(618, 10), 1953 => to_unsigned(130, 10), 1954 => to_unsigned(539, 10), 1955 => to_unsigned(744, 10), 1956 => to_unsigned(375, 10), 1957 => to_unsigned(147, 10), 1958 => to_unsigned(911, 10), 1959 => to_unsigned(839, 10), 1960 => to_unsigned(1004, 10), 1961 => to_unsigned(797, 10), 1962 => to_unsigned(419, 10), 1963 => to_unsigned(737, 10), 1964 => to_unsigned(304, 10), 1965 => to_unsigned(945, 10), 1966 => to_unsigned(848, 10), 1967 => to_unsigned(184, 10), 1968 => to_unsigned(319, 10), 1969 => to_unsigned(472, 10), 1970 => to_unsigned(442, 10), 1971 => to_unsigned(901, 10), 1972 => to_unsigned(819, 10), 1973 => to_unsigned(250, 10), 1974 => to_unsigned(573, 10), 1975 => to_unsigned(106, 10), 1976 => to_unsigned(467, 10), 1977 => to_unsigned(273, 10), 1978 => to_unsigned(45, 10), 1979 => to_unsigned(992, 10), 1980 => to_unsigned(574, 10), 1981 => to_unsigned(22, 10), 1982 => to_unsigned(225, 10), 1983 => to_unsigned(614, 10), 1984 => to_unsigned(649, 10), 1985 => to_unsigned(773, 10), 1986 => to_unsigned(332, 10), 1987 => to_unsigned(573, 10), 1988 => to_unsigned(170, 10), 1989 => to_unsigned(759, 10), 1990 => to_unsigned(400, 10), 1991 => to_unsigned(315, 10), 1992 => to_unsigned(273, 10), 1993 => to_unsigned(196, 10), 1994 => to_unsigned(316, 10), 1995 => to_unsigned(665, 10), 1996 => to_unsigned(142, 10), 1997 => to_unsigned(877, 10), 1998 => to_unsigned(829, 10), 1999 => to_unsigned(181, 10), 2000 => to_unsigned(81, 10), 2001 => to_unsigned(541, 10), 2002 => to_unsigned(198, 10), 2003 => to_unsigned(28, 10), 2004 => to_unsigned(714, 10), 2005 => to_unsigned(645, 10), 2006 => to_unsigned(484, 10), 2007 => to_unsigned(484, 10), 2008 => to_unsigned(340, 10), 2009 => to_unsigned(951, 10), 2010 => to_unsigned(498, 10), 2011 => to_unsigned(178, 10), 2012 => to_unsigned(598, 10), 2013 => to_unsigned(181, 10), 2014 => to_unsigned(778, 10), 2015 => to_unsigned(555, 10), 2016 => to_unsigned(955, 10), 2017 => to_unsigned(414, 10), 2018 => to_unsigned(827, 10), 2019 => to_unsigned(142, 10), 2020 => to_unsigned(1011, 10), 2021 => to_unsigned(432, 10), 2022 => to_unsigned(632, 10), 2023 => to_unsigned(381, 10), 2024 => to_unsigned(56, 10), 2025 => to_unsigned(449, 10), 2026 => to_unsigned(872, 10), 2027 => to_unsigned(903, 10), 2028 => to_unsigned(965, 10), 2029 => to_unsigned(143, 10), 2030 => to_unsigned(631, 10), 2031 => to_unsigned(1001, 10), 2032 => to_unsigned(308, 10), 2033 => to_unsigned(288, 10), 2034 => to_unsigned(87, 10), 2035 => to_unsigned(974, 10), 2036 => to_unsigned(930, 10), 2037 => to_unsigned(541, 10), 2038 => to_unsigned(51, 10), 2039 => to_unsigned(473, 10), 2040 => to_unsigned(437, 10), 2041 => to_unsigned(772, 10), 2042 => to_unsigned(192, 10), 2043 => to_unsigned(891, 10), 2044 => to_unsigned(154, 10), 2045 => to_unsigned(468, 10), 2046 => to_unsigned(389, 10), 2047 => to_unsigned(378, 10)),
        1 => (0 => to_unsigned(570, 10), 1 => to_unsigned(241, 10), 2 => to_unsigned(332, 10), 3 => to_unsigned(597, 10), 4 => to_unsigned(972, 10), 5 => to_unsigned(80, 10), 6 => to_unsigned(599, 10), 7 => to_unsigned(714, 10), 8 => to_unsigned(848, 10), 9 => to_unsigned(85, 10), 10 => to_unsigned(89, 10), 11 => to_unsigned(19, 10), 12 => to_unsigned(482, 10), 13 => to_unsigned(919, 10), 14 => to_unsigned(144, 10), 15 => to_unsigned(364, 10), 16 => to_unsigned(672, 10), 17 => to_unsigned(577, 10), 18 => to_unsigned(346, 10), 19 => to_unsigned(525, 10), 20 => to_unsigned(286, 10), 21 => to_unsigned(163, 10), 22 => to_unsigned(1001, 10), 23 => to_unsigned(300, 10), 24 => to_unsigned(543, 10), 25 => to_unsigned(169, 10), 26 => to_unsigned(952, 10), 27 => to_unsigned(470, 10), 28 => to_unsigned(513, 10), 29 => to_unsigned(510, 10), 30 => to_unsigned(767, 10), 31 => to_unsigned(399, 10), 32 => to_unsigned(415, 10), 33 => to_unsigned(126, 10), 34 => to_unsigned(322, 10), 35 => to_unsigned(717, 10), 36 => to_unsigned(512, 10), 37 => to_unsigned(768, 10), 38 => to_unsigned(10, 10), 39 => to_unsigned(784, 10), 40 => to_unsigned(760, 10), 41 => to_unsigned(523, 10), 42 => to_unsigned(444, 10), 43 => to_unsigned(985, 10), 44 => to_unsigned(278, 10), 45 => to_unsigned(255, 10), 46 => to_unsigned(575, 10), 47 => to_unsigned(837, 10), 48 => to_unsigned(323, 10), 49 => to_unsigned(622, 10), 50 => to_unsigned(252, 10), 51 => to_unsigned(275, 10), 52 => to_unsigned(582, 10), 53 => to_unsigned(307, 10), 54 => to_unsigned(401, 10), 55 => to_unsigned(311, 10), 56 => to_unsigned(400, 10), 57 => to_unsigned(921, 10), 58 => to_unsigned(508, 10), 59 => to_unsigned(482, 10), 60 => to_unsigned(182, 10), 61 => to_unsigned(169, 10), 62 => to_unsigned(977, 10), 63 => to_unsigned(876, 10), 64 => to_unsigned(408, 10), 65 => to_unsigned(266, 10), 66 => to_unsigned(626, 10), 67 => to_unsigned(362, 10), 68 => to_unsigned(282, 10), 69 => to_unsigned(1019, 10), 70 => to_unsigned(55, 10), 71 => to_unsigned(247, 10), 72 => to_unsigned(612, 10), 73 => to_unsigned(380, 10), 74 => to_unsigned(222, 10), 75 => to_unsigned(880, 10), 76 => to_unsigned(722, 10), 77 => to_unsigned(640, 10), 78 => to_unsigned(3, 10), 79 => to_unsigned(190, 10), 80 => to_unsigned(98, 10), 81 => to_unsigned(796, 10), 82 => to_unsigned(511, 10), 83 => to_unsigned(767, 10), 84 => to_unsigned(906, 10), 85 => to_unsigned(593, 10), 86 => to_unsigned(584, 10), 87 => to_unsigned(957, 10), 88 => to_unsigned(917, 10), 89 => to_unsigned(431, 10), 90 => to_unsigned(603, 10), 91 => to_unsigned(78, 10), 92 => to_unsigned(408, 10), 93 => to_unsigned(850, 10), 94 => to_unsigned(802, 10), 95 => to_unsigned(1007, 10), 96 => to_unsigned(1018, 10), 97 => to_unsigned(887, 10), 98 => to_unsigned(979, 10), 99 => to_unsigned(367, 10), 100 => to_unsigned(604, 10), 101 => to_unsigned(971, 10), 102 => to_unsigned(722, 10), 103 => to_unsigned(832, 10), 104 => to_unsigned(422, 10), 105 => to_unsigned(234, 10), 106 => to_unsigned(1007, 10), 107 => to_unsigned(45, 10), 108 => to_unsigned(292, 10), 109 => to_unsigned(513, 10), 110 => to_unsigned(40, 10), 111 => to_unsigned(364, 10), 112 => to_unsigned(95, 10), 113 => to_unsigned(875, 10), 114 => to_unsigned(625, 10), 115 => to_unsigned(352, 10), 116 => to_unsigned(408, 10), 117 => to_unsigned(192, 10), 118 => to_unsigned(157, 10), 119 => to_unsigned(958, 10), 120 => to_unsigned(503, 10), 121 => to_unsigned(108, 10), 122 => to_unsigned(226, 10), 123 => to_unsigned(495, 10), 124 => to_unsigned(1010, 10), 125 => to_unsigned(1004, 10), 126 => to_unsigned(684, 10), 127 => to_unsigned(322, 10), 128 => to_unsigned(530, 10), 129 => to_unsigned(717, 10), 130 => to_unsigned(501, 10), 131 => to_unsigned(200, 10), 132 => to_unsigned(516, 10), 133 => to_unsigned(275, 10), 134 => to_unsigned(905, 10), 135 => to_unsigned(93, 10), 136 => to_unsigned(576, 10), 137 => to_unsigned(294, 10), 138 => to_unsigned(1009, 10), 139 => to_unsigned(534, 10), 140 => to_unsigned(921, 10), 141 => to_unsigned(539, 10), 142 => to_unsigned(657, 10), 143 => to_unsigned(701, 10), 144 => to_unsigned(698, 10), 145 => to_unsigned(246, 10), 146 => to_unsigned(345, 10), 147 => to_unsigned(118, 10), 148 => to_unsigned(118, 10), 149 => to_unsigned(107, 10), 150 => to_unsigned(971, 10), 151 => to_unsigned(454, 10), 152 => to_unsigned(324, 10), 153 => to_unsigned(670, 10), 154 => to_unsigned(648, 10), 155 => to_unsigned(828, 10), 156 => to_unsigned(655, 10), 157 => to_unsigned(531, 10), 158 => to_unsigned(144, 10), 159 => to_unsigned(480, 10), 160 => to_unsigned(860, 10), 161 => to_unsigned(266, 10), 162 => to_unsigned(698, 10), 163 => to_unsigned(157, 10), 164 => to_unsigned(717, 10), 165 => to_unsigned(679, 10), 166 => to_unsigned(995, 10), 167 => to_unsigned(369, 10), 168 => to_unsigned(115, 10), 169 => to_unsigned(299, 10), 170 => to_unsigned(442, 10), 171 => to_unsigned(1003, 10), 172 => to_unsigned(646, 10), 173 => to_unsigned(106, 10), 174 => to_unsigned(518, 10), 175 => to_unsigned(947, 10), 176 => to_unsigned(476, 10), 177 => to_unsigned(41, 10), 178 => to_unsigned(717, 10), 179 => to_unsigned(740, 10), 180 => to_unsigned(678, 10), 181 => to_unsigned(753, 10), 182 => to_unsigned(660, 10), 183 => to_unsigned(113, 10), 184 => to_unsigned(795, 10), 185 => to_unsigned(981, 10), 186 => to_unsigned(99, 10), 187 => to_unsigned(782, 10), 188 => to_unsigned(994, 10), 189 => to_unsigned(882, 10), 190 => to_unsigned(1010, 10), 191 => to_unsigned(1000, 10), 192 => to_unsigned(400, 10), 193 => to_unsigned(316, 10), 194 => to_unsigned(782, 10), 195 => to_unsigned(161, 10), 196 => to_unsigned(821, 10), 197 => to_unsigned(404, 10), 198 => to_unsigned(1006, 10), 199 => to_unsigned(336, 10), 200 => to_unsigned(54, 10), 201 => to_unsigned(94, 10), 202 => to_unsigned(810, 10), 203 => to_unsigned(142, 10), 204 => to_unsigned(882, 10), 205 => to_unsigned(917, 10), 206 => to_unsigned(775, 10), 207 => to_unsigned(185, 10), 208 => to_unsigned(818, 10), 209 => to_unsigned(185, 10), 210 => to_unsigned(673, 10), 211 => to_unsigned(777, 10), 212 => to_unsigned(257, 10), 213 => to_unsigned(968, 10), 214 => to_unsigned(389, 10), 215 => to_unsigned(110, 10), 216 => to_unsigned(556, 10), 217 => to_unsigned(667, 10), 218 => to_unsigned(150, 10), 219 => to_unsigned(771, 10), 220 => to_unsigned(827, 10), 221 => to_unsigned(760, 10), 222 => to_unsigned(979, 10), 223 => to_unsigned(175, 10), 224 => to_unsigned(824, 10), 225 => to_unsigned(459, 10), 226 => to_unsigned(51, 10), 227 => to_unsigned(235, 10), 228 => to_unsigned(68, 10), 229 => to_unsigned(306, 10), 230 => to_unsigned(648, 10), 231 => to_unsigned(100, 10), 232 => to_unsigned(163, 10), 233 => to_unsigned(565, 10), 234 => to_unsigned(463, 10), 235 => to_unsigned(17, 10), 236 => to_unsigned(886, 10), 237 => to_unsigned(469, 10), 238 => to_unsigned(571, 10), 239 => to_unsigned(322, 10), 240 => to_unsigned(987, 10), 241 => to_unsigned(583, 10), 242 => to_unsigned(410, 10), 243 => to_unsigned(0, 10), 244 => to_unsigned(608, 10), 245 => to_unsigned(264, 10), 246 => to_unsigned(319, 10), 247 => to_unsigned(954, 10), 248 => to_unsigned(71, 10), 249 => to_unsigned(442, 10), 250 => to_unsigned(92, 10), 251 => to_unsigned(879, 10), 252 => to_unsigned(283, 10), 253 => to_unsigned(333, 10), 254 => to_unsigned(404, 10), 255 => to_unsigned(703, 10), 256 => to_unsigned(357, 10), 257 => to_unsigned(145, 10), 258 => to_unsigned(880, 10), 259 => to_unsigned(88, 10), 260 => to_unsigned(980, 10), 261 => to_unsigned(68, 10), 262 => to_unsigned(524, 10), 263 => to_unsigned(11, 10), 264 => to_unsigned(522, 10), 265 => to_unsigned(568, 10), 266 => to_unsigned(845, 10), 267 => to_unsigned(58, 10), 268 => to_unsigned(523, 10), 269 => to_unsigned(672, 10), 270 => to_unsigned(220, 10), 271 => to_unsigned(316, 10), 272 => to_unsigned(971, 10), 273 => to_unsigned(423, 10), 274 => to_unsigned(965, 10), 275 => to_unsigned(241, 10), 276 => to_unsigned(627, 10), 277 => to_unsigned(417, 10), 278 => to_unsigned(740, 10), 279 => to_unsigned(189, 10), 280 => to_unsigned(353, 10), 281 => to_unsigned(161, 10), 282 => to_unsigned(518, 10), 283 => to_unsigned(158, 10), 284 => to_unsigned(486, 10), 285 => to_unsigned(859, 10), 286 => to_unsigned(398, 10), 287 => to_unsigned(97, 10), 288 => to_unsigned(986, 10), 289 => to_unsigned(995, 10), 290 => to_unsigned(855, 10), 291 => to_unsigned(468, 10), 292 => to_unsigned(707, 10), 293 => to_unsigned(982, 10), 294 => to_unsigned(325, 10), 295 => to_unsigned(781, 10), 296 => to_unsigned(159, 10), 297 => to_unsigned(755, 10), 298 => to_unsigned(719, 10), 299 => to_unsigned(325, 10), 300 => to_unsigned(820, 10), 301 => to_unsigned(81, 10), 302 => to_unsigned(870, 10), 303 => to_unsigned(479, 10), 304 => to_unsigned(115, 10), 305 => to_unsigned(344, 10), 306 => to_unsigned(854, 10), 307 => to_unsigned(953, 10), 308 => to_unsigned(785, 10), 309 => to_unsigned(635, 10), 310 => to_unsigned(190, 10), 311 => to_unsigned(836, 10), 312 => to_unsigned(107, 10), 313 => to_unsigned(977, 10), 314 => to_unsigned(173, 10), 315 => to_unsigned(182, 10), 316 => to_unsigned(703, 10), 317 => to_unsigned(489, 10), 318 => to_unsigned(838, 10), 319 => to_unsigned(1004, 10), 320 => to_unsigned(187, 10), 321 => to_unsigned(725, 10), 322 => to_unsigned(390, 10), 323 => to_unsigned(812, 10), 324 => to_unsigned(798, 10), 325 => to_unsigned(564, 10), 326 => to_unsigned(406, 10), 327 => to_unsigned(496, 10), 328 => to_unsigned(790, 10), 329 => to_unsigned(938, 10), 330 => to_unsigned(53, 10), 331 => to_unsigned(305, 10), 332 => to_unsigned(90, 10), 333 => to_unsigned(424, 10), 334 => to_unsigned(1015, 10), 335 => to_unsigned(845, 10), 336 => to_unsigned(776, 10), 337 => to_unsigned(303, 10), 338 => to_unsigned(509, 10), 339 => to_unsigned(908, 10), 340 => to_unsigned(984, 10), 341 => to_unsigned(495, 10), 342 => to_unsigned(1023, 10), 343 => to_unsigned(663, 10), 344 => to_unsigned(626, 10), 345 => to_unsigned(805, 10), 346 => to_unsigned(9, 10), 347 => to_unsigned(289, 10), 348 => to_unsigned(1016, 10), 349 => to_unsigned(604, 10), 350 => to_unsigned(481, 10), 351 => to_unsigned(650, 10), 352 => to_unsigned(898, 10), 353 => to_unsigned(219, 10), 354 => to_unsigned(142, 10), 355 => to_unsigned(858, 10), 356 => to_unsigned(771, 10), 357 => to_unsigned(531, 10), 358 => to_unsigned(447, 10), 359 => to_unsigned(716, 10), 360 => to_unsigned(567, 10), 361 => to_unsigned(218, 10), 362 => to_unsigned(842, 10), 363 => to_unsigned(818, 10), 364 => to_unsigned(920, 10), 365 => to_unsigned(996, 10), 366 => to_unsigned(696, 10), 367 => to_unsigned(883, 10), 368 => to_unsigned(938, 10), 369 => to_unsigned(1022, 10), 370 => to_unsigned(997, 10), 371 => to_unsigned(388, 10), 372 => to_unsigned(515, 10), 373 => to_unsigned(964, 10), 374 => to_unsigned(521, 10), 375 => to_unsigned(105, 10), 376 => to_unsigned(975, 10), 377 => to_unsigned(163, 10), 378 => to_unsigned(618, 10), 379 => to_unsigned(380, 10), 380 => to_unsigned(643, 10), 381 => to_unsigned(966, 10), 382 => to_unsigned(78, 10), 383 => to_unsigned(792, 10), 384 => to_unsigned(325, 10), 385 => to_unsigned(808, 10), 386 => to_unsigned(584, 10), 387 => to_unsigned(680, 10), 388 => to_unsigned(142, 10), 389 => to_unsigned(776, 10), 390 => to_unsigned(744, 10), 391 => to_unsigned(624, 10), 392 => to_unsigned(35, 10), 393 => to_unsigned(149, 10), 394 => to_unsigned(643, 10), 395 => to_unsigned(678, 10), 396 => to_unsigned(214, 10), 397 => to_unsigned(197, 10), 398 => to_unsigned(125, 10), 399 => to_unsigned(512, 10), 400 => to_unsigned(48, 10), 401 => to_unsigned(149, 10), 402 => to_unsigned(559, 10), 403 => to_unsigned(608, 10), 404 => to_unsigned(816, 10), 405 => to_unsigned(952, 10), 406 => to_unsigned(903, 10), 407 => to_unsigned(407, 10), 408 => to_unsigned(388, 10), 409 => to_unsigned(542, 10), 410 => to_unsigned(369, 10), 411 => to_unsigned(397, 10), 412 => to_unsigned(690, 10), 413 => to_unsigned(753, 10), 414 => to_unsigned(515, 10), 415 => to_unsigned(954, 10), 416 => to_unsigned(196, 10), 417 => to_unsigned(682, 10), 418 => to_unsigned(665, 10), 419 => to_unsigned(850, 10), 420 => to_unsigned(28, 10), 421 => to_unsigned(848, 10), 422 => to_unsigned(49, 10), 423 => to_unsigned(945, 10), 424 => to_unsigned(398, 10), 425 => to_unsigned(619, 10), 426 => to_unsigned(868, 10), 427 => to_unsigned(714, 10), 428 => to_unsigned(871, 10), 429 => to_unsigned(353, 10), 430 => to_unsigned(574, 10), 431 => to_unsigned(89, 10), 432 => to_unsigned(438, 10), 433 => to_unsigned(757, 10), 434 => to_unsigned(987, 10), 435 => to_unsigned(628, 10), 436 => to_unsigned(335, 10), 437 => to_unsigned(939, 10), 438 => to_unsigned(753, 10), 439 => to_unsigned(626, 10), 440 => to_unsigned(248, 10), 441 => to_unsigned(427, 10), 442 => to_unsigned(809, 10), 443 => to_unsigned(414, 10), 444 => to_unsigned(698, 10), 445 => to_unsigned(725, 10), 446 => to_unsigned(325, 10), 447 => to_unsigned(404, 10), 448 => to_unsigned(925, 10), 449 => to_unsigned(993, 10), 450 => to_unsigned(825, 10), 451 => to_unsigned(255, 10), 452 => to_unsigned(562, 10), 453 => to_unsigned(460, 10), 454 => to_unsigned(844, 10), 455 => to_unsigned(102, 10), 456 => to_unsigned(537, 10), 457 => to_unsigned(518, 10), 458 => to_unsigned(162, 10), 459 => to_unsigned(805, 10), 460 => to_unsigned(938, 10), 461 => to_unsigned(753, 10), 462 => to_unsigned(614, 10), 463 => to_unsigned(816, 10), 464 => to_unsigned(438, 10), 465 => to_unsigned(946, 10), 466 => to_unsigned(95, 10), 467 => to_unsigned(710, 10), 468 => to_unsigned(365, 10), 469 => to_unsigned(776, 10), 470 => to_unsigned(955, 10), 471 => to_unsigned(125, 10), 472 => to_unsigned(670, 10), 473 => to_unsigned(678, 10), 474 => to_unsigned(990, 10), 475 => to_unsigned(889, 10), 476 => to_unsigned(925, 10), 477 => to_unsigned(350, 10), 478 => to_unsigned(514, 10), 479 => to_unsigned(126, 10), 480 => to_unsigned(634, 10), 481 => to_unsigned(212, 10), 482 => to_unsigned(441, 10), 483 => to_unsigned(82, 10), 484 => to_unsigned(756, 10), 485 => to_unsigned(311, 10), 486 => to_unsigned(472, 10), 487 => to_unsigned(731, 10), 488 => to_unsigned(544, 10), 489 => to_unsigned(852, 10), 490 => to_unsigned(165, 10), 491 => to_unsigned(501, 10), 492 => to_unsigned(577, 10), 493 => to_unsigned(766, 10), 494 => to_unsigned(166, 10), 495 => to_unsigned(461, 10), 496 => to_unsigned(13, 10), 497 => to_unsigned(470, 10), 498 => to_unsigned(887, 10), 499 => to_unsigned(837, 10), 500 => to_unsigned(481, 10), 501 => to_unsigned(899, 10), 502 => to_unsigned(681, 10), 503 => to_unsigned(773, 10), 504 => to_unsigned(414, 10), 505 => to_unsigned(388, 10), 506 => to_unsigned(759, 10), 507 => to_unsigned(1004, 10), 508 => to_unsigned(1008, 10), 509 => to_unsigned(868, 10), 510 => to_unsigned(890, 10), 511 => to_unsigned(51, 10), 512 => to_unsigned(614, 10), 513 => to_unsigned(897, 10), 514 => to_unsigned(779, 10), 515 => to_unsigned(946, 10), 516 => to_unsigned(632, 10), 517 => to_unsigned(339, 10), 518 => to_unsigned(468, 10), 519 => to_unsigned(847, 10), 520 => to_unsigned(64, 10), 521 => to_unsigned(1023, 10), 522 => to_unsigned(237, 10), 523 => to_unsigned(437, 10), 524 => to_unsigned(294, 10), 525 => to_unsigned(344, 10), 526 => to_unsigned(921, 10), 527 => to_unsigned(106, 10), 528 => to_unsigned(115, 10), 529 => to_unsigned(974, 10), 530 => to_unsigned(656, 10), 531 => to_unsigned(866, 10), 532 => to_unsigned(925, 10), 533 => to_unsigned(693, 10), 534 => to_unsigned(1009, 10), 535 => to_unsigned(344, 10), 536 => to_unsigned(184, 10), 537 => to_unsigned(921, 10), 538 => to_unsigned(254, 10), 539 => to_unsigned(270, 10), 540 => to_unsigned(92, 10), 541 => to_unsigned(83, 10), 542 => to_unsigned(959, 10), 543 => to_unsigned(136, 10), 544 => to_unsigned(126, 10), 545 => to_unsigned(83, 10), 546 => to_unsigned(764, 10), 547 => to_unsigned(160, 10), 548 => to_unsigned(150, 10), 549 => to_unsigned(272, 10), 550 => to_unsigned(41, 10), 551 => to_unsigned(159, 10), 552 => to_unsigned(708, 10), 553 => to_unsigned(20, 10), 554 => to_unsigned(622, 10), 555 => to_unsigned(77, 10), 556 => to_unsigned(62, 10), 557 => to_unsigned(272, 10), 558 => to_unsigned(973, 10), 559 => to_unsigned(218, 10), 560 => to_unsigned(1016, 10), 561 => to_unsigned(544, 10), 562 => to_unsigned(198, 10), 563 => to_unsigned(381, 10), 564 => to_unsigned(229, 10), 565 => to_unsigned(728, 10), 566 => to_unsigned(777, 10), 567 => to_unsigned(1012, 10), 568 => to_unsigned(469, 10), 569 => to_unsigned(276, 10), 570 => to_unsigned(668, 10), 571 => to_unsigned(847, 10), 572 => to_unsigned(15, 10), 573 => to_unsigned(364, 10), 574 => to_unsigned(524, 10), 575 => to_unsigned(351, 10), 576 => to_unsigned(44, 10), 577 => to_unsigned(814, 10), 578 => to_unsigned(119, 10), 579 => to_unsigned(823, 10), 580 => to_unsigned(589, 10), 581 => to_unsigned(338, 10), 582 => to_unsigned(473, 10), 583 => to_unsigned(900, 10), 584 => to_unsigned(325, 10), 585 => to_unsigned(414, 10), 586 => to_unsigned(264, 10), 587 => to_unsigned(742, 10), 588 => to_unsigned(642, 10), 589 => to_unsigned(929, 10), 590 => to_unsigned(290, 10), 591 => to_unsigned(847, 10), 592 => to_unsigned(546, 10), 593 => to_unsigned(864, 10), 594 => to_unsigned(515, 10), 595 => to_unsigned(570, 10), 596 => to_unsigned(948, 10), 597 => to_unsigned(234, 10), 598 => to_unsigned(57, 10), 599 => to_unsigned(763, 10), 600 => to_unsigned(451, 10), 601 => to_unsigned(853, 10), 602 => to_unsigned(823, 10), 603 => to_unsigned(804, 10), 604 => to_unsigned(957, 10), 605 => to_unsigned(186, 10), 606 => to_unsigned(582, 10), 607 => to_unsigned(85, 10), 608 => to_unsigned(377, 10), 609 => to_unsigned(782, 10), 610 => to_unsigned(373, 10), 611 => to_unsigned(14, 10), 612 => to_unsigned(721, 10), 613 => to_unsigned(350, 10), 614 => to_unsigned(59, 10), 615 => to_unsigned(467, 10), 616 => to_unsigned(876, 10), 617 => to_unsigned(493, 10), 618 => to_unsigned(610, 10), 619 => to_unsigned(352, 10), 620 => to_unsigned(608, 10), 621 => to_unsigned(477, 10), 622 => to_unsigned(54, 10), 623 => to_unsigned(23, 10), 624 => to_unsigned(326, 10), 625 => to_unsigned(362, 10), 626 => to_unsigned(55, 10), 627 => to_unsigned(991, 10), 628 => to_unsigned(48, 10), 629 => to_unsigned(662, 10), 630 => to_unsigned(86, 10), 631 => to_unsigned(950, 10), 632 => to_unsigned(1003, 10), 633 => to_unsigned(352, 10), 634 => to_unsigned(897, 10), 635 => to_unsigned(509, 10), 636 => to_unsigned(852, 10), 637 => to_unsigned(660, 10), 638 => to_unsigned(653, 10), 639 => to_unsigned(318, 10), 640 => to_unsigned(966, 10), 641 => to_unsigned(357, 10), 642 => to_unsigned(574, 10), 643 => to_unsigned(176, 10), 644 => to_unsigned(802, 10), 645 => to_unsigned(229, 10), 646 => to_unsigned(486, 10), 647 => to_unsigned(980, 10), 648 => to_unsigned(1005, 10), 649 => to_unsigned(546, 10), 650 => to_unsigned(307, 10), 651 => to_unsigned(138, 10), 652 => to_unsigned(597, 10), 653 => to_unsigned(350, 10), 654 => to_unsigned(170, 10), 655 => to_unsigned(897, 10), 656 => to_unsigned(518, 10), 657 => to_unsigned(156, 10), 658 => to_unsigned(844, 10), 659 => to_unsigned(944, 10), 660 => to_unsigned(315, 10), 661 => to_unsigned(434, 10), 662 => to_unsigned(191, 10), 663 => to_unsigned(331, 10), 664 => to_unsigned(746, 10), 665 => to_unsigned(692, 10), 666 => to_unsigned(373, 10), 667 => to_unsigned(76, 10), 668 => to_unsigned(751, 10), 669 => to_unsigned(48, 10), 670 => to_unsigned(389, 10), 671 => to_unsigned(302, 10), 672 => to_unsigned(759, 10), 673 => to_unsigned(852, 10), 674 => to_unsigned(527, 10), 675 => to_unsigned(16, 10), 676 => to_unsigned(883, 10), 677 => to_unsigned(492, 10), 678 => to_unsigned(320, 10), 679 => to_unsigned(409, 10), 680 => to_unsigned(359, 10), 681 => to_unsigned(356, 10), 682 => to_unsigned(360, 10), 683 => to_unsigned(191, 10), 684 => to_unsigned(37, 10), 685 => to_unsigned(879, 10), 686 => to_unsigned(797, 10), 687 => to_unsigned(425, 10), 688 => to_unsigned(331, 10), 689 => to_unsigned(937, 10), 690 => to_unsigned(90, 10), 691 => to_unsigned(646, 10), 692 => to_unsigned(726, 10), 693 => to_unsigned(488, 10), 694 => to_unsigned(225, 10), 695 => to_unsigned(364, 10), 696 => to_unsigned(285, 10), 697 => to_unsigned(850, 10), 698 => to_unsigned(986, 10), 699 => to_unsigned(587, 10), 700 => to_unsigned(1013, 10), 701 => to_unsigned(433, 10), 702 => to_unsigned(981, 10), 703 => to_unsigned(136, 10), 704 => to_unsigned(362, 10), 705 => to_unsigned(429, 10), 706 => to_unsigned(1001, 10), 707 => to_unsigned(944, 10), 708 => to_unsigned(160, 10), 709 => to_unsigned(410, 10), 710 => to_unsigned(271, 10), 711 => to_unsigned(690, 10), 712 => to_unsigned(208, 10), 713 => to_unsigned(640, 10), 714 => to_unsigned(585, 10), 715 => to_unsigned(616, 10), 716 => to_unsigned(903, 10), 717 => to_unsigned(221, 10), 718 => to_unsigned(483, 10), 719 => to_unsigned(384, 10), 720 => to_unsigned(1008, 10), 721 => to_unsigned(928, 10), 722 => to_unsigned(992, 10), 723 => to_unsigned(398, 10), 724 => to_unsigned(562, 10), 725 => to_unsigned(71, 10), 726 => to_unsigned(610, 10), 727 => to_unsigned(280, 10), 728 => to_unsigned(802, 10), 729 => to_unsigned(656, 10), 730 => to_unsigned(778, 10), 731 => to_unsigned(566, 10), 732 => to_unsigned(754, 10), 733 => to_unsigned(9, 10), 734 => to_unsigned(395, 10), 735 => to_unsigned(1004, 10), 736 => to_unsigned(660, 10), 737 => to_unsigned(446, 10), 738 => to_unsigned(531, 10), 739 => to_unsigned(429, 10), 740 => to_unsigned(340, 10), 741 => to_unsigned(992, 10), 742 => to_unsigned(242, 10), 743 => to_unsigned(278, 10), 744 => to_unsigned(983, 10), 745 => to_unsigned(241, 10), 746 => to_unsigned(861, 10), 747 => to_unsigned(855, 10), 748 => to_unsigned(63, 10), 749 => to_unsigned(944, 10), 750 => to_unsigned(454, 10), 751 => to_unsigned(629, 10), 752 => to_unsigned(434, 10), 753 => to_unsigned(183, 10), 754 => to_unsigned(325, 10), 755 => to_unsigned(654, 10), 756 => to_unsigned(75, 10), 757 => to_unsigned(26, 10), 758 => to_unsigned(716, 10), 759 => to_unsigned(806, 10), 760 => to_unsigned(931, 10), 761 => to_unsigned(813, 10), 762 => to_unsigned(933, 10), 763 => to_unsigned(33, 10), 764 => to_unsigned(923, 10), 765 => to_unsigned(299, 10), 766 => to_unsigned(318, 10), 767 => to_unsigned(344, 10), 768 => to_unsigned(555, 10), 769 => to_unsigned(804, 10), 770 => to_unsigned(104, 10), 771 => to_unsigned(557, 10), 772 => to_unsigned(672, 10), 773 => to_unsigned(130, 10), 774 => to_unsigned(258, 10), 775 => to_unsigned(204, 10), 776 => to_unsigned(791, 10), 777 => to_unsigned(597, 10), 778 => to_unsigned(496, 10), 779 => to_unsigned(903, 10), 780 => to_unsigned(610, 10), 781 => to_unsigned(479, 10), 782 => to_unsigned(323, 10), 783 => to_unsigned(954, 10), 784 => to_unsigned(454, 10), 785 => to_unsigned(924, 10), 786 => to_unsigned(296, 10), 787 => to_unsigned(466, 10), 788 => to_unsigned(944, 10), 789 => to_unsigned(564, 10), 790 => to_unsigned(716, 10), 791 => to_unsigned(193, 10), 792 => to_unsigned(141, 10), 793 => to_unsigned(456, 10), 794 => to_unsigned(30, 10), 795 => to_unsigned(719, 10), 796 => to_unsigned(56, 10), 797 => to_unsigned(49, 10), 798 => to_unsigned(997, 10), 799 => to_unsigned(860, 10), 800 => to_unsigned(229, 10), 801 => to_unsigned(608, 10), 802 => to_unsigned(795, 10), 803 => to_unsigned(733, 10), 804 => to_unsigned(857, 10), 805 => to_unsigned(676, 10), 806 => to_unsigned(139, 10), 807 => to_unsigned(82, 10), 808 => to_unsigned(825, 10), 809 => to_unsigned(716, 10), 810 => to_unsigned(213, 10), 811 => to_unsigned(838, 10), 812 => to_unsigned(969, 10), 813 => to_unsigned(485, 10), 814 => to_unsigned(421, 10), 815 => to_unsigned(555, 10), 816 => to_unsigned(256, 10), 817 => to_unsigned(105, 10), 818 => to_unsigned(965, 10), 819 => to_unsigned(346, 10), 820 => to_unsigned(36, 10), 821 => to_unsigned(397, 10), 822 => to_unsigned(14, 10), 823 => to_unsigned(563, 10), 824 => to_unsigned(551, 10), 825 => to_unsigned(572, 10), 826 => to_unsigned(658, 10), 827 => to_unsigned(507, 10), 828 => to_unsigned(377, 10), 829 => to_unsigned(936, 10), 830 => to_unsigned(389, 10), 831 => to_unsigned(766, 10), 832 => to_unsigned(214, 10), 833 => to_unsigned(630, 10), 834 => to_unsigned(776, 10), 835 => to_unsigned(760, 10), 836 => to_unsigned(227, 10), 837 => to_unsigned(782, 10), 838 => to_unsigned(363, 10), 839 => to_unsigned(691, 10), 840 => to_unsigned(969, 10), 841 => to_unsigned(365, 10), 842 => to_unsigned(105, 10), 843 => to_unsigned(956, 10), 844 => to_unsigned(656, 10), 845 => to_unsigned(618, 10), 846 => to_unsigned(786, 10), 847 => to_unsigned(302, 10), 848 => to_unsigned(292, 10), 849 => to_unsigned(349, 10), 850 => to_unsigned(1010, 10), 851 => to_unsigned(449, 10), 852 => to_unsigned(999, 10), 853 => to_unsigned(469, 10), 854 => to_unsigned(762, 10), 855 => to_unsigned(817, 10), 856 => to_unsigned(291, 10), 857 => to_unsigned(343, 10), 858 => to_unsigned(708, 10), 859 => to_unsigned(509, 10), 860 => to_unsigned(833, 10), 861 => to_unsigned(758, 10), 862 => to_unsigned(533, 10), 863 => to_unsigned(947, 10), 864 => to_unsigned(287, 10), 865 => to_unsigned(355, 10), 866 => to_unsigned(134, 10), 867 => to_unsigned(514, 10), 868 => to_unsigned(655, 10), 869 => to_unsigned(699, 10), 870 => to_unsigned(1013, 10), 871 => to_unsigned(698, 10), 872 => to_unsigned(250, 10), 873 => to_unsigned(551, 10), 874 => to_unsigned(916, 10), 875 => to_unsigned(288, 10), 876 => to_unsigned(216, 10), 877 => to_unsigned(930, 10), 878 => to_unsigned(710, 10), 879 => to_unsigned(827, 10), 880 => to_unsigned(438, 10), 881 => to_unsigned(756, 10), 882 => to_unsigned(744, 10), 883 => to_unsigned(137, 10), 884 => to_unsigned(43, 10), 885 => to_unsigned(525, 10), 886 => to_unsigned(201, 10), 887 => to_unsigned(120, 10), 888 => to_unsigned(852, 10), 889 => to_unsigned(845, 10), 890 => to_unsigned(758, 10), 891 => to_unsigned(141, 10), 892 => to_unsigned(500, 10), 893 => to_unsigned(716, 10), 894 => to_unsigned(469, 10), 895 => to_unsigned(634, 10), 896 => to_unsigned(293, 10), 897 => to_unsigned(204, 10), 898 => to_unsigned(78, 10), 899 => to_unsigned(457, 10), 900 => to_unsigned(871, 10), 901 => to_unsigned(283, 10), 902 => to_unsigned(485, 10), 903 => to_unsigned(990, 10), 904 => to_unsigned(787, 10), 905 => to_unsigned(356, 10), 906 => to_unsigned(277, 10), 907 => to_unsigned(6, 10), 908 => to_unsigned(611, 10), 909 => to_unsigned(834, 10), 910 => to_unsigned(757, 10), 911 => to_unsigned(294, 10), 912 => to_unsigned(531, 10), 913 => to_unsigned(772, 10), 914 => to_unsigned(720, 10), 915 => to_unsigned(209, 10), 916 => to_unsigned(678, 10), 917 => to_unsigned(589, 10), 918 => to_unsigned(382, 10), 919 => to_unsigned(747, 10), 920 => to_unsigned(942, 10), 921 => to_unsigned(677, 10), 922 => to_unsigned(281, 10), 923 => to_unsigned(525, 10), 924 => to_unsigned(981, 10), 925 => to_unsigned(444, 10), 926 => to_unsigned(293, 10), 927 => to_unsigned(298, 10), 928 => to_unsigned(361, 10), 929 => to_unsigned(744, 10), 930 => to_unsigned(260, 10), 931 => to_unsigned(602, 10), 932 => to_unsigned(953, 10), 933 => to_unsigned(982, 10), 934 => to_unsigned(334, 10), 935 => to_unsigned(241, 10), 936 => to_unsigned(846, 10), 937 => to_unsigned(42, 10), 938 => to_unsigned(723, 10), 939 => to_unsigned(921, 10), 940 => to_unsigned(862, 10), 941 => to_unsigned(176, 10), 942 => to_unsigned(36, 10), 943 => to_unsigned(907, 10), 944 => to_unsigned(950, 10), 945 => to_unsigned(734, 10), 946 => to_unsigned(570, 10), 947 => to_unsigned(534, 10), 948 => to_unsigned(577, 10), 949 => to_unsigned(875, 10), 950 => to_unsigned(628, 10), 951 => to_unsigned(410, 10), 952 => to_unsigned(976, 10), 953 => to_unsigned(656, 10), 954 => to_unsigned(736, 10), 955 => to_unsigned(208, 10), 956 => to_unsigned(837, 10), 957 => to_unsigned(138, 10), 958 => to_unsigned(971, 10), 959 => to_unsigned(533, 10), 960 => to_unsigned(228, 10), 961 => to_unsigned(419, 10), 962 => to_unsigned(752, 10), 963 => to_unsigned(60, 10), 964 => to_unsigned(726, 10), 965 => to_unsigned(480, 10), 966 => to_unsigned(441, 10), 967 => to_unsigned(480, 10), 968 => to_unsigned(529, 10), 969 => to_unsigned(77, 10), 970 => to_unsigned(403, 10), 971 => to_unsigned(853, 10), 972 => to_unsigned(759, 10), 973 => to_unsigned(746, 10), 974 => to_unsigned(580, 10), 975 => to_unsigned(600, 10), 976 => to_unsigned(343, 10), 977 => to_unsigned(897, 10), 978 => to_unsigned(903, 10), 979 => to_unsigned(554, 10), 980 => to_unsigned(74, 10), 981 => to_unsigned(769, 10), 982 => to_unsigned(790, 10), 983 => to_unsigned(306, 10), 984 => to_unsigned(967, 10), 985 => to_unsigned(649, 10), 986 => to_unsigned(220, 10), 987 => to_unsigned(763, 10), 988 => to_unsigned(812, 10), 989 => to_unsigned(891, 10), 990 => to_unsigned(233, 10), 991 => to_unsigned(814, 10), 992 => to_unsigned(915, 10), 993 => to_unsigned(250, 10), 994 => to_unsigned(103, 10), 995 => to_unsigned(453, 10), 996 => to_unsigned(90, 10), 997 => to_unsigned(264, 10), 998 => to_unsigned(569, 10), 999 => to_unsigned(44, 10), 1000 => to_unsigned(85, 10), 1001 => to_unsigned(145, 10), 1002 => to_unsigned(645, 10), 1003 => to_unsigned(974, 10), 1004 => to_unsigned(352, 10), 1005 => to_unsigned(293, 10), 1006 => to_unsigned(667, 10), 1007 => to_unsigned(990, 10), 1008 => to_unsigned(61, 10), 1009 => to_unsigned(828, 10), 1010 => to_unsigned(188, 10), 1011 => to_unsigned(442, 10), 1012 => to_unsigned(184, 10), 1013 => to_unsigned(966, 10), 1014 => to_unsigned(204, 10), 1015 => to_unsigned(587, 10), 1016 => to_unsigned(155, 10), 1017 => to_unsigned(628, 10), 1018 => to_unsigned(209, 10), 1019 => to_unsigned(722, 10), 1020 => to_unsigned(207, 10), 1021 => to_unsigned(772, 10), 1022 => to_unsigned(528, 10), 1023 => to_unsigned(891, 10), 1024 => to_unsigned(359, 10), 1025 => to_unsigned(584, 10), 1026 => to_unsigned(139, 10), 1027 => to_unsigned(937, 10), 1028 => to_unsigned(42, 10), 1029 => to_unsigned(958, 10), 1030 => to_unsigned(780, 10), 1031 => to_unsigned(125, 10), 1032 => to_unsigned(804, 10), 1033 => to_unsigned(534, 10), 1034 => to_unsigned(890, 10), 1035 => to_unsigned(981, 10), 1036 => to_unsigned(124, 10), 1037 => to_unsigned(683, 10), 1038 => to_unsigned(636, 10), 1039 => to_unsigned(318, 10), 1040 => to_unsigned(639, 10), 1041 => to_unsigned(329, 10), 1042 => to_unsigned(376, 10), 1043 => to_unsigned(123, 10), 1044 => to_unsigned(844, 10), 1045 => to_unsigned(977, 10), 1046 => to_unsigned(215, 10), 1047 => to_unsigned(692, 10), 1048 => to_unsigned(55, 10), 1049 => to_unsigned(143, 10), 1050 => to_unsigned(387, 10), 1051 => to_unsigned(351, 10), 1052 => to_unsigned(58, 10), 1053 => to_unsigned(253, 10), 1054 => to_unsigned(303, 10), 1055 => to_unsigned(189, 10), 1056 => to_unsigned(139, 10), 1057 => to_unsigned(416, 10), 1058 => to_unsigned(618, 10), 1059 => to_unsigned(463, 10), 1060 => to_unsigned(921, 10), 1061 => to_unsigned(143, 10), 1062 => to_unsigned(833, 10), 1063 => to_unsigned(605, 10), 1064 => to_unsigned(528, 10), 1065 => to_unsigned(29, 10), 1066 => to_unsigned(312, 10), 1067 => to_unsigned(356, 10), 1068 => to_unsigned(605, 10), 1069 => to_unsigned(448, 10), 1070 => to_unsigned(573, 10), 1071 => to_unsigned(759, 10), 1072 => to_unsigned(295, 10), 1073 => to_unsigned(854, 10), 1074 => to_unsigned(258, 10), 1075 => to_unsigned(357, 10), 1076 => to_unsigned(688, 10), 1077 => to_unsigned(254, 10), 1078 => to_unsigned(787, 10), 1079 => to_unsigned(711, 10), 1080 => to_unsigned(910, 10), 1081 => to_unsigned(482, 10), 1082 => to_unsigned(926, 10), 1083 => to_unsigned(387, 10), 1084 => to_unsigned(586, 10), 1085 => to_unsigned(632, 10), 1086 => to_unsigned(236, 10), 1087 => to_unsigned(534, 10), 1088 => to_unsigned(815, 10), 1089 => to_unsigned(746, 10), 1090 => to_unsigned(822, 10), 1091 => to_unsigned(238, 10), 1092 => to_unsigned(983, 10), 1093 => to_unsigned(944, 10), 1094 => to_unsigned(127, 10), 1095 => to_unsigned(73, 10), 1096 => to_unsigned(545, 10), 1097 => to_unsigned(881, 10), 1098 => to_unsigned(218, 10), 1099 => to_unsigned(136, 10), 1100 => to_unsigned(157, 10), 1101 => to_unsigned(348, 10), 1102 => to_unsigned(993, 10), 1103 => to_unsigned(177, 10), 1104 => to_unsigned(360, 10), 1105 => to_unsigned(245, 10), 1106 => to_unsigned(182, 10), 1107 => to_unsigned(940, 10), 1108 => to_unsigned(892, 10), 1109 => to_unsigned(146, 10), 1110 => to_unsigned(462, 10), 1111 => to_unsigned(770, 10), 1112 => to_unsigned(1000, 10), 1113 => to_unsigned(650, 10), 1114 => to_unsigned(217, 10), 1115 => to_unsigned(326, 10), 1116 => to_unsigned(156, 10), 1117 => to_unsigned(53, 10), 1118 => to_unsigned(476, 10), 1119 => to_unsigned(400, 10), 1120 => to_unsigned(743, 10), 1121 => to_unsigned(85, 10), 1122 => to_unsigned(86, 10), 1123 => to_unsigned(61, 10), 1124 => to_unsigned(504, 10), 1125 => to_unsigned(722, 10), 1126 => to_unsigned(128, 10), 1127 => to_unsigned(968, 10), 1128 => to_unsigned(369, 10), 1129 => to_unsigned(322, 10), 1130 => to_unsigned(699, 10), 1131 => to_unsigned(1014, 10), 1132 => to_unsigned(9, 10), 1133 => to_unsigned(291, 10), 1134 => to_unsigned(845, 10), 1135 => to_unsigned(362, 10), 1136 => to_unsigned(442, 10), 1137 => to_unsigned(604, 10), 1138 => to_unsigned(428, 10), 1139 => to_unsigned(917, 10), 1140 => to_unsigned(0, 10), 1141 => to_unsigned(723, 10), 1142 => to_unsigned(456, 10), 1143 => to_unsigned(290, 10), 1144 => to_unsigned(954, 10), 1145 => to_unsigned(88, 10), 1146 => to_unsigned(819, 10), 1147 => to_unsigned(330, 10), 1148 => to_unsigned(500, 10), 1149 => to_unsigned(109, 10), 1150 => to_unsigned(908, 10), 1151 => to_unsigned(773, 10), 1152 => to_unsigned(996, 10), 1153 => to_unsigned(681, 10), 1154 => to_unsigned(884, 10), 1155 => to_unsigned(584, 10), 1156 => to_unsigned(194, 10), 1157 => to_unsigned(631, 10), 1158 => to_unsigned(242, 10), 1159 => to_unsigned(728, 10), 1160 => to_unsigned(745, 10), 1161 => to_unsigned(874, 10), 1162 => to_unsigned(666, 10), 1163 => to_unsigned(594, 10), 1164 => to_unsigned(37, 10), 1165 => to_unsigned(42, 10), 1166 => to_unsigned(766, 10), 1167 => to_unsigned(207, 10), 1168 => to_unsigned(145, 10), 1169 => to_unsigned(360, 10), 1170 => to_unsigned(143, 10), 1171 => to_unsigned(241, 10), 1172 => to_unsigned(1008, 10), 1173 => to_unsigned(128, 10), 1174 => to_unsigned(617, 10), 1175 => to_unsigned(992, 10), 1176 => to_unsigned(366, 10), 1177 => to_unsigned(887, 10), 1178 => to_unsigned(726, 10), 1179 => to_unsigned(675, 10), 1180 => to_unsigned(398, 10), 1181 => to_unsigned(125, 10), 1182 => to_unsigned(544, 10), 1183 => to_unsigned(288, 10), 1184 => to_unsigned(717, 10), 1185 => to_unsigned(314, 10), 1186 => to_unsigned(149, 10), 1187 => to_unsigned(150, 10), 1188 => to_unsigned(522, 10), 1189 => to_unsigned(533, 10), 1190 => to_unsigned(375, 10), 1191 => to_unsigned(979, 10), 1192 => to_unsigned(641, 10), 1193 => to_unsigned(937, 10), 1194 => to_unsigned(739, 10), 1195 => to_unsigned(976, 10), 1196 => to_unsigned(456, 10), 1197 => to_unsigned(3, 10), 1198 => to_unsigned(118, 10), 1199 => to_unsigned(725, 10), 1200 => to_unsigned(271, 10), 1201 => to_unsigned(24, 10), 1202 => to_unsigned(413, 10), 1203 => to_unsigned(983, 10), 1204 => to_unsigned(448, 10), 1205 => to_unsigned(748, 10), 1206 => to_unsigned(896, 10), 1207 => to_unsigned(951, 10), 1208 => to_unsigned(191, 10), 1209 => to_unsigned(33, 10), 1210 => to_unsigned(647, 10), 1211 => to_unsigned(155, 10), 1212 => to_unsigned(470, 10), 1213 => to_unsigned(90, 10), 1214 => to_unsigned(725, 10), 1215 => to_unsigned(484, 10), 1216 => to_unsigned(820, 10), 1217 => to_unsigned(565, 10), 1218 => to_unsigned(51, 10), 1219 => to_unsigned(89, 10), 1220 => to_unsigned(219, 10), 1221 => to_unsigned(777, 10), 1222 => to_unsigned(569, 10), 1223 => to_unsigned(182, 10), 1224 => to_unsigned(688, 10), 1225 => to_unsigned(413, 10), 1226 => to_unsigned(346, 10), 1227 => to_unsigned(393, 10), 1228 => to_unsigned(688, 10), 1229 => to_unsigned(925, 10), 1230 => to_unsigned(884, 10), 1231 => to_unsigned(683, 10), 1232 => to_unsigned(906, 10), 1233 => to_unsigned(1023, 10), 1234 => to_unsigned(422, 10), 1235 => to_unsigned(1001, 10), 1236 => to_unsigned(698, 10), 1237 => to_unsigned(406, 10), 1238 => to_unsigned(272, 10), 1239 => to_unsigned(980, 10), 1240 => to_unsigned(101, 10), 1241 => to_unsigned(684, 10), 1242 => to_unsigned(411, 10), 1243 => to_unsigned(266, 10), 1244 => to_unsigned(365, 10), 1245 => to_unsigned(167, 10), 1246 => to_unsigned(45, 10), 1247 => to_unsigned(428, 10), 1248 => to_unsigned(937, 10), 1249 => to_unsigned(605, 10), 1250 => to_unsigned(635, 10), 1251 => to_unsigned(1021, 10), 1252 => to_unsigned(133, 10), 1253 => to_unsigned(642, 10), 1254 => to_unsigned(304, 10), 1255 => to_unsigned(530, 10), 1256 => to_unsigned(996, 10), 1257 => to_unsigned(102, 10), 1258 => to_unsigned(607, 10), 1259 => to_unsigned(560, 10), 1260 => to_unsigned(823, 10), 1261 => to_unsigned(445, 10), 1262 => to_unsigned(136, 10), 1263 => to_unsigned(470, 10), 1264 => to_unsigned(934, 10), 1265 => to_unsigned(19, 10), 1266 => to_unsigned(762, 10), 1267 => to_unsigned(87, 10), 1268 => to_unsigned(645, 10), 1269 => to_unsigned(702, 10), 1270 => to_unsigned(284, 10), 1271 => to_unsigned(375, 10), 1272 => to_unsigned(801, 10), 1273 => to_unsigned(705, 10), 1274 => to_unsigned(58, 10), 1275 => to_unsigned(67, 10), 1276 => to_unsigned(945, 10), 1277 => to_unsigned(340, 10), 1278 => to_unsigned(718, 10), 1279 => to_unsigned(134, 10), 1280 => to_unsigned(939, 10), 1281 => to_unsigned(757, 10), 1282 => to_unsigned(875, 10), 1283 => to_unsigned(828, 10), 1284 => to_unsigned(667, 10), 1285 => to_unsigned(146, 10), 1286 => to_unsigned(605, 10), 1287 => to_unsigned(177, 10), 1288 => to_unsigned(897, 10), 1289 => to_unsigned(587, 10), 1290 => to_unsigned(477, 10), 1291 => to_unsigned(438, 10), 1292 => to_unsigned(173, 10), 1293 => to_unsigned(767, 10), 1294 => to_unsigned(375, 10), 1295 => to_unsigned(11, 10), 1296 => to_unsigned(924, 10), 1297 => to_unsigned(923, 10), 1298 => to_unsigned(951, 10), 1299 => to_unsigned(534, 10), 1300 => to_unsigned(154, 10), 1301 => to_unsigned(885, 10), 1302 => to_unsigned(675, 10), 1303 => to_unsigned(366, 10), 1304 => to_unsigned(86, 10), 1305 => to_unsigned(472, 10), 1306 => to_unsigned(88, 10), 1307 => to_unsigned(845, 10), 1308 => to_unsigned(486, 10), 1309 => to_unsigned(839, 10), 1310 => to_unsigned(77, 10), 1311 => to_unsigned(782, 10), 1312 => to_unsigned(795, 10), 1313 => to_unsigned(583, 10), 1314 => to_unsigned(341, 10), 1315 => to_unsigned(372, 10), 1316 => to_unsigned(455, 10), 1317 => to_unsigned(152, 10), 1318 => to_unsigned(303, 10), 1319 => to_unsigned(469, 10), 1320 => to_unsigned(122, 10), 1321 => to_unsigned(473, 10), 1322 => to_unsigned(125, 10), 1323 => to_unsigned(115, 10), 1324 => to_unsigned(805, 10), 1325 => to_unsigned(944, 10), 1326 => to_unsigned(969, 10), 1327 => to_unsigned(826, 10), 1328 => to_unsigned(564, 10), 1329 => to_unsigned(391, 10), 1330 => to_unsigned(513, 10), 1331 => to_unsigned(683, 10), 1332 => to_unsigned(889, 10), 1333 => to_unsigned(131, 10), 1334 => to_unsigned(871, 10), 1335 => to_unsigned(31, 10), 1336 => to_unsigned(20, 10), 1337 => to_unsigned(469, 10), 1338 => to_unsigned(528, 10), 1339 => to_unsigned(332, 10), 1340 => to_unsigned(315, 10), 1341 => to_unsigned(405, 10), 1342 => to_unsigned(70, 10), 1343 => to_unsigned(375, 10), 1344 => to_unsigned(521, 10), 1345 => to_unsigned(294, 10), 1346 => to_unsigned(330, 10), 1347 => to_unsigned(816, 10), 1348 => to_unsigned(798, 10), 1349 => to_unsigned(152, 10), 1350 => to_unsigned(169, 10), 1351 => to_unsigned(50, 10), 1352 => to_unsigned(72, 10), 1353 => to_unsigned(495, 10), 1354 => to_unsigned(807, 10), 1355 => to_unsigned(122, 10), 1356 => to_unsigned(193, 10), 1357 => to_unsigned(971, 10), 1358 => to_unsigned(627, 10), 1359 => to_unsigned(444, 10), 1360 => to_unsigned(731, 10), 1361 => to_unsigned(744, 10), 1362 => to_unsigned(37, 10), 1363 => to_unsigned(161, 10), 1364 => to_unsigned(32, 10), 1365 => to_unsigned(333, 10), 1366 => to_unsigned(644, 10), 1367 => to_unsigned(355, 10), 1368 => to_unsigned(817, 10), 1369 => to_unsigned(797, 10), 1370 => to_unsigned(129, 10), 1371 => to_unsigned(190, 10), 1372 => to_unsigned(565, 10), 1373 => to_unsigned(10, 10), 1374 => to_unsigned(198, 10), 1375 => to_unsigned(602, 10), 1376 => to_unsigned(41, 10), 1377 => to_unsigned(507, 10), 1378 => to_unsigned(798, 10), 1379 => to_unsigned(628, 10), 1380 => to_unsigned(716, 10), 1381 => to_unsigned(645, 10), 1382 => to_unsigned(535, 10), 1383 => to_unsigned(1014, 10), 1384 => to_unsigned(224, 10), 1385 => to_unsigned(447, 10), 1386 => to_unsigned(928, 10), 1387 => to_unsigned(581, 10), 1388 => to_unsigned(226, 10), 1389 => to_unsigned(152, 10), 1390 => to_unsigned(793, 10), 1391 => to_unsigned(391, 10), 1392 => to_unsigned(465, 10), 1393 => to_unsigned(984, 10), 1394 => to_unsigned(462, 10), 1395 => to_unsigned(401, 10), 1396 => to_unsigned(820, 10), 1397 => to_unsigned(645, 10), 1398 => to_unsigned(299, 10), 1399 => to_unsigned(929, 10), 1400 => to_unsigned(940, 10), 1401 => to_unsigned(421, 10), 1402 => to_unsigned(660, 10), 1403 => to_unsigned(741, 10), 1404 => to_unsigned(385, 10), 1405 => to_unsigned(524, 10), 1406 => to_unsigned(293, 10), 1407 => to_unsigned(875, 10), 1408 => to_unsigned(208, 10), 1409 => to_unsigned(174, 10), 1410 => to_unsigned(618, 10), 1411 => to_unsigned(228, 10), 1412 => to_unsigned(738, 10), 1413 => to_unsigned(64, 10), 1414 => to_unsigned(419, 10), 1415 => to_unsigned(178, 10), 1416 => to_unsigned(398, 10), 1417 => to_unsigned(601, 10), 1418 => to_unsigned(300, 10), 1419 => to_unsigned(46, 10), 1420 => to_unsigned(645, 10), 1421 => to_unsigned(829, 10), 1422 => to_unsigned(28, 10), 1423 => to_unsigned(716, 10), 1424 => to_unsigned(176, 10), 1425 => to_unsigned(742, 10), 1426 => to_unsigned(455, 10), 1427 => to_unsigned(723, 10), 1428 => to_unsigned(41, 10), 1429 => to_unsigned(469, 10), 1430 => to_unsigned(168, 10), 1431 => to_unsigned(255, 10), 1432 => to_unsigned(25, 10), 1433 => to_unsigned(832, 10), 1434 => to_unsigned(598, 10), 1435 => to_unsigned(299, 10), 1436 => to_unsigned(38, 10), 1437 => to_unsigned(245, 10), 1438 => to_unsigned(537, 10), 1439 => to_unsigned(383, 10), 1440 => to_unsigned(568, 10), 1441 => to_unsigned(428, 10), 1442 => to_unsigned(476, 10), 1443 => to_unsigned(769, 10), 1444 => to_unsigned(194, 10), 1445 => to_unsigned(438, 10), 1446 => to_unsigned(138, 10), 1447 => to_unsigned(749, 10), 1448 => to_unsigned(877, 10), 1449 => to_unsigned(182, 10), 1450 => to_unsigned(299, 10), 1451 => to_unsigned(269, 10), 1452 => to_unsigned(988, 10), 1453 => to_unsigned(749, 10), 1454 => to_unsigned(1, 10), 1455 => to_unsigned(767, 10), 1456 => to_unsigned(764, 10), 1457 => to_unsigned(501, 10), 1458 => to_unsigned(805, 10), 1459 => to_unsigned(740, 10), 1460 => to_unsigned(870, 10), 1461 => to_unsigned(434, 10), 1462 => to_unsigned(633, 10), 1463 => to_unsigned(482, 10), 1464 => to_unsigned(872, 10), 1465 => to_unsigned(296, 10), 1466 => to_unsigned(482, 10), 1467 => to_unsigned(239, 10), 1468 => to_unsigned(154, 10), 1469 => to_unsigned(235, 10), 1470 => to_unsigned(729, 10), 1471 => to_unsigned(601, 10), 1472 => to_unsigned(569, 10), 1473 => to_unsigned(190, 10), 1474 => to_unsigned(646, 10), 1475 => to_unsigned(911, 10), 1476 => to_unsigned(570, 10), 1477 => to_unsigned(1015, 10), 1478 => to_unsigned(46, 10), 1479 => to_unsigned(350, 10), 1480 => to_unsigned(903, 10), 1481 => to_unsigned(205, 10), 1482 => to_unsigned(727, 10), 1483 => to_unsigned(236, 10), 1484 => to_unsigned(27, 10), 1485 => to_unsigned(842, 10), 1486 => to_unsigned(954, 10), 1487 => to_unsigned(420, 10), 1488 => to_unsigned(665, 10), 1489 => to_unsigned(1014, 10), 1490 => to_unsigned(334, 10), 1491 => to_unsigned(737, 10), 1492 => to_unsigned(888, 10), 1493 => to_unsigned(425, 10), 1494 => to_unsigned(183, 10), 1495 => to_unsigned(999, 10), 1496 => to_unsigned(870, 10), 1497 => to_unsigned(799, 10), 1498 => to_unsigned(633, 10), 1499 => to_unsigned(339, 10), 1500 => to_unsigned(522, 10), 1501 => to_unsigned(183, 10), 1502 => to_unsigned(409, 10), 1503 => to_unsigned(934, 10), 1504 => to_unsigned(712, 10), 1505 => to_unsigned(166, 10), 1506 => to_unsigned(136, 10), 1507 => to_unsigned(348, 10), 1508 => to_unsigned(564, 10), 1509 => to_unsigned(67, 10), 1510 => to_unsigned(328, 10), 1511 => to_unsigned(348, 10), 1512 => to_unsigned(938, 10), 1513 => to_unsigned(617, 10), 1514 => to_unsigned(190, 10), 1515 => to_unsigned(910, 10), 1516 => to_unsigned(273, 10), 1517 => to_unsigned(1001, 10), 1518 => to_unsigned(145, 10), 1519 => to_unsigned(650, 10), 1520 => to_unsigned(708, 10), 1521 => to_unsigned(895, 10), 1522 => to_unsigned(733, 10), 1523 => to_unsigned(544, 10), 1524 => to_unsigned(870, 10), 1525 => to_unsigned(696, 10), 1526 => to_unsigned(483, 10), 1527 => to_unsigned(77, 10), 1528 => to_unsigned(669, 10), 1529 => to_unsigned(958, 10), 1530 => to_unsigned(211, 10), 1531 => to_unsigned(236, 10), 1532 => to_unsigned(11, 10), 1533 => to_unsigned(677, 10), 1534 => to_unsigned(355, 10), 1535 => to_unsigned(771, 10), 1536 => to_unsigned(578, 10), 1537 => to_unsigned(122, 10), 1538 => to_unsigned(273, 10), 1539 => to_unsigned(193, 10), 1540 => to_unsigned(310, 10), 1541 => to_unsigned(257, 10), 1542 => to_unsigned(947, 10), 1543 => to_unsigned(779, 10), 1544 => to_unsigned(925, 10), 1545 => to_unsigned(130, 10), 1546 => to_unsigned(280, 10), 1547 => to_unsigned(695, 10), 1548 => to_unsigned(412, 10), 1549 => to_unsigned(285, 10), 1550 => to_unsigned(684, 10), 1551 => to_unsigned(196, 10), 1552 => to_unsigned(317, 10), 1553 => to_unsigned(798, 10), 1554 => to_unsigned(792, 10), 1555 => to_unsigned(935, 10), 1556 => to_unsigned(349, 10), 1557 => to_unsigned(532, 10), 1558 => to_unsigned(628, 10), 1559 => to_unsigned(854, 10), 1560 => to_unsigned(919, 10), 1561 => to_unsigned(267, 10), 1562 => to_unsigned(948, 10), 1563 => to_unsigned(605, 10), 1564 => to_unsigned(396, 10), 1565 => to_unsigned(750, 10), 1566 => to_unsigned(161, 10), 1567 => to_unsigned(3, 10), 1568 => to_unsigned(327, 10), 1569 => to_unsigned(826, 10), 1570 => to_unsigned(171, 10), 1571 => to_unsigned(357, 10), 1572 => to_unsigned(908, 10), 1573 => to_unsigned(24, 10), 1574 => to_unsigned(241, 10), 1575 => to_unsigned(986, 10), 1576 => to_unsigned(757, 10), 1577 => to_unsigned(15, 10), 1578 => to_unsigned(117, 10), 1579 => to_unsigned(662, 10), 1580 => to_unsigned(483, 10), 1581 => to_unsigned(353, 10), 1582 => to_unsigned(890, 10), 1583 => to_unsigned(592, 10), 1584 => to_unsigned(620, 10), 1585 => to_unsigned(125, 10), 1586 => to_unsigned(247, 10), 1587 => to_unsigned(192, 10), 1588 => to_unsigned(886, 10), 1589 => to_unsigned(196, 10), 1590 => to_unsigned(518, 10), 1591 => to_unsigned(434, 10), 1592 => to_unsigned(377, 10), 1593 => to_unsigned(926, 10), 1594 => to_unsigned(762, 10), 1595 => to_unsigned(723, 10), 1596 => to_unsigned(528, 10), 1597 => to_unsigned(81, 10), 1598 => to_unsigned(413, 10), 1599 => to_unsigned(365, 10), 1600 => to_unsigned(588, 10), 1601 => to_unsigned(330, 10), 1602 => to_unsigned(401, 10), 1603 => to_unsigned(501, 10), 1604 => to_unsigned(694, 10), 1605 => to_unsigned(994, 10), 1606 => to_unsigned(808, 10), 1607 => to_unsigned(472, 10), 1608 => to_unsigned(27, 10), 1609 => to_unsigned(546, 10), 1610 => to_unsigned(442, 10), 1611 => to_unsigned(782, 10), 1612 => to_unsigned(776, 10), 1613 => to_unsigned(52, 10), 1614 => to_unsigned(812, 10), 1615 => to_unsigned(914, 10), 1616 => to_unsigned(475, 10), 1617 => to_unsigned(218, 10), 1618 => to_unsigned(1010, 10), 1619 => to_unsigned(727, 10), 1620 => to_unsigned(455, 10), 1621 => to_unsigned(970, 10), 1622 => to_unsigned(962, 10), 1623 => to_unsigned(21, 10), 1624 => to_unsigned(716, 10), 1625 => to_unsigned(102, 10), 1626 => to_unsigned(395, 10), 1627 => to_unsigned(662, 10), 1628 => to_unsigned(956, 10), 1629 => to_unsigned(679, 10), 1630 => to_unsigned(461, 10), 1631 => to_unsigned(1017, 10), 1632 => to_unsigned(289, 10), 1633 => to_unsigned(1001, 10), 1634 => to_unsigned(984, 10), 1635 => to_unsigned(757, 10), 1636 => to_unsigned(251, 10), 1637 => to_unsigned(695, 10), 1638 => to_unsigned(471, 10), 1639 => to_unsigned(599, 10), 1640 => to_unsigned(220, 10), 1641 => to_unsigned(270, 10), 1642 => to_unsigned(989, 10), 1643 => to_unsigned(189, 10), 1644 => to_unsigned(427, 10), 1645 => to_unsigned(167, 10), 1646 => to_unsigned(961, 10), 1647 => to_unsigned(348, 10), 1648 => to_unsigned(757, 10), 1649 => to_unsigned(432, 10), 1650 => to_unsigned(574, 10), 1651 => to_unsigned(626, 10), 1652 => to_unsigned(758, 10), 1653 => to_unsigned(478, 10), 1654 => to_unsigned(143, 10), 1655 => to_unsigned(351, 10), 1656 => to_unsigned(412, 10), 1657 => to_unsigned(264, 10), 1658 => to_unsigned(356, 10), 1659 => to_unsigned(876, 10), 1660 => to_unsigned(467, 10), 1661 => to_unsigned(527, 10), 1662 => to_unsigned(1014, 10), 1663 => to_unsigned(82, 10), 1664 => to_unsigned(873, 10), 1665 => to_unsigned(699, 10), 1666 => to_unsigned(320, 10), 1667 => to_unsigned(576, 10), 1668 => to_unsigned(567, 10), 1669 => to_unsigned(689, 10), 1670 => to_unsigned(317, 10), 1671 => to_unsigned(961, 10), 1672 => to_unsigned(330, 10), 1673 => to_unsigned(222, 10), 1674 => to_unsigned(906, 10), 1675 => to_unsigned(419, 10), 1676 => to_unsigned(514, 10), 1677 => to_unsigned(769, 10), 1678 => to_unsigned(457, 10), 1679 => to_unsigned(1014, 10), 1680 => to_unsigned(938, 10), 1681 => to_unsigned(112, 10), 1682 => to_unsigned(884, 10), 1683 => to_unsigned(451, 10), 1684 => to_unsigned(494, 10), 1685 => to_unsigned(363, 10), 1686 => to_unsigned(36, 10), 1687 => to_unsigned(525, 10), 1688 => to_unsigned(163, 10), 1689 => to_unsigned(245, 10), 1690 => to_unsigned(783, 10), 1691 => to_unsigned(690, 10), 1692 => to_unsigned(878, 10), 1693 => to_unsigned(969, 10), 1694 => to_unsigned(871, 10), 1695 => to_unsigned(978, 10), 1696 => to_unsigned(962, 10), 1697 => to_unsigned(941, 10), 1698 => to_unsigned(553, 10), 1699 => to_unsigned(4, 10), 1700 => to_unsigned(764, 10), 1701 => to_unsigned(108, 10), 1702 => to_unsigned(462, 10), 1703 => to_unsigned(911, 10), 1704 => to_unsigned(108, 10), 1705 => to_unsigned(980, 10), 1706 => to_unsigned(473, 10), 1707 => to_unsigned(554, 10), 1708 => to_unsigned(978, 10), 1709 => to_unsigned(854, 10), 1710 => to_unsigned(916, 10), 1711 => to_unsigned(382, 10), 1712 => to_unsigned(491, 10), 1713 => to_unsigned(885, 10), 1714 => to_unsigned(302, 10), 1715 => to_unsigned(828, 10), 1716 => to_unsigned(1002, 10), 1717 => to_unsigned(818, 10), 1718 => to_unsigned(450, 10), 1719 => to_unsigned(967, 10), 1720 => to_unsigned(944, 10), 1721 => to_unsigned(914, 10), 1722 => to_unsigned(77, 10), 1723 => to_unsigned(321, 10), 1724 => to_unsigned(307, 10), 1725 => to_unsigned(372, 10), 1726 => to_unsigned(608, 10), 1727 => to_unsigned(451, 10), 1728 => to_unsigned(1014, 10), 1729 => to_unsigned(868, 10), 1730 => to_unsigned(176, 10), 1731 => to_unsigned(1008, 10), 1732 => to_unsigned(541, 10), 1733 => to_unsigned(67, 10), 1734 => to_unsigned(581, 10), 1735 => to_unsigned(667, 10), 1736 => to_unsigned(394, 10), 1737 => to_unsigned(52, 10), 1738 => to_unsigned(238, 10), 1739 => to_unsigned(774, 10), 1740 => to_unsigned(780, 10), 1741 => to_unsigned(321, 10), 1742 => to_unsigned(323, 10), 1743 => to_unsigned(703, 10), 1744 => to_unsigned(8, 10), 1745 => to_unsigned(356, 10), 1746 => to_unsigned(395, 10), 1747 => to_unsigned(465, 10), 1748 => to_unsigned(872, 10), 1749 => to_unsigned(34, 10), 1750 => to_unsigned(259, 10), 1751 => to_unsigned(673, 10), 1752 => to_unsigned(659, 10), 1753 => to_unsigned(643, 10), 1754 => to_unsigned(237, 10), 1755 => to_unsigned(93, 10), 1756 => to_unsigned(282, 10), 1757 => to_unsigned(731, 10), 1758 => to_unsigned(359, 10), 1759 => to_unsigned(499, 10), 1760 => to_unsigned(1008, 10), 1761 => to_unsigned(837, 10), 1762 => to_unsigned(662, 10), 1763 => to_unsigned(468, 10), 1764 => to_unsigned(589, 10), 1765 => to_unsigned(218, 10), 1766 => to_unsigned(927, 10), 1767 => to_unsigned(242, 10), 1768 => to_unsigned(38, 10), 1769 => to_unsigned(901, 10), 1770 => to_unsigned(689, 10), 1771 => to_unsigned(742, 10), 1772 => to_unsigned(137, 10), 1773 => to_unsigned(231, 10), 1774 => to_unsigned(349, 10), 1775 => to_unsigned(876, 10), 1776 => to_unsigned(184, 10), 1777 => to_unsigned(189, 10), 1778 => to_unsigned(648, 10), 1779 => to_unsigned(992, 10), 1780 => to_unsigned(946, 10), 1781 => to_unsigned(656, 10), 1782 => to_unsigned(405, 10), 1783 => to_unsigned(735, 10), 1784 => to_unsigned(107, 10), 1785 => to_unsigned(504, 10), 1786 => to_unsigned(248, 10), 1787 => to_unsigned(938, 10), 1788 => to_unsigned(965, 10), 1789 => to_unsigned(242, 10), 1790 => to_unsigned(131, 10), 1791 => to_unsigned(59, 10), 1792 => to_unsigned(88, 10), 1793 => to_unsigned(478, 10), 1794 => to_unsigned(11, 10), 1795 => to_unsigned(633, 10), 1796 => to_unsigned(748, 10), 1797 => to_unsigned(425, 10), 1798 => to_unsigned(547, 10), 1799 => to_unsigned(247, 10), 1800 => to_unsigned(538, 10), 1801 => to_unsigned(627, 10), 1802 => to_unsigned(176, 10), 1803 => to_unsigned(130, 10), 1804 => to_unsigned(390, 10), 1805 => to_unsigned(305, 10), 1806 => to_unsigned(623, 10), 1807 => to_unsigned(11, 10), 1808 => to_unsigned(42, 10), 1809 => to_unsigned(533, 10), 1810 => to_unsigned(126, 10), 1811 => to_unsigned(789, 10), 1812 => to_unsigned(80, 10), 1813 => to_unsigned(776, 10), 1814 => to_unsigned(215, 10), 1815 => to_unsigned(871, 10), 1816 => to_unsigned(1008, 10), 1817 => to_unsigned(725, 10), 1818 => to_unsigned(960, 10), 1819 => to_unsigned(485, 10), 1820 => to_unsigned(239, 10), 1821 => to_unsigned(523, 10), 1822 => to_unsigned(675, 10), 1823 => to_unsigned(738, 10), 1824 => to_unsigned(346, 10), 1825 => to_unsigned(544, 10), 1826 => to_unsigned(97, 10), 1827 => to_unsigned(107, 10), 1828 => to_unsigned(764, 10), 1829 => to_unsigned(470, 10), 1830 => to_unsigned(403, 10), 1831 => to_unsigned(1000, 10), 1832 => to_unsigned(486, 10), 1833 => to_unsigned(565, 10), 1834 => to_unsigned(744, 10), 1835 => to_unsigned(56, 10), 1836 => to_unsigned(509, 10), 1837 => to_unsigned(701, 10), 1838 => to_unsigned(441, 10), 1839 => to_unsigned(66, 10), 1840 => to_unsigned(604, 10), 1841 => to_unsigned(544, 10), 1842 => to_unsigned(263, 10), 1843 => to_unsigned(253, 10), 1844 => to_unsigned(655, 10), 1845 => to_unsigned(619, 10), 1846 => to_unsigned(863, 10), 1847 => to_unsigned(1009, 10), 1848 => to_unsigned(734, 10), 1849 => to_unsigned(428, 10), 1850 => to_unsigned(469, 10), 1851 => to_unsigned(209, 10), 1852 => to_unsigned(205, 10), 1853 => to_unsigned(482, 10), 1854 => to_unsigned(816, 10), 1855 => to_unsigned(987, 10), 1856 => to_unsigned(200, 10), 1857 => to_unsigned(676, 10), 1858 => to_unsigned(468, 10), 1859 => to_unsigned(612, 10), 1860 => to_unsigned(666, 10), 1861 => to_unsigned(823, 10), 1862 => to_unsigned(37, 10), 1863 => to_unsigned(178, 10), 1864 => to_unsigned(620, 10), 1865 => to_unsigned(674, 10), 1866 => to_unsigned(10, 10), 1867 => to_unsigned(735, 10), 1868 => to_unsigned(340, 10), 1869 => to_unsigned(783, 10), 1870 => to_unsigned(875, 10), 1871 => to_unsigned(45, 10), 1872 => to_unsigned(889, 10), 1873 => to_unsigned(682, 10), 1874 => to_unsigned(279, 10), 1875 => to_unsigned(444, 10), 1876 => to_unsigned(942, 10), 1877 => to_unsigned(779, 10), 1878 => to_unsigned(917, 10), 1879 => to_unsigned(522, 10), 1880 => to_unsigned(961, 10), 1881 => to_unsigned(579, 10), 1882 => to_unsigned(307, 10), 1883 => to_unsigned(889, 10), 1884 => to_unsigned(292, 10), 1885 => to_unsigned(305, 10), 1886 => to_unsigned(481, 10), 1887 => to_unsigned(892, 10), 1888 => to_unsigned(452, 10), 1889 => to_unsigned(712, 10), 1890 => to_unsigned(323, 10), 1891 => to_unsigned(867, 10), 1892 => to_unsigned(847, 10), 1893 => to_unsigned(820, 10), 1894 => to_unsigned(350, 10), 1895 => to_unsigned(168, 10), 1896 => to_unsigned(895, 10), 1897 => to_unsigned(849, 10), 1898 => to_unsigned(801, 10), 1899 => to_unsigned(530, 10), 1900 => to_unsigned(639, 10), 1901 => to_unsigned(323, 10), 1902 => to_unsigned(1017, 10), 1903 => to_unsigned(533, 10), 1904 => to_unsigned(696, 10), 1905 => to_unsigned(563, 10), 1906 => to_unsigned(500, 10), 1907 => to_unsigned(237, 10), 1908 => to_unsigned(726, 10), 1909 => to_unsigned(464, 10), 1910 => to_unsigned(718, 10), 1911 => to_unsigned(729, 10), 1912 => to_unsigned(525, 10), 1913 => to_unsigned(387, 10), 1914 => to_unsigned(985, 10), 1915 => to_unsigned(762, 10), 1916 => to_unsigned(465, 10), 1917 => to_unsigned(460, 10), 1918 => to_unsigned(29, 10), 1919 => to_unsigned(686, 10), 1920 => to_unsigned(173, 10), 1921 => to_unsigned(217, 10), 1922 => to_unsigned(325, 10), 1923 => to_unsigned(492, 10), 1924 => to_unsigned(520, 10), 1925 => to_unsigned(942, 10), 1926 => to_unsigned(249, 10), 1927 => to_unsigned(176, 10), 1928 => to_unsigned(250, 10), 1929 => to_unsigned(704, 10), 1930 => to_unsigned(66, 10), 1931 => to_unsigned(61, 10), 1932 => to_unsigned(393, 10), 1933 => to_unsigned(11, 10), 1934 => to_unsigned(319, 10), 1935 => to_unsigned(799, 10), 1936 => to_unsigned(918, 10), 1937 => to_unsigned(801, 10), 1938 => to_unsigned(447, 10), 1939 => to_unsigned(943, 10), 1940 => to_unsigned(84, 10), 1941 => to_unsigned(713, 10), 1942 => to_unsigned(854, 10), 1943 => to_unsigned(347, 10), 1944 => to_unsigned(329, 10), 1945 => to_unsigned(147, 10), 1946 => to_unsigned(983, 10), 1947 => to_unsigned(185, 10), 1948 => to_unsigned(951, 10), 1949 => to_unsigned(820, 10), 1950 => to_unsigned(252, 10), 1951 => to_unsigned(984, 10), 1952 => to_unsigned(372, 10), 1953 => to_unsigned(217, 10), 1954 => to_unsigned(626, 10), 1955 => to_unsigned(198, 10), 1956 => to_unsigned(819, 10), 1957 => to_unsigned(291, 10), 1958 => to_unsigned(592, 10), 1959 => to_unsigned(479, 10), 1960 => to_unsigned(545, 10), 1961 => to_unsigned(389, 10), 1962 => to_unsigned(700, 10), 1963 => to_unsigned(909, 10), 1964 => to_unsigned(267, 10), 1965 => to_unsigned(363, 10), 1966 => to_unsigned(683, 10), 1967 => to_unsigned(965, 10), 1968 => to_unsigned(458, 10), 1969 => to_unsigned(210, 10), 1970 => to_unsigned(834, 10), 1971 => to_unsigned(702, 10), 1972 => to_unsigned(119, 10), 1973 => to_unsigned(656, 10), 1974 => to_unsigned(256, 10), 1975 => to_unsigned(269, 10), 1976 => to_unsigned(48, 10), 1977 => to_unsigned(918, 10), 1978 => to_unsigned(929, 10), 1979 => to_unsigned(768, 10), 1980 => to_unsigned(490, 10), 1981 => to_unsigned(585, 10), 1982 => to_unsigned(665, 10), 1983 => to_unsigned(104, 10), 1984 => to_unsigned(313, 10), 1985 => to_unsigned(570, 10), 1986 => to_unsigned(450, 10), 1987 => to_unsigned(526, 10), 1988 => to_unsigned(374, 10), 1989 => to_unsigned(826, 10), 1990 => to_unsigned(924, 10), 1991 => to_unsigned(725, 10), 1992 => to_unsigned(962, 10), 1993 => to_unsigned(406, 10), 1994 => to_unsigned(509, 10), 1995 => to_unsigned(200, 10), 1996 => to_unsigned(239, 10), 1997 => to_unsigned(464, 10), 1998 => to_unsigned(291, 10), 1999 => to_unsigned(493, 10), 2000 => to_unsigned(923, 10), 2001 => to_unsigned(866, 10), 2002 => to_unsigned(313, 10), 2003 => to_unsigned(647, 10), 2004 => to_unsigned(925, 10), 2005 => to_unsigned(394, 10), 2006 => to_unsigned(605, 10), 2007 => to_unsigned(71, 10), 2008 => to_unsigned(496, 10), 2009 => to_unsigned(135, 10), 2010 => to_unsigned(833, 10), 2011 => to_unsigned(409, 10), 2012 => to_unsigned(909, 10), 2013 => to_unsigned(205, 10), 2014 => to_unsigned(192, 10), 2015 => to_unsigned(809, 10), 2016 => to_unsigned(684, 10), 2017 => to_unsigned(147, 10), 2018 => to_unsigned(323, 10), 2019 => to_unsigned(889, 10), 2020 => to_unsigned(167, 10), 2021 => to_unsigned(117, 10), 2022 => to_unsigned(321, 10), 2023 => to_unsigned(81, 10), 2024 => to_unsigned(59, 10), 2025 => to_unsigned(246, 10), 2026 => to_unsigned(738, 10), 2027 => to_unsigned(106, 10), 2028 => to_unsigned(261, 10), 2029 => to_unsigned(834, 10), 2030 => to_unsigned(843, 10), 2031 => to_unsigned(63, 10), 2032 => to_unsigned(747, 10), 2033 => to_unsigned(965, 10), 2034 => to_unsigned(458, 10), 2035 => to_unsigned(1012, 10), 2036 => to_unsigned(644, 10), 2037 => to_unsigned(301, 10), 2038 => to_unsigned(383, 10), 2039 => to_unsigned(288, 10), 2040 => to_unsigned(308, 10), 2041 => to_unsigned(944, 10), 2042 => to_unsigned(723, 10), 2043 => to_unsigned(342, 10), 2044 => to_unsigned(68, 10), 2045 => to_unsigned(405, 10), 2046 => to_unsigned(995, 10), 2047 => to_unsigned(460, 10)),
        2 => (0 => to_unsigned(904, 10), 1 => to_unsigned(350, 10), 2 => to_unsigned(231, 10), 3 => to_unsigned(865, 10), 4 => to_unsigned(651, 10), 5 => to_unsigned(324, 10), 6 => to_unsigned(147, 10), 7 => to_unsigned(879, 10), 8 => to_unsigned(630, 10), 9 => to_unsigned(373, 10), 10 => to_unsigned(955, 10), 11 => to_unsigned(170, 10), 12 => to_unsigned(708, 10), 13 => to_unsigned(886, 10), 14 => to_unsigned(754, 10), 15 => to_unsigned(843, 10), 16 => to_unsigned(343, 10), 17 => to_unsigned(151, 10), 18 => to_unsigned(579, 10), 19 => to_unsigned(820, 10), 20 => to_unsigned(210, 10), 21 => to_unsigned(370, 10), 22 => to_unsigned(51, 10), 23 => to_unsigned(975, 10), 24 => to_unsigned(199, 10), 25 => to_unsigned(324, 10), 26 => to_unsigned(465, 10), 27 => to_unsigned(927, 10), 28 => to_unsigned(985, 10), 29 => to_unsigned(41, 10), 30 => to_unsigned(857, 10), 31 => to_unsigned(806, 10), 32 => to_unsigned(587, 10), 33 => to_unsigned(443, 10), 34 => to_unsigned(879, 10), 35 => to_unsigned(467, 10), 36 => to_unsigned(751, 10), 37 => to_unsigned(593, 10), 38 => to_unsigned(662, 10), 39 => to_unsigned(392, 10), 40 => to_unsigned(961, 10), 41 => to_unsigned(622, 10), 42 => to_unsigned(9, 10), 43 => to_unsigned(53, 10), 44 => to_unsigned(835, 10), 45 => to_unsigned(165, 10), 46 => to_unsigned(857, 10), 47 => to_unsigned(732, 10), 48 => to_unsigned(601, 10), 49 => to_unsigned(622, 10), 50 => to_unsigned(319, 10), 51 => to_unsigned(365, 10), 52 => to_unsigned(767, 10), 53 => to_unsigned(858, 10), 54 => to_unsigned(213, 10), 55 => to_unsigned(671, 10), 56 => to_unsigned(274, 10), 57 => to_unsigned(357, 10), 58 => to_unsigned(489, 10), 59 => to_unsigned(869, 10), 60 => to_unsigned(807, 10), 61 => to_unsigned(970, 10), 62 => to_unsigned(662, 10), 63 => to_unsigned(325, 10), 64 => to_unsigned(836, 10), 65 => to_unsigned(97, 10), 66 => to_unsigned(505, 10), 67 => to_unsigned(744, 10), 68 => to_unsigned(490, 10), 69 => to_unsigned(349, 10), 70 => to_unsigned(300, 10), 71 => to_unsigned(182, 10), 72 => to_unsigned(148, 10), 73 => to_unsigned(965, 10), 74 => to_unsigned(122, 10), 75 => to_unsigned(111, 10), 76 => to_unsigned(655, 10), 77 => to_unsigned(880, 10), 78 => to_unsigned(804, 10), 79 => to_unsigned(29, 10), 80 => to_unsigned(245, 10), 81 => to_unsigned(718, 10), 82 => to_unsigned(239, 10), 83 => to_unsigned(689, 10), 84 => to_unsigned(169, 10), 85 => to_unsigned(116, 10), 86 => to_unsigned(608, 10), 87 => to_unsigned(752, 10), 88 => to_unsigned(730, 10), 89 => to_unsigned(870, 10), 90 => to_unsigned(630, 10), 91 => to_unsigned(379, 10), 92 => to_unsigned(704, 10), 93 => to_unsigned(665, 10), 94 => to_unsigned(26, 10), 95 => to_unsigned(15, 10), 96 => to_unsigned(646, 10), 97 => to_unsigned(292, 10), 98 => to_unsigned(237, 10), 99 => to_unsigned(15, 10), 100 => to_unsigned(263, 10), 101 => to_unsigned(804, 10), 102 => to_unsigned(199, 10), 103 => to_unsigned(93, 10), 104 => to_unsigned(760, 10), 105 => to_unsigned(609, 10), 106 => to_unsigned(582, 10), 107 => to_unsigned(534, 10), 108 => to_unsigned(25, 10), 109 => to_unsigned(99, 10), 110 => to_unsigned(550, 10), 111 => to_unsigned(585, 10), 112 => to_unsigned(457, 10), 113 => to_unsigned(320, 10), 114 => to_unsigned(544, 10), 115 => to_unsigned(109, 10), 116 => to_unsigned(172, 10), 117 => to_unsigned(677, 10), 118 => to_unsigned(92, 10), 119 => to_unsigned(330, 10), 120 => to_unsigned(22, 10), 121 => to_unsigned(200, 10), 122 => to_unsigned(837, 10), 123 => to_unsigned(465, 10), 124 => to_unsigned(787, 10), 125 => to_unsigned(56, 10), 126 => to_unsigned(411, 10), 127 => to_unsigned(562, 10), 128 => to_unsigned(124, 10), 129 => to_unsigned(980, 10), 130 => to_unsigned(334, 10), 131 => to_unsigned(726, 10), 132 => to_unsigned(982, 10), 133 => to_unsigned(909, 10), 134 => to_unsigned(134, 10), 135 => to_unsigned(638, 10), 136 => to_unsigned(223, 10), 137 => to_unsigned(415, 10), 138 => to_unsigned(264, 10), 139 => to_unsigned(202, 10), 140 => to_unsigned(400, 10), 141 => to_unsigned(197, 10), 142 => to_unsigned(976, 10), 143 => to_unsigned(378, 10), 144 => to_unsigned(456, 10), 145 => to_unsigned(842, 10), 146 => to_unsigned(833, 10), 147 => to_unsigned(646, 10), 148 => to_unsigned(652, 10), 149 => to_unsigned(576, 10), 150 => to_unsigned(324, 10), 151 => to_unsigned(447, 10), 152 => to_unsigned(185, 10), 153 => to_unsigned(957, 10), 154 => to_unsigned(319, 10), 155 => to_unsigned(165, 10), 156 => to_unsigned(1017, 10), 157 => to_unsigned(258, 10), 158 => to_unsigned(506, 10), 159 => to_unsigned(427, 10), 160 => to_unsigned(479, 10), 161 => to_unsigned(389, 10), 162 => to_unsigned(57, 10), 163 => to_unsigned(402, 10), 164 => to_unsigned(647, 10), 165 => to_unsigned(233, 10), 166 => to_unsigned(98, 10), 167 => to_unsigned(307, 10), 168 => to_unsigned(205, 10), 169 => to_unsigned(189, 10), 170 => to_unsigned(54, 10), 171 => to_unsigned(19, 10), 172 => to_unsigned(739, 10), 173 => to_unsigned(787, 10), 174 => to_unsigned(466, 10), 175 => to_unsigned(761, 10), 176 => to_unsigned(879, 10), 177 => to_unsigned(1002, 10), 178 => to_unsigned(756, 10), 179 => to_unsigned(991, 10), 180 => to_unsigned(634, 10), 181 => to_unsigned(527, 10), 182 => to_unsigned(981, 10), 183 => to_unsigned(817, 10), 184 => to_unsigned(659, 10), 185 => to_unsigned(507, 10), 186 => to_unsigned(702, 10), 187 => to_unsigned(532, 10), 188 => to_unsigned(126, 10), 189 => to_unsigned(803, 10), 190 => to_unsigned(689, 10), 191 => to_unsigned(906, 10), 192 => to_unsigned(877, 10), 193 => to_unsigned(679, 10), 194 => to_unsigned(12, 10), 195 => to_unsigned(397, 10), 196 => to_unsigned(916, 10), 197 => to_unsigned(245, 10), 198 => to_unsigned(190, 10), 199 => to_unsigned(571, 10), 200 => to_unsigned(178, 10), 201 => to_unsigned(446, 10), 202 => to_unsigned(837, 10), 203 => to_unsigned(852, 10), 204 => to_unsigned(827, 10), 205 => to_unsigned(861, 10), 206 => to_unsigned(941, 10), 207 => to_unsigned(454, 10), 208 => to_unsigned(186, 10), 209 => to_unsigned(857, 10), 210 => to_unsigned(420, 10), 211 => to_unsigned(685, 10), 212 => to_unsigned(451, 10), 213 => to_unsigned(277, 10), 214 => to_unsigned(838, 10), 215 => to_unsigned(838, 10), 216 => to_unsigned(860, 10), 217 => to_unsigned(553, 10), 218 => to_unsigned(934, 10), 219 => to_unsigned(904, 10), 220 => to_unsigned(724, 10), 221 => to_unsigned(784, 10), 222 => to_unsigned(499, 10), 223 => to_unsigned(640, 10), 224 => to_unsigned(749, 10), 225 => to_unsigned(295, 10), 226 => to_unsigned(619, 10), 227 => to_unsigned(453, 10), 228 => to_unsigned(726, 10), 229 => to_unsigned(462, 10), 230 => to_unsigned(678, 10), 231 => to_unsigned(396, 10), 232 => to_unsigned(237, 10), 233 => to_unsigned(621, 10), 234 => to_unsigned(719, 10), 235 => to_unsigned(316, 10), 236 => to_unsigned(943, 10), 237 => to_unsigned(86, 10), 238 => to_unsigned(259, 10), 239 => to_unsigned(566, 10), 240 => to_unsigned(63, 10), 241 => to_unsigned(914, 10), 242 => to_unsigned(553, 10), 243 => to_unsigned(523, 10), 244 => to_unsigned(500, 10), 245 => to_unsigned(10, 10), 246 => to_unsigned(145, 10), 247 => to_unsigned(974, 10), 248 => to_unsigned(697, 10), 249 => to_unsigned(869, 10), 250 => to_unsigned(211, 10), 251 => to_unsigned(988, 10), 252 => to_unsigned(88, 10), 253 => to_unsigned(826, 10), 254 => to_unsigned(213, 10), 255 => to_unsigned(1001, 10), 256 => to_unsigned(770, 10), 257 => to_unsigned(812, 10), 258 => to_unsigned(391, 10), 259 => to_unsigned(746, 10), 260 => to_unsigned(760, 10), 261 => to_unsigned(1018, 10), 262 => to_unsigned(325, 10), 263 => to_unsigned(761, 10), 264 => to_unsigned(871, 10), 265 => to_unsigned(840, 10), 266 => to_unsigned(183, 10), 267 => to_unsigned(685, 10), 268 => to_unsigned(354, 10), 269 => to_unsigned(652, 10), 270 => to_unsigned(798, 10), 271 => to_unsigned(322, 10), 272 => to_unsigned(242, 10), 273 => to_unsigned(210, 10), 274 => to_unsigned(273, 10), 275 => to_unsigned(507, 10), 276 => to_unsigned(952, 10), 277 => to_unsigned(199, 10), 278 => to_unsigned(931, 10), 279 => to_unsigned(396, 10), 280 => to_unsigned(554, 10), 281 => to_unsigned(1017, 10), 282 => to_unsigned(190, 10), 283 => to_unsigned(404, 10), 284 => to_unsigned(641, 10), 285 => to_unsigned(519, 10), 286 => to_unsigned(766, 10), 287 => to_unsigned(438, 10), 288 => to_unsigned(719, 10), 289 => to_unsigned(925, 10), 290 => to_unsigned(253, 10), 291 => to_unsigned(452, 10), 292 => to_unsigned(140, 10), 293 => to_unsigned(839, 10), 294 => to_unsigned(71, 10), 295 => to_unsigned(819, 10), 296 => to_unsigned(498, 10), 297 => to_unsigned(618, 10), 298 => to_unsigned(908, 10), 299 => to_unsigned(708, 10), 300 => to_unsigned(778, 10), 301 => to_unsigned(1020, 10), 302 => to_unsigned(447, 10), 303 => to_unsigned(126, 10), 304 => to_unsigned(251, 10), 305 => to_unsigned(119, 10), 306 => to_unsigned(315, 10), 307 => to_unsigned(735, 10), 308 => to_unsigned(525, 10), 309 => to_unsigned(88, 10), 310 => to_unsigned(471, 10), 311 => to_unsigned(123, 10), 312 => to_unsigned(300, 10), 313 => to_unsigned(522, 10), 314 => to_unsigned(213, 10), 315 => to_unsigned(746, 10), 316 => to_unsigned(1000, 10), 317 => to_unsigned(889, 10), 318 => to_unsigned(242, 10), 319 => to_unsigned(902, 10), 320 => to_unsigned(980, 10), 321 => to_unsigned(556, 10), 322 => to_unsigned(260, 10), 323 => to_unsigned(351, 10), 324 => to_unsigned(863, 10), 325 => to_unsigned(871, 10), 326 => to_unsigned(988, 10), 327 => to_unsigned(16, 10), 328 => to_unsigned(577, 10), 329 => to_unsigned(747, 10), 330 => to_unsigned(992, 10), 331 => to_unsigned(194, 10), 332 => to_unsigned(119, 10), 333 => to_unsigned(157, 10), 334 => to_unsigned(330, 10), 335 => to_unsigned(152, 10), 336 => to_unsigned(776, 10), 337 => to_unsigned(815, 10), 338 => to_unsigned(94, 10), 339 => to_unsigned(793, 10), 340 => to_unsigned(521, 10), 341 => to_unsigned(328, 10), 342 => to_unsigned(764, 10), 343 => to_unsigned(759, 10), 344 => to_unsigned(195, 10), 345 => to_unsigned(170, 10), 346 => to_unsigned(485, 10), 347 => to_unsigned(269, 10), 348 => to_unsigned(31, 10), 349 => to_unsigned(46, 10), 350 => to_unsigned(661, 10), 351 => to_unsigned(384, 10), 352 => to_unsigned(637, 10), 353 => to_unsigned(963, 10), 354 => to_unsigned(763, 10), 355 => to_unsigned(826, 10), 356 => to_unsigned(838, 10), 357 => to_unsigned(460, 10), 358 => to_unsigned(856, 10), 359 => to_unsigned(382, 10), 360 => to_unsigned(309, 10), 361 => to_unsigned(15, 10), 362 => to_unsigned(900, 10), 363 => to_unsigned(440, 10), 364 => to_unsigned(393, 10), 365 => to_unsigned(541, 10), 366 => to_unsigned(29, 10), 367 => to_unsigned(538, 10), 368 => to_unsigned(4, 10), 369 => to_unsigned(155, 10), 370 => to_unsigned(541, 10), 371 => to_unsigned(400, 10), 372 => to_unsigned(112, 10), 373 => to_unsigned(270, 10), 374 => to_unsigned(900, 10), 375 => to_unsigned(585, 10), 376 => to_unsigned(462, 10), 377 => to_unsigned(267, 10), 378 => to_unsigned(23, 10), 379 => to_unsigned(754, 10), 380 => to_unsigned(246, 10), 381 => to_unsigned(88, 10), 382 => to_unsigned(149, 10), 383 => to_unsigned(617, 10), 384 => to_unsigned(193, 10), 385 => to_unsigned(32, 10), 386 => to_unsigned(716, 10), 387 => to_unsigned(512, 10), 388 => to_unsigned(479, 10), 389 => to_unsigned(36, 10), 390 => to_unsigned(667, 10), 391 => to_unsigned(516, 10), 392 => to_unsigned(572, 10), 393 => to_unsigned(950, 10), 394 => to_unsigned(111, 10), 395 => to_unsigned(294, 10), 396 => to_unsigned(434, 10), 397 => to_unsigned(418, 10), 398 => to_unsigned(323, 10), 399 => to_unsigned(595, 10), 400 => to_unsigned(358, 10), 401 => to_unsigned(996, 10), 402 => to_unsigned(565, 10), 403 => to_unsigned(445, 10), 404 => to_unsigned(881, 10), 405 => to_unsigned(379, 10), 406 => to_unsigned(467, 10), 407 => to_unsigned(772, 10), 408 => to_unsigned(857, 10), 409 => to_unsigned(341, 10), 410 => to_unsigned(995, 10), 411 => to_unsigned(932, 10), 412 => to_unsigned(477, 10), 413 => to_unsigned(274, 10), 414 => to_unsigned(257, 10), 415 => to_unsigned(955, 10), 416 => to_unsigned(154, 10), 417 => to_unsigned(628, 10), 418 => to_unsigned(285, 10), 419 => to_unsigned(664, 10), 420 => to_unsigned(54, 10), 421 => to_unsigned(450, 10), 422 => to_unsigned(49, 10), 423 => to_unsigned(219, 10), 424 => to_unsigned(690, 10), 425 => to_unsigned(888, 10), 426 => to_unsigned(877, 10), 427 => to_unsigned(93, 10), 428 => to_unsigned(122, 10), 429 => to_unsigned(331, 10), 430 => to_unsigned(566, 10), 431 => to_unsigned(512, 10), 432 => to_unsigned(712, 10), 433 => to_unsigned(219, 10), 434 => to_unsigned(264, 10), 435 => to_unsigned(678, 10), 436 => to_unsigned(746, 10), 437 => to_unsigned(692, 10), 438 => to_unsigned(336, 10), 439 => to_unsigned(653, 10), 440 => to_unsigned(696, 10), 441 => to_unsigned(675, 10), 442 => to_unsigned(155, 10), 443 => to_unsigned(23, 10), 444 => to_unsigned(943, 10), 445 => to_unsigned(885, 10), 446 => to_unsigned(911, 10), 447 => to_unsigned(178, 10), 448 => to_unsigned(888, 10), 449 => to_unsigned(317, 10), 450 => to_unsigned(648, 10), 451 => to_unsigned(721, 10), 452 => to_unsigned(464, 10), 453 => to_unsigned(920, 10), 454 => to_unsigned(244, 10), 455 => to_unsigned(567, 10), 456 => to_unsigned(270, 10), 457 => to_unsigned(336, 10), 458 => to_unsigned(840, 10), 459 => to_unsigned(761, 10), 460 => to_unsigned(571, 10), 461 => to_unsigned(87, 10), 462 => to_unsigned(917, 10), 463 => to_unsigned(202, 10), 464 => to_unsigned(929, 10), 465 => to_unsigned(824, 10), 466 => to_unsigned(992, 10), 467 => to_unsigned(549, 10), 468 => to_unsigned(742, 10), 469 => to_unsigned(110, 10), 470 => to_unsigned(975, 10), 471 => to_unsigned(433, 10), 472 => to_unsigned(617, 10), 473 => to_unsigned(204, 10), 474 => to_unsigned(178, 10), 475 => to_unsigned(593, 10), 476 => to_unsigned(459, 10), 477 => to_unsigned(804, 10), 478 => to_unsigned(824, 10), 479 => to_unsigned(154, 10), 480 => to_unsigned(730, 10), 481 => to_unsigned(635, 10), 482 => to_unsigned(613, 10), 483 => to_unsigned(937, 10), 484 => to_unsigned(534, 10), 485 => to_unsigned(454, 10), 486 => to_unsigned(660, 10), 487 => to_unsigned(826, 10), 488 => to_unsigned(395, 10), 489 => to_unsigned(808, 10), 490 => to_unsigned(193, 10), 491 => to_unsigned(62, 10), 492 => to_unsigned(281, 10), 493 => to_unsigned(456, 10), 494 => to_unsigned(1001, 10), 495 => to_unsigned(196, 10), 496 => to_unsigned(635, 10), 497 => to_unsigned(127, 10), 498 => to_unsigned(619, 10), 499 => to_unsigned(570, 10), 500 => to_unsigned(389, 10), 501 => to_unsigned(834, 10), 502 => to_unsigned(692, 10), 503 => to_unsigned(727, 10), 504 => to_unsigned(204, 10), 505 => to_unsigned(442, 10), 506 => to_unsigned(340, 10), 507 => to_unsigned(696, 10), 508 => to_unsigned(125, 10), 509 => to_unsigned(61, 10), 510 => to_unsigned(894, 10), 511 => to_unsigned(296, 10), 512 => to_unsigned(237, 10), 513 => to_unsigned(190, 10), 514 => to_unsigned(971, 10), 515 => to_unsigned(919, 10), 516 => to_unsigned(896, 10), 517 => to_unsigned(873, 10), 518 => to_unsigned(755, 10), 519 => to_unsigned(346, 10), 520 => to_unsigned(729, 10), 521 => to_unsigned(164, 10), 522 => to_unsigned(430, 10), 523 => to_unsigned(313, 10), 524 => to_unsigned(1023, 10), 525 => to_unsigned(541, 10), 526 => to_unsigned(233, 10), 527 => to_unsigned(533, 10), 528 => to_unsigned(650, 10), 529 => to_unsigned(503, 10), 530 => to_unsigned(884, 10), 531 => to_unsigned(976, 10), 532 => to_unsigned(752, 10), 533 => to_unsigned(473, 10), 534 => to_unsigned(769, 10), 535 => to_unsigned(114, 10), 536 => to_unsigned(365, 10), 537 => to_unsigned(307, 10), 538 => to_unsigned(170, 10), 539 => to_unsigned(649, 10), 540 => to_unsigned(1010, 10), 541 => to_unsigned(70, 10), 542 => to_unsigned(181, 10), 543 => to_unsigned(70, 10), 544 => to_unsigned(267, 10), 545 => to_unsigned(577, 10), 546 => to_unsigned(199, 10), 547 => to_unsigned(340, 10), 548 => to_unsigned(105, 10), 549 => to_unsigned(739, 10), 550 => to_unsigned(807, 10), 551 => to_unsigned(494, 10), 552 => to_unsigned(642, 10), 553 => to_unsigned(547, 10), 554 => to_unsigned(129, 10), 555 => to_unsigned(651, 10), 556 => to_unsigned(912, 10), 557 => to_unsigned(249, 10), 558 => to_unsigned(990, 10), 559 => to_unsigned(943, 10), 560 => to_unsigned(400, 10), 561 => to_unsigned(978, 10), 562 => to_unsigned(747, 10), 563 => to_unsigned(1017, 10), 564 => to_unsigned(485, 10), 565 => to_unsigned(331, 10), 566 => to_unsigned(315, 10), 567 => to_unsigned(729, 10), 568 => to_unsigned(536, 10), 569 => to_unsigned(446, 10), 570 => to_unsigned(233, 10), 571 => to_unsigned(107, 10), 572 => to_unsigned(281, 10), 573 => to_unsigned(218, 10), 574 => to_unsigned(1012, 10), 575 => to_unsigned(145, 10), 576 => to_unsigned(41, 10), 577 => to_unsigned(342, 10), 578 => to_unsigned(910, 10), 579 => to_unsigned(324, 10), 580 => to_unsigned(531, 10), 581 => to_unsigned(715, 10), 582 => to_unsigned(607, 10), 583 => to_unsigned(371, 10), 584 => to_unsigned(756, 10), 585 => to_unsigned(133, 10), 586 => to_unsigned(357, 10), 587 => to_unsigned(757, 10), 588 => to_unsigned(816, 10), 589 => to_unsigned(451, 10), 590 => to_unsigned(609, 10), 591 => to_unsigned(497, 10), 592 => to_unsigned(622, 10), 593 => to_unsigned(760, 10), 594 => to_unsigned(497, 10), 595 => to_unsigned(30, 10), 596 => to_unsigned(386, 10), 597 => to_unsigned(870, 10), 598 => to_unsigned(311, 10), 599 => to_unsigned(438, 10), 600 => to_unsigned(55, 10), 601 => to_unsigned(24, 10), 602 => to_unsigned(503, 10), 603 => to_unsigned(14, 10), 604 => to_unsigned(769, 10), 605 => to_unsigned(950, 10), 606 => to_unsigned(180, 10), 607 => to_unsigned(660, 10), 608 => to_unsigned(661, 10), 609 => to_unsigned(327, 10), 610 => to_unsigned(406, 10), 611 => to_unsigned(89, 10), 612 => to_unsigned(900, 10), 613 => to_unsigned(507, 10), 614 => to_unsigned(336, 10), 615 => to_unsigned(501, 10), 616 => to_unsigned(39, 10), 617 => to_unsigned(534, 10), 618 => to_unsigned(300, 10), 619 => to_unsigned(616, 10), 620 => to_unsigned(616, 10), 621 => to_unsigned(680, 10), 622 => to_unsigned(577, 10), 623 => to_unsigned(968, 10), 624 => to_unsigned(115, 10), 625 => to_unsigned(42, 10), 626 => to_unsigned(245, 10), 627 => to_unsigned(648, 10), 628 => to_unsigned(439, 10), 629 => to_unsigned(455, 10), 630 => to_unsigned(319, 10), 631 => to_unsigned(540, 10), 632 => to_unsigned(616, 10), 633 => to_unsigned(358, 10), 634 => to_unsigned(516, 10), 635 => to_unsigned(340, 10), 636 => to_unsigned(611, 10), 637 => to_unsigned(438, 10), 638 => to_unsigned(491, 10), 639 => to_unsigned(628, 10), 640 => to_unsigned(250, 10), 641 => to_unsigned(839, 10), 642 => to_unsigned(937, 10), 643 => to_unsigned(205, 10), 644 => to_unsigned(957, 10), 645 => to_unsigned(568, 10), 646 => to_unsigned(659, 10), 647 => to_unsigned(32, 10), 648 => to_unsigned(73, 10), 649 => to_unsigned(94, 10), 650 => to_unsigned(631, 10), 651 => to_unsigned(933, 10), 652 => to_unsigned(108, 10), 653 => to_unsigned(383, 10), 654 => to_unsigned(845, 10), 655 => to_unsigned(238, 10), 656 => to_unsigned(350, 10), 657 => to_unsigned(833, 10), 658 => to_unsigned(588, 10), 659 => to_unsigned(1014, 10), 660 => to_unsigned(132, 10), 661 => to_unsigned(89, 10), 662 => to_unsigned(362, 10), 663 => to_unsigned(27, 10), 664 => to_unsigned(9, 10), 665 => to_unsigned(72, 10), 666 => to_unsigned(445, 10), 667 => to_unsigned(355, 10), 668 => to_unsigned(408, 10), 669 => to_unsigned(481, 10), 670 => to_unsigned(521, 10), 671 => to_unsigned(383, 10), 672 => to_unsigned(113, 10), 673 => to_unsigned(580, 10), 674 => to_unsigned(785, 10), 675 => to_unsigned(1010, 10), 676 => to_unsigned(490, 10), 677 => to_unsigned(66, 10), 678 => to_unsigned(917, 10), 679 => to_unsigned(118, 10), 680 => to_unsigned(267, 10), 681 => to_unsigned(610, 10), 682 => to_unsigned(796, 10), 683 => to_unsigned(125, 10), 684 => to_unsigned(989, 10), 685 => to_unsigned(483, 10), 686 => to_unsigned(660, 10), 687 => to_unsigned(67, 10), 688 => to_unsigned(191, 10), 689 => to_unsigned(926, 10), 690 => to_unsigned(496, 10), 691 => to_unsigned(156, 10), 692 => to_unsigned(741, 10), 693 => to_unsigned(474, 10), 694 => to_unsigned(724, 10), 695 => to_unsigned(35, 10), 696 => to_unsigned(690, 10), 697 => to_unsigned(558, 10), 698 => to_unsigned(83, 10), 699 => to_unsigned(413, 10), 700 => to_unsigned(738, 10), 701 => to_unsigned(606, 10), 702 => to_unsigned(48, 10), 703 => to_unsigned(284, 10), 704 => to_unsigned(975, 10), 705 => to_unsigned(164, 10), 706 => to_unsigned(625, 10), 707 => to_unsigned(778, 10), 708 => to_unsigned(965, 10), 709 => to_unsigned(659, 10), 710 => to_unsigned(130, 10), 711 => to_unsigned(381, 10), 712 => to_unsigned(241, 10), 713 => to_unsigned(710, 10), 714 => to_unsigned(960, 10), 715 => to_unsigned(57, 10), 716 => to_unsigned(158, 10), 717 => to_unsigned(900, 10), 718 => to_unsigned(512, 10), 719 => to_unsigned(854, 10), 720 => to_unsigned(983, 10), 721 => to_unsigned(10, 10), 722 => to_unsigned(902, 10), 723 => to_unsigned(958, 10), 724 => to_unsigned(992, 10), 725 => to_unsigned(323, 10), 726 => to_unsigned(548, 10), 727 => to_unsigned(737, 10), 728 => to_unsigned(638, 10), 729 => to_unsigned(224, 10), 730 => to_unsigned(6, 10), 731 => to_unsigned(709, 10), 732 => to_unsigned(101, 10), 733 => to_unsigned(831, 10), 734 => to_unsigned(79, 10), 735 => to_unsigned(483, 10), 736 => to_unsigned(857, 10), 737 => to_unsigned(19, 10), 738 => to_unsigned(385, 10), 739 => to_unsigned(1003, 10), 740 => to_unsigned(536, 10), 741 => to_unsigned(630, 10), 742 => to_unsigned(213, 10), 743 => to_unsigned(226, 10), 744 => to_unsigned(654, 10), 745 => to_unsigned(628, 10), 746 => to_unsigned(386, 10), 747 => to_unsigned(583, 10), 748 => to_unsigned(101, 10), 749 => to_unsigned(279, 10), 750 => to_unsigned(694, 10), 751 => to_unsigned(422, 10), 752 => to_unsigned(287, 10), 753 => to_unsigned(705, 10), 754 => to_unsigned(1023, 10), 755 => to_unsigned(103, 10), 756 => to_unsigned(443, 10), 757 => to_unsigned(762, 10), 758 => to_unsigned(17, 10), 759 => to_unsigned(52, 10), 760 => to_unsigned(461, 10), 761 => to_unsigned(798, 10), 762 => to_unsigned(867, 10), 763 => to_unsigned(313, 10), 764 => to_unsigned(854, 10), 765 => to_unsigned(211, 10), 766 => to_unsigned(251, 10), 767 => to_unsigned(412, 10), 768 => to_unsigned(326, 10), 769 => to_unsigned(193, 10), 770 => to_unsigned(505, 10), 771 => to_unsigned(5, 10), 772 => to_unsigned(523, 10), 773 => to_unsigned(53, 10), 774 => to_unsigned(920, 10), 775 => to_unsigned(346, 10), 776 => to_unsigned(760, 10), 777 => to_unsigned(815, 10), 778 => to_unsigned(321, 10), 779 => to_unsigned(869, 10), 780 => to_unsigned(682, 10), 781 => to_unsigned(447, 10), 782 => to_unsigned(160, 10), 783 => to_unsigned(523, 10), 784 => to_unsigned(914, 10), 785 => to_unsigned(639, 10), 786 => to_unsigned(536, 10), 787 => to_unsigned(132, 10), 788 => to_unsigned(903, 10), 789 => to_unsigned(544, 10), 790 => to_unsigned(399, 10), 791 => to_unsigned(1, 10), 792 => to_unsigned(369, 10), 793 => to_unsigned(88, 10), 794 => to_unsigned(933, 10), 795 => to_unsigned(886, 10), 796 => to_unsigned(593, 10), 797 => to_unsigned(372, 10), 798 => to_unsigned(31, 10), 799 => to_unsigned(927, 10), 800 => to_unsigned(456, 10), 801 => to_unsigned(961, 10), 802 => to_unsigned(372, 10), 803 => to_unsigned(753, 10), 804 => to_unsigned(52, 10), 805 => to_unsigned(256, 10), 806 => to_unsigned(669, 10), 807 => to_unsigned(824, 10), 808 => to_unsigned(897, 10), 809 => to_unsigned(153, 10), 810 => to_unsigned(745, 10), 811 => to_unsigned(834, 10), 812 => to_unsigned(44, 10), 813 => to_unsigned(786, 10), 814 => to_unsigned(724, 10), 815 => to_unsigned(231, 10), 816 => to_unsigned(993, 10), 817 => to_unsigned(509, 10), 818 => to_unsigned(819, 10), 819 => to_unsigned(845, 10), 820 => to_unsigned(287, 10), 821 => to_unsigned(885, 10), 822 => to_unsigned(132, 10), 823 => to_unsigned(680, 10), 824 => to_unsigned(995, 10), 825 => to_unsigned(376, 10), 826 => to_unsigned(119, 10), 827 => to_unsigned(883, 10), 828 => to_unsigned(610, 10), 829 => to_unsigned(382, 10), 830 => to_unsigned(407, 10), 831 => to_unsigned(606, 10), 832 => to_unsigned(312, 10), 833 => to_unsigned(441, 10), 834 => to_unsigned(829, 10), 835 => to_unsigned(3, 10), 836 => to_unsigned(333, 10), 837 => to_unsigned(686, 10), 838 => to_unsigned(283, 10), 839 => to_unsigned(494, 10), 840 => to_unsigned(96, 10), 841 => to_unsigned(257, 10), 842 => to_unsigned(3, 10), 843 => to_unsigned(98, 10), 844 => to_unsigned(740, 10), 845 => to_unsigned(267, 10), 846 => to_unsigned(699, 10), 847 => to_unsigned(103, 10), 848 => to_unsigned(470, 10), 849 => to_unsigned(401, 10), 850 => to_unsigned(156, 10), 851 => to_unsigned(679, 10), 852 => to_unsigned(66, 10), 853 => to_unsigned(820, 10), 854 => to_unsigned(857, 10), 855 => to_unsigned(656, 10), 856 => to_unsigned(684, 10), 857 => to_unsigned(623, 10), 858 => to_unsigned(752, 10), 859 => to_unsigned(118, 10), 860 => to_unsigned(343, 10), 861 => to_unsigned(245, 10), 862 => to_unsigned(746, 10), 863 => to_unsigned(132, 10), 864 => to_unsigned(844, 10), 865 => to_unsigned(455, 10), 866 => to_unsigned(1002, 10), 867 => to_unsigned(535, 10), 868 => to_unsigned(88, 10), 869 => to_unsigned(447, 10), 870 => to_unsigned(209, 10), 871 => to_unsigned(756, 10), 872 => to_unsigned(939, 10), 873 => to_unsigned(732, 10), 874 => to_unsigned(453, 10), 875 => to_unsigned(362, 10), 876 => to_unsigned(342, 10), 877 => to_unsigned(912, 10), 878 => to_unsigned(815, 10), 879 => to_unsigned(1018, 10), 880 => to_unsigned(617, 10), 881 => to_unsigned(642, 10), 882 => to_unsigned(709, 10), 883 => to_unsigned(683, 10), 884 => to_unsigned(406, 10), 885 => to_unsigned(753, 10), 886 => to_unsigned(275, 10), 887 => to_unsigned(724, 10), 888 => to_unsigned(550, 10), 889 => to_unsigned(338, 10), 890 => to_unsigned(649, 10), 891 => to_unsigned(87, 10), 892 => to_unsigned(835, 10), 893 => to_unsigned(430, 10), 894 => to_unsigned(134, 10), 895 => to_unsigned(140, 10), 896 => to_unsigned(235, 10), 897 => to_unsigned(137, 10), 898 => to_unsigned(26, 10), 899 => to_unsigned(1005, 10), 900 => to_unsigned(457, 10), 901 => to_unsigned(651, 10), 902 => to_unsigned(453, 10), 903 => to_unsigned(256, 10), 904 => to_unsigned(967, 10), 905 => to_unsigned(438, 10), 906 => to_unsigned(829, 10), 907 => to_unsigned(469, 10), 908 => to_unsigned(713, 10), 909 => to_unsigned(412, 10), 910 => to_unsigned(80, 10), 911 => to_unsigned(46, 10), 912 => to_unsigned(308, 10), 913 => to_unsigned(980, 10), 914 => to_unsigned(635, 10), 915 => to_unsigned(808, 10), 916 => to_unsigned(885, 10), 917 => to_unsigned(606, 10), 918 => to_unsigned(526, 10), 919 => to_unsigned(552, 10), 920 => to_unsigned(980, 10), 921 => to_unsigned(385, 10), 922 => to_unsigned(684, 10), 923 => to_unsigned(540, 10), 924 => to_unsigned(505, 10), 925 => to_unsigned(395, 10), 926 => to_unsigned(997, 10), 927 => to_unsigned(701, 10), 928 => to_unsigned(507, 10), 929 => to_unsigned(706, 10), 930 => to_unsigned(289, 10), 931 => to_unsigned(635, 10), 932 => to_unsigned(536, 10), 933 => to_unsigned(260, 10), 934 => to_unsigned(932, 10), 935 => to_unsigned(178, 10), 936 => to_unsigned(828, 10), 937 => to_unsigned(92, 10), 938 => to_unsigned(645, 10), 939 => to_unsigned(989, 10), 940 => to_unsigned(434, 10), 941 => to_unsigned(599, 10), 942 => to_unsigned(293, 10), 943 => to_unsigned(519, 10), 944 => to_unsigned(718, 10), 945 => to_unsigned(96, 10), 946 => to_unsigned(866, 10), 947 => to_unsigned(621, 10), 948 => to_unsigned(707, 10), 949 => to_unsigned(360, 10), 950 => to_unsigned(966, 10), 951 => to_unsigned(100, 10), 952 => to_unsigned(748, 10), 953 => to_unsigned(929, 10), 954 => to_unsigned(446, 10), 955 => to_unsigned(572, 10), 956 => to_unsigned(244, 10), 957 => to_unsigned(389, 10), 958 => to_unsigned(644, 10), 959 => to_unsigned(363, 10), 960 => to_unsigned(172, 10), 961 => to_unsigned(916, 10), 962 => to_unsigned(34, 10), 963 => to_unsigned(313, 10), 964 => to_unsigned(1019, 10), 965 => to_unsigned(126, 10), 966 => to_unsigned(352, 10), 967 => to_unsigned(626, 10), 968 => to_unsigned(151, 10), 969 => to_unsigned(340, 10), 970 => to_unsigned(780, 10), 971 => to_unsigned(501, 10), 972 => to_unsigned(88, 10), 973 => to_unsigned(142, 10), 974 => to_unsigned(462, 10), 975 => to_unsigned(378, 10), 976 => to_unsigned(534, 10), 977 => to_unsigned(134, 10), 978 => to_unsigned(1017, 10), 979 => to_unsigned(868, 10), 980 => to_unsigned(188, 10), 981 => to_unsigned(509, 10), 982 => to_unsigned(241, 10), 983 => to_unsigned(758, 10), 984 => to_unsigned(372, 10), 985 => to_unsigned(812, 10), 986 => to_unsigned(852, 10), 987 => to_unsigned(619, 10), 988 => to_unsigned(648, 10), 989 => to_unsigned(379, 10), 990 => to_unsigned(315, 10), 991 => to_unsigned(575, 10), 992 => to_unsigned(468, 10), 993 => to_unsigned(200, 10), 994 => to_unsigned(322, 10), 995 => to_unsigned(803, 10), 996 => to_unsigned(441, 10), 997 => to_unsigned(461, 10), 998 => to_unsigned(233, 10), 999 => to_unsigned(332, 10), 1000 => to_unsigned(1005, 10), 1001 => to_unsigned(370, 10), 1002 => to_unsigned(825, 10), 1003 => to_unsigned(562, 10), 1004 => to_unsigned(278, 10), 1005 => to_unsigned(132, 10), 1006 => to_unsigned(42, 10), 1007 => to_unsigned(954, 10), 1008 => to_unsigned(42, 10), 1009 => to_unsigned(488, 10), 1010 => to_unsigned(493, 10), 1011 => to_unsigned(875, 10), 1012 => to_unsigned(544, 10), 1013 => to_unsigned(374, 10), 1014 => to_unsigned(965, 10), 1015 => to_unsigned(619, 10), 1016 => to_unsigned(136, 10), 1017 => to_unsigned(704, 10), 1018 => to_unsigned(303, 10), 1019 => to_unsigned(348, 10), 1020 => to_unsigned(695, 10), 1021 => to_unsigned(856, 10), 1022 => to_unsigned(916, 10), 1023 => to_unsigned(267, 10), 1024 => to_unsigned(385, 10), 1025 => to_unsigned(601, 10), 1026 => to_unsigned(311, 10), 1027 => to_unsigned(879, 10), 1028 => to_unsigned(37, 10), 1029 => to_unsigned(928, 10), 1030 => to_unsigned(305, 10), 1031 => to_unsigned(75, 10), 1032 => to_unsigned(325, 10), 1033 => to_unsigned(400, 10), 1034 => to_unsigned(808, 10), 1035 => to_unsigned(908, 10), 1036 => to_unsigned(496, 10), 1037 => to_unsigned(983, 10), 1038 => to_unsigned(235, 10), 1039 => to_unsigned(601, 10), 1040 => to_unsigned(680, 10), 1041 => to_unsigned(234, 10), 1042 => to_unsigned(833, 10), 1043 => to_unsigned(217, 10), 1044 => to_unsigned(918, 10), 1045 => to_unsigned(321, 10), 1046 => to_unsigned(183, 10), 1047 => to_unsigned(333, 10), 1048 => to_unsigned(149, 10), 1049 => to_unsigned(358, 10), 1050 => to_unsigned(124, 10), 1051 => to_unsigned(163, 10), 1052 => to_unsigned(314, 10), 1053 => to_unsigned(608, 10), 1054 => to_unsigned(143, 10), 1055 => to_unsigned(630, 10), 1056 => to_unsigned(711, 10), 1057 => to_unsigned(695, 10), 1058 => to_unsigned(393, 10), 1059 => to_unsigned(969, 10), 1060 => to_unsigned(793, 10), 1061 => to_unsigned(255, 10), 1062 => to_unsigned(754, 10), 1063 => to_unsigned(731, 10), 1064 => to_unsigned(693, 10), 1065 => to_unsigned(984, 10), 1066 => to_unsigned(738, 10), 1067 => to_unsigned(429, 10), 1068 => to_unsigned(920, 10), 1069 => to_unsigned(847, 10), 1070 => to_unsigned(514, 10), 1071 => to_unsigned(300, 10), 1072 => to_unsigned(511, 10), 1073 => to_unsigned(382, 10), 1074 => to_unsigned(772, 10), 1075 => to_unsigned(391, 10), 1076 => to_unsigned(25, 10), 1077 => to_unsigned(974, 10), 1078 => to_unsigned(925, 10), 1079 => to_unsigned(341, 10), 1080 => to_unsigned(332, 10), 1081 => to_unsigned(658, 10), 1082 => to_unsigned(502, 10), 1083 => to_unsigned(752, 10), 1084 => to_unsigned(494, 10), 1085 => to_unsigned(523, 10), 1086 => to_unsigned(869, 10), 1087 => to_unsigned(11, 10), 1088 => to_unsigned(513, 10), 1089 => to_unsigned(207, 10), 1090 => to_unsigned(756, 10), 1091 => to_unsigned(912, 10), 1092 => to_unsigned(411, 10), 1093 => to_unsigned(717, 10), 1094 => to_unsigned(679, 10), 1095 => to_unsigned(543, 10), 1096 => to_unsigned(356, 10), 1097 => to_unsigned(713, 10), 1098 => to_unsigned(679, 10), 1099 => to_unsigned(209, 10), 1100 => to_unsigned(814, 10), 1101 => to_unsigned(584, 10), 1102 => to_unsigned(548, 10), 1103 => to_unsigned(290, 10), 1104 => to_unsigned(171, 10), 1105 => to_unsigned(775, 10), 1106 => to_unsigned(122, 10), 1107 => to_unsigned(675, 10), 1108 => to_unsigned(890, 10), 1109 => to_unsigned(409, 10), 1110 => to_unsigned(395, 10), 1111 => to_unsigned(34, 10), 1112 => to_unsigned(535, 10), 1113 => to_unsigned(103, 10), 1114 => to_unsigned(444, 10), 1115 => to_unsigned(401, 10), 1116 => to_unsigned(689, 10), 1117 => to_unsigned(692, 10), 1118 => to_unsigned(981, 10), 1119 => to_unsigned(474, 10), 1120 => to_unsigned(110, 10), 1121 => to_unsigned(762, 10), 1122 => to_unsigned(203, 10), 1123 => to_unsigned(889, 10), 1124 => to_unsigned(34, 10), 1125 => to_unsigned(246, 10), 1126 => to_unsigned(130, 10), 1127 => to_unsigned(73, 10), 1128 => to_unsigned(367, 10), 1129 => to_unsigned(420, 10), 1130 => to_unsigned(637, 10), 1131 => to_unsigned(385, 10), 1132 => to_unsigned(186, 10), 1133 => to_unsigned(319, 10), 1134 => to_unsigned(311, 10), 1135 => to_unsigned(573, 10), 1136 => to_unsigned(457, 10), 1137 => to_unsigned(811, 10), 1138 => to_unsigned(843, 10), 1139 => to_unsigned(788, 10), 1140 => to_unsigned(773, 10), 1141 => to_unsigned(36, 10), 1142 => to_unsigned(619, 10), 1143 => to_unsigned(56, 10), 1144 => to_unsigned(979, 10), 1145 => to_unsigned(950, 10), 1146 => to_unsigned(711, 10), 1147 => to_unsigned(946, 10), 1148 => to_unsigned(826, 10), 1149 => to_unsigned(931, 10), 1150 => to_unsigned(6, 10), 1151 => to_unsigned(545, 10), 1152 => to_unsigned(216, 10), 1153 => to_unsigned(259, 10), 1154 => to_unsigned(729, 10), 1155 => to_unsigned(657, 10), 1156 => to_unsigned(744, 10), 1157 => to_unsigned(943, 10), 1158 => to_unsigned(588, 10), 1159 => to_unsigned(1004, 10), 1160 => to_unsigned(751, 10), 1161 => to_unsigned(305, 10), 1162 => to_unsigned(565, 10), 1163 => to_unsigned(523, 10), 1164 => to_unsigned(648, 10), 1165 => to_unsigned(1014, 10), 1166 => to_unsigned(733, 10), 1167 => to_unsigned(817, 10), 1168 => to_unsigned(536, 10), 1169 => to_unsigned(668, 10), 1170 => to_unsigned(288, 10), 1171 => to_unsigned(339, 10), 1172 => to_unsigned(302, 10), 1173 => to_unsigned(840, 10), 1174 => to_unsigned(888, 10), 1175 => to_unsigned(345, 10), 1176 => to_unsigned(144, 10), 1177 => to_unsigned(460, 10), 1178 => to_unsigned(246, 10), 1179 => to_unsigned(366, 10), 1180 => to_unsigned(163, 10), 1181 => to_unsigned(894, 10), 1182 => to_unsigned(235, 10), 1183 => to_unsigned(126, 10), 1184 => to_unsigned(615, 10), 1185 => to_unsigned(312, 10), 1186 => to_unsigned(547, 10), 1187 => to_unsigned(29, 10), 1188 => to_unsigned(846, 10), 1189 => to_unsigned(717, 10), 1190 => to_unsigned(109, 10), 1191 => to_unsigned(394, 10), 1192 => to_unsigned(912, 10), 1193 => to_unsigned(387, 10), 1194 => to_unsigned(767, 10), 1195 => to_unsigned(277, 10), 1196 => to_unsigned(542, 10), 1197 => to_unsigned(667, 10), 1198 => to_unsigned(615, 10), 1199 => to_unsigned(650, 10), 1200 => to_unsigned(311, 10), 1201 => to_unsigned(864, 10), 1202 => to_unsigned(265, 10), 1203 => to_unsigned(474, 10), 1204 => to_unsigned(605, 10), 1205 => to_unsigned(1007, 10), 1206 => to_unsigned(891, 10), 1207 => to_unsigned(435, 10), 1208 => to_unsigned(20, 10), 1209 => to_unsigned(924, 10), 1210 => to_unsigned(558, 10), 1211 => to_unsigned(887, 10), 1212 => to_unsigned(920, 10), 1213 => to_unsigned(800, 10), 1214 => to_unsigned(907, 10), 1215 => to_unsigned(63, 10), 1216 => to_unsigned(196, 10), 1217 => to_unsigned(523, 10), 1218 => to_unsigned(539, 10), 1219 => to_unsigned(168, 10), 1220 => to_unsigned(781, 10), 1221 => to_unsigned(766, 10), 1222 => to_unsigned(58, 10), 1223 => to_unsigned(128, 10), 1224 => to_unsigned(164, 10), 1225 => to_unsigned(804, 10), 1226 => to_unsigned(75, 10), 1227 => to_unsigned(661, 10), 1228 => to_unsigned(374, 10), 1229 => to_unsigned(460, 10), 1230 => to_unsigned(733, 10), 1231 => to_unsigned(182, 10), 1232 => to_unsigned(750, 10), 1233 => to_unsigned(1014, 10), 1234 => to_unsigned(984, 10), 1235 => to_unsigned(650, 10), 1236 => to_unsigned(663, 10), 1237 => to_unsigned(770, 10), 1238 => to_unsigned(607, 10), 1239 => to_unsigned(358, 10), 1240 => to_unsigned(476, 10), 1241 => to_unsigned(699, 10), 1242 => to_unsigned(804, 10), 1243 => to_unsigned(375, 10), 1244 => to_unsigned(44, 10), 1245 => to_unsigned(812, 10), 1246 => to_unsigned(342, 10), 1247 => to_unsigned(964, 10), 1248 => to_unsigned(328, 10), 1249 => to_unsigned(902, 10), 1250 => to_unsigned(590, 10), 1251 => to_unsigned(148, 10), 1252 => to_unsigned(440, 10), 1253 => to_unsigned(834, 10), 1254 => to_unsigned(595, 10), 1255 => to_unsigned(371, 10), 1256 => to_unsigned(45, 10), 1257 => to_unsigned(580, 10), 1258 => to_unsigned(255, 10), 1259 => to_unsigned(838, 10), 1260 => to_unsigned(696, 10), 1261 => to_unsigned(104, 10), 1262 => to_unsigned(852, 10), 1263 => to_unsigned(568, 10), 1264 => to_unsigned(673, 10), 1265 => to_unsigned(409, 10), 1266 => to_unsigned(640, 10), 1267 => to_unsigned(905, 10), 1268 => to_unsigned(90, 10), 1269 => to_unsigned(981, 10), 1270 => to_unsigned(717, 10), 1271 => to_unsigned(976, 10), 1272 => to_unsigned(409, 10), 1273 => to_unsigned(906, 10), 1274 => to_unsigned(891, 10), 1275 => to_unsigned(955, 10), 1276 => to_unsigned(831, 10), 1277 => to_unsigned(261, 10), 1278 => to_unsigned(138, 10), 1279 => to_unsigned(924, 10), 1280 => to_unsigned(914, 10), 1281 => to_unsigned(107, 10), 1282 => to_unsigned(702, 10), 1283 => to_unsigned(661, 10), 1284 => to_unsigned(826, 10), 1285 => to_unsigned(687, 10), 1286 => to_unsigned(356, 10), 1287 => to_unsigned(591, 10), 1288 => to_unsigned(450, 10), 1289 => to_unsigned(889, 10), 1290 => to_unsigned(457, 10), 1291 => to_unsigned(57, 10), 1292 => to_unsigned(915, 10), 1293 => to_unsigned(104, 10), 1294 => to_unsigned(697, 10), 1295 => to_unsigned(487, 10), 1296 => to_unsigned(306, 10), 1297 => to_unsigned(750, 10), 1298 => to_unsigned(669, 10), 1299 => to_unsigned(775, 10), 1300 => to_unsigned(523, 10), 1301 => to_unsigned(599, 10), 1302 => to_unsigned(374, 10), 1303 => to_unsigned(72, 10), 1304 => to_unsigned(663, 10), 1305 => to_unsigned(836, 10), 1306 => to_unsigned(384, 10), 1307 => to_unsigned(282, 10), 1308 => to_unsigned(501, 10), 1309 => to_unsigned(340, 10), 1310 => to_unsigned(704, 10), 1311 => to_unsigned(337, 10), 1312 => to_unsigned(223, 10), 1313 => to_unsigned(948, 10), 1314 => to_unsigned(709, 10), 1315 => to_unsigned(775, 10), 1316 => to_unsigned(997, 10), 1317 => to_unsigned(503, 10), 1318 => to_unsigned(293, 10), 1319 => to_unsigned(20, 10), 1320 => to_unsigned(620, 10), 1321 => to_unsigned(361, 10), 1322 => to_unsigned(84, 10), 1323 => to_unsigned(158, 10), 1324 => to_unsigned(399, 10), 1325 => to_unsigned(934, 10), 1326 => to_unsigned(156, 10), 1327 => to_unsigned(305, 10), 1328 => to_unsigned(597, 10), 1329 => to_unsigned(494, 10), 1330 => to_unsigned(985, 10), 1331 => to_unsigned(911, 10), 1332 => to_unsigned(432, 10), 1333 => to_unsigned(99, 10), 1334 => to_unsigned(268, 10), 1335 => to_unsigned(632, 10), 1336 => to_unsigned(23, 10), 1337 => to_unsigned(872, 10), 1338 => to_unsigned(677, 10), 1339 => to_unsigned(368, 10), 1340 => to_unsigned(203, 10), 1341 => to_unsigned(465, 10), 1342 => to_unsigned(472, 10), 1343 => to_unsigned(396, 10), 1344 => to_unsigned(503, 10), 1345 => to_unsigned(426, 10), 1346 => to_unsigned(572, 10), 1347 => to_unsigned(411, 10), 1348 => to_unsigned(992, 10), 1349 => to_unsigned(902, 10), 1350 => to_unsigned(826, 10), 1351 => to_unsigned(630, 10), 1352 => to_unsigned(813, 10), 1353 => to_unsigned(620, 10), 1354 => to_unsigned(744, 10), 1355 => to_unsigned(1001, 10), 1356 => to_unsigned(406, 10), 1357 => to_unsigned(140, 10), 1358 => to_unsigned(341, 10), 1359 => to_unsigned(384, 10), 1360 => to_unsigned(874, 10), 1361 => to_unsigned(156, 10), 1362 => to_unsigned(555, 10), 1363 => to_unsigned(739, 10), 1364 => to_unsigned(1008, 10), 1365 => to_unsigned(449, 10), 1366 => to_unsigned(657, 10), 1367 => to_unsigned(375, 10), 1368 => to_unsigned(25, 10), 1369 => to_unsigned(399, 10), 1370 => to_unsigned(717, 10), 1371 => to_unsigned(119, 10), 1372 => to_unsigned(127, 10), 1373 => to_unsigned(277, 10), 1374 => to_unsigned(2, 10), 1375 => to_unsigned(486, 10), 1376 => to_unsigned(654, 10), 1377 => to_unsigned(20, 10), 1378 => to_unsigned(881, 10), 1379 => to_unsigned(535, 10), 1380 => to_unsigned(34, 10), 1381 => to_unsigned(614, 10), 1382 => to_unsigned(246, 10), 1383 => to_unsigned(328, 10), 1384 => to_unsigned(790, 10), 1385 => to_unsigned(7, 10), 1386 => to_unsigned(820, 10), 1387 => to_unsigned(235, 10), 1388 => to_unsigned(831, 10), 1389 => to_unsigned(1, 10), 1390 => to_unsigned(968, 10), 1391 => to_unsigned(412, 10), 1392 => to_unsigned(987, 10), 1393 => to_unsigned(226, 10), 1394 => to_unsigned(157, 10), 1395 => to_unsigned(954, 10), 1396 => to_unsigned(222, 10), 1397 => to_unsigned(905, 10), 1398 => to_unsigned(60, 10), 1399 => to_unsigned(848, 10), 1400 => to_unsigned(1014, 10), 1401 => to_unsigned(631, 10), 1402 => to_unsigned(232, 10), 1403 => to_unsigned(413, 10), 1404 => to_unsigned(176, 10), 1405 => to_unsigned(857, 10), 1406 => to_unsigned(993, 10), 1407 => to_unsigned(321, 10), 1408 => to_unsigned(929, 10), 1409 => to_unsigned(978, 10), 1410 => to_unsigned(284, 10), 1411 => to_unsigned(816, 10), 1412 => to_unsigned(747, 10), 1413 => to_unsigned(616, 10), 1414 => to_unsigned(565, 10), 1415 => to_unsigned(850, 10), 1416 => to_unsigned(326, 10), 1417 => to_unsigned(547, 10), 1418 => to_unsigned(873, 10), 1419 => to_unsigned(393, 10), 1420 => to_unsigned(280, 10), 1421 => to_unsigned(898, 10), 1422 => to_unsigned(27, 10), 1423 => to_unsigned(880, 10), 1424 => to_unsigned(190, 10), 1425 => to_unsigned(578, 10), 1426 => to_unsigned(79, 10), 1427 => to_unsigned(642, 10), 1428 => to_unsigned(587, 10), 1429 => to_unsigned(795, 10), 1430 => to_unsigned(995, 10), 1431 => to_unsigned(111, 10), 1432 => to_unsigned(878, 10), 1433 => to_unsigned(271, 10), 1434 => to_unsigned(36, 10), 1435 => to_unsigned(343, 10), 1436 => to_unsigned(909, 10), 1437 => to_unsigned(306, 10), 1438 => to_unsigned(329, 10), 1439 => to_unsigned(59, 10), 1440 => to_unsigned(636, 10), 1441 => to_unsigned(659, 10), 1442 => to_unsigned(598, 10), 1443 => to_unsigned(758, 10), 1444 => to_unsigned(101, 10), 1445 => to_unsigned(420, 10), 1446 => to_unsigned(828, 10), 1447 => to_unsigned(655, 10), 1448 => to_unsigned(937, 10), 1449 => to_unsigned(187, 10), 1450 => to_unsigned(94, 10), 1451 => to_unsigned(525, 10), 1452 => to_unsigned(1002, 10), 1453 => to_unsigned(580, 10), 1454 => to_unsigned(578, 10), 1455 => to_unsigned(278, 10), 1456 => to_unsigned(470, 10), 1457 => to_unsigned(971, 10), 1458 => to_unsigned(892, 10), 1459 => to_unsigned(598, 10), 1460 => to_unsigned(605, 10), 1461 => to_unsigned(420, 10), 1462 => to_unsigned(98, 10), 1463 => to_unsigned(480, 10), 1464 => to_unsigned(608, 10), 1465 => to_unsigned(920, 10), 1466 => to_unsigned(824, 10), 1467 => to_unsigned(922, 10), 1468 => to_unsigned(279, 10), 1469 => to_unsigned(104, 10), 1470 => to_unsigned(374, 10), 1471 => to_unsigned(756, 10), 1472 => to_unsigned(722, 10), 1473 => to_unsigned(835, 10), 1474 => to_unsigned(984, 10), 1475 => to_unsigned(338, 10), 1476 => to_unsigned(629, 10), 1477 => to_unsigned(25, 10), 1478 => to_unsigned(799, 10), 1479 => to_unsigned(440, 10), 1480 => to_unsigned(553, 10), 1481 => to_unsigned(268, 10), 1482 => to_unsigned(562, 10), 1483 => to_unsigned(799, 10), 1484 => to_unsigned(160, 10), 1485 => to_unsigned(47, 10), 1486 => to_unsigned(264, 10), 1487 => to_unsigned(903, 10), 1488 => to_unsigned(105, 10), 1489 => to_unsigned(373, 10), 1490 => to_unsigned(666, 10), 1491 => to_unsigned(590, 10), 1492 => to_unsigned(222, 10), 1493 => to_unsigned(40, 10), 1494 => to_unsigned(686, 10), 1495 => to_unsigned(650, 10), 1496 => to_unsigned(843, 10), 1497 => to_unsigned(126, 10), 1498 => to_unsigned(968, 10), 1499 => to_unsigned(943, 10), 1500 => to_unsigned(401, 10), 1501 => to_unsigned(545, 10), 1502 => to_unsigned(35, 10), 1503 => to_unsigned(638, 10), 1504 => to_unsigned(928, 10), 1505 => to_unsigned(755, 10), 1506 => to_unsigned(945, 10), 1507 => to_unsigned(906, 10), 1508 => to_unsigned(846, 10), 1509 => to_unsigned(644, 10), 1510 => to_unsigned(630, 10), 1511 => to_unsigned(960, 10), 1512 => to_unsigned(805, 10), 1513 => to_unsigned(290, 10), 1514 => to_unsigned(53, 10), 1515 => to_unsigned(596, 10), 1516 => to_unsigned(965, 10), 1517 => to_unsigned(638, 10), 1518 => to_unsigned(399, 10), 1519 => to_unsigned(525, 10), 1520 => to_unsigned(710, 10), 1521 => to_unsigned(620, 10), 1522 => to_unsigned(495, 10), 1523 => to_unsigned(302, 10), 1524 => to_unsigned(114, 10), 1525 => to_unsigned(764, 10), 1526 => to_unsigned(195, 10), 1527 => to_unsigned(488, 10), 1528 => to_unsigned(245, 10), 1529 => to_unsigned(172, 10), 1530 => to_unsigned(51, 10), 1531 => to_unsigned(781, 10), 1532 => to_unsigned(781, 10), 1533 => to_unsigned(391, 10), 1534 => to_unsigned(474, 10), 1535 => to_unsigned(690, 10), 1536 => to_unsigned(864, 10), 1537 => to_unsigned(870, 10), 1538 => to_unsigned(794, 10), 1539 => to_unsigned(332, 10), 1540 => to_unsigned(815, 10), 1541 => to_unsigned(111, 10), 1542 => to_unsigned(241, 10), 1543 => to_unsigned(701, 10), 1544 => to_unsigned(407, 10), 1545 => to_unsigned(2, 10), 1546 => to_unsigned(435, 10), 1547 => to_unsigned(979, 10), 1548 => to_unsigned(211, 10), 1549 => to_unsigned(731, 10), 1550 => to_unsigned(137, 10), 1551 => to_unsigned(420, 10), 1552 => to_unsigned(978, 10), 1553 => to_unsigned(288, 10), 1554 => to_unsigned(913, 10), 1555 => to_unsigned(389, 10), 1556 => to_unsigned(670, 10), 1557 => to_unsigned(158, 10), 1558 => to_unsigned(1017, 10), 1559 => to_unsigned(821, 10), 1560 => to_unsigned(769, 10), 1561 => to_unsigned(122, 10), 1562 => to_unsigned(444, 10), 1563 => to_unsigned(73, 10), 1564 => to_unsigned(482, 10), 1565 => to_unsigned(652, 10), 1566 => to_unsigned(697, 10), 1567 => to_unsigned(694, 10), 1568 => to_unsigned(638, 10), 1569 => to_unsigned(200, 10), 1570 => to_unsigned(38, 10), 1571 => to_unsigned(55, 10), 1572 => to_unsigned(574, 10), 1573 => to_unsigned(986, 10), 1574 => to_unsigned(316, 10), 1575 => to_unsigned(395, 10), 1576 => to_unsigned(1011, 10), 1577 => to_unsigned(817, 10), 1578 => to_unsigned(893, 10), 1579 => to_unsigned(452, 10), 1580 => to_unsigned(133, 10), 1581 => to_unsigned(301, 10), 1582 => to_unsigned(289, 10), 1583 => to_unsigned(756, 10), 1584 => to_unsigned(856, 10), 1585 => to_unsigned(972, 10), 1586 => to_unsigned(861, 10), 1587 => to_unsigned(192, 10), 1588 => to_unsigned(219, 10), 1589 => to_unsigned(69, 10), 1590 => to_unsigned(1000, 10), 1591 => to_unsigned(429, 10), 1592 => to_unsigned(850, 10), 1593 => to_unsigned(690, 10), 1594 => to_unsigned(34, 10), 1595 => to_unsigned(506, 10), 1596 => to_unsigned(63, 10), 1597 => to_unsigned(529, 10), 1598 => to_unsigned(909, 10), 1599 => to_unsigned(85, 10), 1600 => to_unsigned(485, 10), 1601 => to_unsigned(970, 10), 1602 => to_unsigned(579, 10), 1603 => to_unsigned(913, 10), 1604 => to_unsigned(122, 10), 1605 => to_unsigned(178, 10), 1606 => to_unsigned(227, 10), 1607 => to_unsigned(588, 10), 1608 => to_unsigned(367, 10), 1609 => to_unsigned(176, 10), 1610 => to_unsigned(450, 10), 1611 => to_unsigned(657, 10), 1612 => to_unsigned(540, 10), 1613 => to_unsigned(272, 10), 1614 => to_unsigned(4, 10), 1615 => to_unsigned(32, 10), 1616 => to_unsigned(689, 10), 1617 => to_unsigned(81, 10), 1618 => to_unsigned(967, 10), 1619 => to_unsigned(18, 10), 1620 => to_unsigned(312, 10), 1621 => to_unsigned(70, 10), 1622 => to_unsigned(962, 10), 1623 => to_unsigned(568, 10), 1624 => to_unsigned(466, 10), 1625 => to_unsigned(870, 10), 1626 => to_unsigned(824, 10), 1627 => to_unsigned(656, 10), 1628 => to_unsigned(742, 10), 1629 => to_unsigned(151, 10), 1630 => to_unsigned(793, 10), 1631 => to_unsigned(822, 10), 1632 => to_unsigned(556, 10), 1633 => to_unsigned(884, 10), 1634 => to_unsigned(87, 10), 1635 => to_unsigned(339, 10), 1636 => to_unsigned(684, 10), 1637 => to_unsigned(927, 10), 1638 => to_unsigned(94, 10), 1639 => to_unsigned(961, 10), 1640 => to_unsigned(97, 10), 1641 => to_unsigned(24, 10), 1642 => to_unsigned(982, 10), 1643 => to_unsigned(929, 10), 1644 => to_unsigned(723, 10), 1645 => to_unsigned(926, 10), 1646 => to_unsigned(1021, 10), 1647 => to_unsigned(602, 10), 1648 => to_unsigned(546, 10), 1649 => to_unsigned(980, 10), 1650 => to_unsigned(1008, 10), 1651 => to_unsigned(740, 10), 1652 => to_unsigned(81, 10), 1653 => to_unsigned(528, 10), 1654 => to_unsigned(303, 10), 1655 => to_unsigned(826, 10), 1656 => to_unsigned(731, 10), 1657 => to_unsigned(857, 10), 1658 => to_unsigned(674, 10), 1659 => to_unsigned(227, 10), 1660 => to_unsigned(507, 10), 1661 => to_unsigned(870, 10), 1662 => to_unsigned(390, 10), 1663 => to_unsigned(30, 10), 1664 => to_unsigned(824, 10), 1665 => to_unsigned(849, 10), 1666 => to_unsigned(845, 10), 1667 => to_unsigned(304, 10), 1668 => to_unsigned(948, 10), 1669 => to_unsigned(493, 10), 1670 => to_unsigned(379, 10), 1671 => to_unsigned(629, 10), 1672 => to_unsigned(130, 10), 1673 => to_unsigned(26, 10), 1674 => to_unsigned(636, 10), 1675 => to_unsigned(951, 10), 1676 => to_unsigned(152, 10), 1677 => to_unsigned(1007, 10), 1678 => to_unsigned(284, 10), 1679 => to_unsigned(968, 10), 1680 => to_unsigned(503, 10), 1681 => to_unsigned(228, 10), 1682 => to_unsigned(204, 10), 1683 => to_unsigned(37, 10), 1684 => to_unsigned(895, 10), 1685 => to_unsigned(1001, 10), 1686 => to_unsigned(965, 10), 1687 => to_unsigned(129, 10), 1688 => to_unsigned(233, 10), 1689 => to_unsigned(808, 10), 1690 => to_unsigned(338, 10), 1691 => to_unsigned(248, 10), 1692 => to_unsigned(170, 10), 1693 => to_unsigned(341, 10), 1694 => to_unsigned(64, 10), 1695 => to_unsigned(336, 10), 1696 => to_unsigned(681, 10), 1697 => to_unsigned(236, 10), 1698 => to_unsigned(39, 10), 1699 => to_unsigned(223, 10), 1700 => to_unsigned(613, 10), 1701 => to_unsigned(108, 10), 1702 => to_unsigned(472, 10), 1703 => to_unsigned(115, 10), 1704 => to_unsigned(539, 10), 1705 => to_unsigned(869, 10), 1706 => to_unsigned(589, 10), 1707 => to_unsigned(668, 10), 1708 => to_unsigned(58, 10), 1709 => to_unsigned(993, 10), 1710 => to_unsigned(961, 10), 1711 => to_unsigned(534, 10), 1712 => to_unsigned(77, 10), 1713 => to_unsigned(270, 10), 1714 => to_unsigned(996, 10), 1715 => to_unsigned(89, 10), 1716 => to_unsigned(416, 10), 1717 => to_unsigned(198, 10), 1718 => to_unsigned(273, 10), 1719 => to_unsigned(39, 10), 1720 => to_unsigned(4, 10), 1721 => to_unsigned(628, 10), 1722 => to_unsigned(154, 10), 1723 => to_unsigned(94, 10), 1724 => to_unsigned(136, 10), 1725 => to_unsigned(142, 10), 1726 => to_unsigned(184, 10), 1727 => to_unsigned(90, 10), 1728 => to_unsigned(785, 10), 1729 => to_unsigned(980, 10), 1730 => to_unsigned(28, 10), 1731 => to_unsigned(811, 10), 1732 => to_unsigned(259, 10), 1733 => to_unsigned(448, 10), 1734 => to_unsigned(12, 10), 1735 => to_unsigned(595, 10), 1736 => to_unsigned(62, 10), 1737 => to_unsigned(638, 10), 1738 => to_unsigned(567, 10), 1739 => to_unsigned(703, 10), 1740 => to_unsigned(442, 10), 1741 => to_unsigned(340, 10), 1742 => to_unsigned(521, 10), 1743 => to_unsigned(936, 10), 1744 => to_unsigned(817, 10), 1745 => to_unsigned(195, 10), 1746 => to_unsigned(607, 10), 1747 => to_unsigned(269, 10), 1748 => to_unsigned(108, 10), 1749 => to_unsigned(343, 10), 1750 => to_unsigned(274, 10), 1751 => to_unsigned(255, 10), 1752 => to_unsigned(572, 10), 1753 => to_unsigned(327, 10), 1754 => to_unsigned(684, 10), 1755 => to_unsigned(432, 10), 1756 => to_unsigned(811, 10), 1757 => to_unsigned(982, 10), 1758 => to_unsigned(489, 10), 1759 => to_unsigned(695, 10), 1760 => to_unsigned(683, 10), 1761 => to_unsigned(52, 10), 1762 => to_unsigned(181, 10), 1763 => to_unsigned(406, 10), 1764 => to_unsigned(322, 10), 1765 => to_unsigned(1006, 10), 1766 => to_unsigned(566, 10), 1767 => to_unsigned(965, 10), 1768 => to_unsigned(591, 10), 1769 => to_unsigned(1023, 10), 1770 => to_unsigned(903, 10), 1771 => to_unsigned(889, 10), 1772 => to_unsigned(225, 10), 1773 => to_unsigned(986, 10), 1774 => to_unsigned(918, 10), 1775 => to_unsigned(674, 10), 1776 => to_unsigned(220, 10), 1777 => to_unsigned(260, 10), 1778 => to_unsigned(1001, 10), 1779 => to_unsigned(999, 10), 1780 => to_unsigned(439, 10), 1781 => to_unsigned(73, 10), 1782 => to_unsigned(80, 10), 1783 => to_unsigned(956, 10), 1784 => to_unsigned(282, 10), 1785 => to_unsigned(805, 10), 1786 => to_unsigned(894, 10), 1787 => to_unsigned(45, 10), 1788 => to_unsigned(890, 10), 1789 => to_unsigned(486, 10), 1790 => to_unsigned(324, 10), 1791 => to_unsigned(395, 10), 1792 => to_unsigned(701, 10), 1793 => to_unsigned(402, 10), 1794 => to_unsigned(992, 10), 1795 => to_unsigned(215, 10), 1796 => to_unsigned(400, 10), 1797 => to_unsigned(127, 10), 1798 => to_unsigned(141, 10), 1799 => to_unsigned(259, 10), 1800 => to_unsigned(240, 10), 1801 => to_unsigned(396, 10), 1802 => to_unsigned(123, 10), 1803 => to_unsigned(945, 10), 1804 => to_unsigned(839, 10), 1805 => to_unsigned(860, 10), 1806 => to_unsigned(282, 10), 1807 => to_unsigned(620, 10), 1808 => to_unsigned(91, 10), 1809 => to_unsigned(392, 10), 1810 => to_unsigned(869, 10), 1811 => to_unsigned(157, 10), 1812 => to_unsigned(613, 10), 1813 => to_unsigned(229, 10), 1814 => to_unsigned(441, 10), 1815 => to_unsigned(699, 10), 1816 => to_unsigned(48, 10), 1817 => to_unsigned(143, 10), 1818 => to_unsigned(1017, 10), 1819 => to_unsigned(737, 10), 1820 => to_unsigned(518, 10), 1821 => to_unsigned(199, 10), 1822 => to_unsigned(455, 10), 1823 => to_unsigned(164, 10), 1824 => to_unsigned(148, 10), 1825 => to_unsigned(424, 10), 1826 => to_unsigned(176, 10), 1827 => to_unsigned(235, 10), 1828 => to_unsigned(84, 10), 1829 => to_unsigned(417, 10), 1830 => to_unsigned(675, 10), 1831 => to_unsigned(214, 10), 1832 => to_unsigned(570, 10), 1833 => to_unsigned(909, 10), 1834 => to_unsigned(942, 10), 1835 => to_unsigned(451, 10), 1836 => to_unsigned(370, 10), 1837 => to_unsigned(842, 10), 1838 => to_unsigned(32, 10), 1839 => to_unsigned(896, 10), 1840 => to_unsigned(264, 10), 1841 => to_unsigned(62, 10), 1842 => to_unsigned(419, 10), 1843 => to_unsigned(706, 10), 1844 => to_unsigned(10, 10), 1845 => to_unsigned(176, 10), 1846 => to_unsigned(287, 10), 1847 => to_unsigned(941, 10), 1848 => to_unsigned(979, 10), 1849 => to_unsigned(446, 10), 1850 => to_unsigned(501, 10), 1851 => to_unsigned(339, 10), 1852 => to_unsigned(867, 10), 1853 => to_unsigned(646, 10), 1854 => to_unsigned(440, 10), 1855 => to_unsigned(467, 10), 1856 => to_unsigned(315, 10), 1857 => to_unsigned(230, 10), 1858 => to_unsigned(502, 10), 1859 => to_unsigned(956, 10), 1860 => to_unsigned(849, 10), 1861 => to_unsigned(318, 10), 1862 => to_unsigned(282, 10), 1863 => to_unsigned(250, 10), 1864 => to_unsigned(770, 10), 1865 => to_unsigned(875, 10), 1866 => to_unsigned(344, 10), 1867 => to_unsigned(473, 10), 1868 => to_unsigned(808, 10), 1869 => to_unsigned(499, 10), 1870 => to_unsigned(113, 10), 1871 => to_unsigned(340, 10), 1872 => to_unsigned(970, 10), 1873 => to_unsigned(691, 10), 1874 => to_unsigned(914, 10), 1875 => to_unsigned(189, 10), 1876 => to_unsigned(741, 10), 1877 => to_unsigned(839, 10), 1878 => to_unsigned(236, 10), 1879 => to_unsigned(516, 10), 1880 => to_unsigned(161, 10), 1881 => to_unsigned(903, 10), 1882 => to_unsigned(553, 10), 1883 => to_unsigned(770, 10), 1884 => to_unsigned(446, 10), 1885 => to_unsigned(938, 10), 1886 => to_unsigned(760, 10), 1887 => to_unsigned(924, 10), 1888 => to_unsigned(537, 10), 1889 => to_unsigned(56, 10), 1890 => to_unsigned(25, 10), 1891 => to_unsigned(982, 10), 1892 => to_unsigned(433, 10), 1893 => to_unsigned(181, 10), 1894 => to_unsigned(221, 10), 1895 => to_unsigned(958, 10), 1896 => to_unsigned(218, 10), 1897 => to_unsigned(958, 10), 1898 => to_unsigned(829, 10), 1899 => to_unsigned(371, 10), 1900 => to_unsigned(829, 10), 1901 => to_unsigned(638, 10), 1902 => to_unsigned(120, 10), 1903 => to_unsigned(600, 10), 1904 => to_unsigned(123, 10), 1905 => to_unsigned(275, 10), 1906 => to_unsigned(736, 10), 1907 => to_unsigned(809, 10), 1908 => to_unsigned(880, 10), 1909 => to_unsigned(1008, 10), 1910 => to_unsigned(535, 10), 1911 => to_unsigned(53, 10), 1912 => to_unsigned(524, 10), 1913 => to_unsigned(736, 10), 1914 => to_unsigned(78, 10), 1915 => to_unsigned(937, 10), 1916 => to_unsigned(305, 10), 1917 => to_unsigned(540, 10), 1918 => to_unsigned(952, 10), 1919 => to_unsigned(551, 10), 1920 => to_unsigned(473, 10), 1921 => to_unsigned(73, 10), 1922 => to_unsigned(460, 10), 1923 => to_unsigned(753, 10), 1924 => to_unsigned(269, 10), 1925 => to_unsigned(1016, 10), 1926 => to_unsigned(805, 10), 1927 => to_unsigned(475, 10), 1928 => to_unsigned(840, 10), 1929 => to_unsigned(553, 10), 1930 => to_unsigned(574, 10), 1931 => to_unsigned(808, 10), 1932 => to_unsigned(545, 10), 1933 => to_unsigned(765, 10), 1934 => to_unsigned(0, 10), 1935 => to_unsigned(15, 10), 1936 => to_unsigned(294, 10), 1937 => to_unsigned(419, 10), 1938 => to_unsigned(275, 10), 1939 => to_unsigned(484, 10), 1940 => to_unsigned(806, 10), 1941 => to_unsigned(865, 10), 1942 => to_unsigned(103, 10), 1943 => to_unsigned(461, 10), 1944 => to_unsigned(548, 10), 1945 => to_unsigned(619, 10), 1946 => to_unsigned(320, 10), 1947 => to_unsigned(168, 10), 1948 => to_unsigned(394, 10), 1949 => to_unsigned(295, 10), 1950 => to_unsigned(232, 10), 1951 => to_unsigned(274, 10), 1952 => to_unsigned(366, 10), 1953 => to_unsigned(940, 10), 1954 => to_unsigned(422, 10), 1955 => to_unsigned(3, 10), 1956 => to_unsigned(739, 10), 1957 => to_unsigned(997, 10), 1958 => to_unsigned(253, 10), 1959 => to_unsigned(754, 10), 1960 => to_unsigned(767, 10), 1961 => to_unsigned(334, 10), 1962 => to_unsigned(978, 10), 1963 => to_unsigned(593, 10), 1964 => to_unsigned(245, 10), 1965 => to_unsigned(133, 10), 1966 => to_unsigned(73, 10), 1967 => to_unsigned(819, 10), 1968 => to_unsigned(591, 10), 1969 => to_unsigned(458, 10), 1970 => to_unsigned(934, 10), 1971 => to_unsigned(884, 10), 1972 => to_unsigned(158, 10), 1973 => to_unsigned(645, 10), 1974 => to_unsigned(203, 10), 1975 => to_unsigned(278, 10), 1976 => to_unsigned(489, 10), 1977 => to_unsigned(892, 10), 1978 => to_unsigned(599, 10), 1979 => to_unsigned(921, 10), 1980 => to_unsigned(789, 10), 1981 => to_unsigned(71, 10), 1982 => to_unsigned(945, 10), 1983 => to_unsigned(529, 10), 1984 => to_unsigned(862, 10), 1985 => to_unsigned(714, 10), 1986 => to_unsigned(897, 10), 1987 => to_unsigned(329, 10), 1988 => to_unsigned(367, 10), 1989 => to_unsigned(648, 10), 1990 => to_unsigned(901, 10), 1991 => to_unsigned(970, 10), 1992 => to_unsigned(996, 10), 1993 => to_unsigned(605, 10), 1994 => to_unsigned(430, 10), 1995 => to_unsigned(440, 10), 1996 => to_unsigned(699, 10), 1997 => to_unsigned(369, 10), 1998 => to_unsigned(288, 10), 1999 => to_unsigned(225, 10), 2000 => to_unsigned(511, 10), 2001 => to_unsigned(653, 10), 2002 => to_unsigned(277, 10), 2003 => to_unsigned(890, 10), 2004 => to_unsigned(538, 10), 2005 => to_unsigned(636, 10), 2006 => to_unsigned(904, 10), 2007 => to_unsigned(925, 10), 2008 => to_unsigned(748, 10), 2009 => to_unsigned(698, 10), 2010 => to_unsigned(962, 10), 2011 => to_unsigned(279, 10), 2012 => to_unsigned(258, 10), 2013 => to_unsigned(725, 10), 2014 => to_unsigned(827, 10), 2015 => to_unsigned(731, 10), 2016 => to_unsigned(537, 10), 2017 => to_unsigned(192, 10), 2018 => to_unsigned(403, 10), 2019 => to_unsigned(131, 10), 2020 => to_unsigned(628, 10), 2021 => to_unsigned(941, 10), 2022 => to_unsigned(483, 10), 2023 => to_unsigned(1015, 10), 2024 => to_unsigned(962, 10), 2025 => to_unsigned(707, 10), 2026 => to_unsigned(229, 10), 2027 => to_unsigned(449, 10), 2028 => to_unsigned(243, 10), 2029 => to_unsigned(585, 10), 2030 => to_unsigned(96, 10), 2031 => to_unsigned(230, 10), 2032 => to_unsigned(181, 10), 2033 => to_unsigned(602, 10), 2034 => to_unsigned(620, 10), 2035 => to_unsigned(515, 10), 2036 => to_unsigned(615, 10), 2037 => to_unsigned(319, 10), 2038 => to_unsigned(543, 10), 2039 => to_unsigned(166, 10), 2040 => to_unsigned(124, 10), 2041 => to_unsigned(510, 10), 2042 => to_unsigned(100, 10), 2043 => to_unsigned(284, 10), 2044 => to_unsigned(772, 10), 2045 => to_unsigned(178, 10), 2046 => to_unsigned(319, 10), 2047 => to_unsigned(393, 10))
    );

begin

	-- Generate main clock signal
    clock_gen : process
        constant clock_period : time := 20 ns;
	begin
		wait for clock_period / 2;
		clock <= not clock;
	end process clock_gen;

    test : process
        constant fragment_size : integer := vnir_row_width / vnir_lvds_n_channels;
        variable tests_passed : boolean := true;
    begin
        wait until rising_edge(clock);

        config.window_blue <= (lo => 0, hi => 0);
        config.window_red  <= (lo => 1, hi => 1);
        config.window_nir  <= (lo => 2, hi => 2);
        read_config <= '1';
        wait until rising_edge(clock);
        read_config <= '0';

        report "Uploading started";
        start <= '1';
        wait until rising_edge(clock);
        start <= '0';

        fragment_available <= '1';
        for w in 0 to 2 loop
            for f in 0 to fragment_size-1 loop
                for i in 0 to vnir_lvds_n_channels-1 loop
                    fragment(i) <= data(w)(f + fragment_size * i);
                    -- fragment(i) <= to_unsigned(f, 10);
                end loop;
                wait until rising_edge(clock);
            end loop;
        end loop;
        fragment_available <= '0';
        report "Uploading finished";

        wait until rising_edge(clock);
        wait until rising_edge(clock);
        wait until rising_edge(clock);

        wait until rising_edge(clock);
        tests_passed := tests_passed and test_report(rows_available = '1', "rows available");
        tests_passed := tests_passed and test_report(rows.nir = data(0), "NIR row");
        tests_passed := tests_passed and test_report(rows.blue = data(1), "blue row");
        tests_passed := tests_passed and test_report(rows.red = data(2), "red row");

        test_end(tests_passed);
        wait;
    end process test;

    row_collector_component : row_collector port map (
        clock => clock,
        config => config,
        read_config => read_config,
        start => start,
        fragment => fragment,
        fragment_available => fragment_available,
        rows => rows,
        rows_available => rows_available
    );

end tests;
